* Substrate SPICE library
* This is a generated file. Be careful when editing manually: this file may be overwritten.


.SUBCKT sram_sp_hstrap BR VDD VSS BL VNB VPB

  X0 BL VNB BL VNB sky130_fd_pr__special_nfet_pass l=0.140 nf=1 w=0.140

  X1 BL VNB BL VNB sky130_fd_pr__special_nfet_pass l=0.140 nf=1 w=0.140


.ENDS sram_sp_hstrap

.SUBCKT sky130_fd_sc_hs__mux2_4 A0 A1 S VGND VNB VPB VPWR X

  X0 a_27_368# S VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X1 a_722_391# A0 a_193_241# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X2 a_722_391# S VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X3 VGND a_27_368# a_937_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X4 a_193_241# A1 a_936_391# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X5 a_709_119# S VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X6 a_709_119# A1 a_193_241# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X7 X a_193_241# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X8 X a_193_241# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 VPWR a_27_368# a_936_391# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X10 X a_193_241# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X11 a_193_241# A0 a_722_391# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X12 a_937_119# A0 a_193_241# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X13 a_936_391# a_27_368# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X14 VGND a_193_241# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X15 VPWR a_193_241# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X16 VPWR S a_722_391# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X17 a_936_391# A1 a_193_241# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X18 a_193_241# A0 a_937_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X19 a_193_241# A1 a_709_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X20 X a_193_241# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X21 VGND a_193_241# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X22 a_27_368# S VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X23 a_937_119# a_27_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X24 VPWR a_193_241# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X25 VGND S a_709_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640


.ENDS sky130_fd_sc_hs__mux2_4

.SUBCKT sky130_fd_sc_hs__mux2_4_wrapper A0 A1 S VGND VNB VPB VPWR X

  X0 A0 A1 S VGND VNB VPB VPWR X sky130_fd_sc_hs__mux2_4

.ENDS sky130_fd_sc_hs__mux2_4_wrapper

.SUBCKT mos_w2000_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=2.000


.ENDS mos_w2000_l150_m1_nf1_id0

.SUBCKT mos_w2500_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.500


.ENDS mos_w2500_l150_m1_nf1_id1

.SUBCKT nand2 vdd vss a b y

  Xn1 x a vss vss mos_w2000_l150_m1_nf1_id0
  Xn2 y b x vss mos_w2000_l150_m1_nf1_id0
  Xp1 y a vdd vdd mos_w2500_l150_m1_nf1_id1
  Xp2 y b vdd vdd mos_w2500_l150_m1_nf1_id1

.ENDS nand2

.SUBCKT mos_w2180_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.180


.ENDS mos_w2180_l150_m1_nf1_id1

.SUBCKT mos_w880_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.880


.ENDS mos_w880_l150_m1_nf1_id0

.SUBCKT folded_inv_8 vdd vss a y

  XMP0 y a vdd vdd mos_w2180_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w880_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w2180_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w880_l150_m1_nf1_id0

.ENDS folded_inv_8

.SUBCKT and2_1 vdd a b y yb vss

  X0 vdd vss a b yb nand2
  X0_1 vdd vss yb y folded_inv_8

.ENDS and2_1

.SUBCKT mos_w700_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.700


.ENDS mos_w700_l150_m1_nf1_id1

.SUBCKT mos_w700_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.700


.ENDS mos_w700_l150_m1_nf1_id0

.SUBCKT multi_finger_inv_10 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_10

.SUBCKT multi_finger_inv_11 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP19 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN7 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_11

.SUBCKT multi_finger_inv_12 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP19 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP20 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP21 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP22 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP23 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP24 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP25 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP26 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP27 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP28 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP29 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP30 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP31 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP32 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP33 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP34 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP35 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN7 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN8 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN9 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN10 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN11 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN12 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN13 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_12

.SUBCKT multi_finger_inv_13 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP19 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP20 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP21 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP22 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP23 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP24 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP25 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP26 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP27 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP28 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP29 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP30 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP31 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP32 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP33 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP34 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP35 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP36 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP37 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP38 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP39 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP40 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP41 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP42 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP43 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP44 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP45 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP46 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP47 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP48 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP49 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP50 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP51 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP52 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP53 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP54 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP55 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP56 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP57 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP58 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP59 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP60 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP61 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP62 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP63 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP64 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN7 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN8 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN9 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN10 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN11 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN12 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN13 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN14 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN15 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN16 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN17 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN18 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN19 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN20 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN21 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN22 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN23 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN24 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN25 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_13

.SUBCKT multi_finger_inv_14 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP19 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP20 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP21 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP22 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP23 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP24 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP25 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP26 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP27 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP28 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP29 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP30 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP31 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP32 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP33 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP34 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP35 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP36 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP37 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP38 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP39 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP40 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP41 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP42 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP43 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP44 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP45 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP46 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP47 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP48 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP49 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP50 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP51 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP52 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP53 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP54 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP55 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP56 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP57 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP58 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP59 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP60 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP61 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP62 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP63 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP64 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP65 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP66 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP67 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP68 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP69 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP70 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP71 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP72 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP73 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP74 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP75 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP76 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP77 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP78 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP79 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP80 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP81 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP82 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP83 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP84 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP85 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP86 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP87 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP88 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP89 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP90 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP91 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP92 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP93 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP94 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP95 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP96 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP97 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP98 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP99 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP100 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP101 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP102 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP103 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP104 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP105 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP106 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP107 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP108 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP109 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP110 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP111 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP112 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP113 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP114 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP115 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP116 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN7 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN8 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN9 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN10 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN11 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN12 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN13 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN14 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN15 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN16 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN17 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN18 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN19 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN20 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN21 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN22 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN23 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN24 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN25 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN26 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN27 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN28 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN29 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN30 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN31 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN32 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN33 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN34 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN35 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN36 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN37 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN38 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN39 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN40 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN41 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN42 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN43 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN44 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN45 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN46 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_14

.SUBCKT multi_finger_inv_15 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP19 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP20 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP21 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP22 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP23 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP24 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP25 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP26 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP27 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP28 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP29 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP30 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP31 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP32 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP33 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP34 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP35 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP36 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP37 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP38 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP39 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP40 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP41 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP42 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP43 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP44 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP45 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP46 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP47 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP48 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP49 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP50 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP51 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP52 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP53 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP54 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP55 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP56 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP57 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP58 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP59 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP60 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP61 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP62 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP63 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP64 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP65 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP66 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP67 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP68 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP69 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP70 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP71 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP72 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP73 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP74 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP75 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP76 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP77 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP78 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP79 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP80 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP81 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP82 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP83 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP84 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP85 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP86 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP87 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP88 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP89 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP90 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP91 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP92 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP93 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP94 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP95 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP96 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP97 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP98 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP99 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP100 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP101 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP102 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP103 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP104 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP105 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP106 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP107 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP108 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP109 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP110 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP111 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP112 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP113 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP114 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP115 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP116 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP117 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP118 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP119 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP120 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP121 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP122 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP123 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP124 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP125 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP126 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP127 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP128 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP129 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP130 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP131 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP132 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP133 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP134 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP135 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP136 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP137 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP138 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP139 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP140 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP141 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP142 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP143 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP144 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP145 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP146 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP147 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP148 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP149 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP150 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP151 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP152 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP153 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP154 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP155 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP156 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP157 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP158 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP159 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP160 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP161 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP162 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP163 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP164 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP165 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP166 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP167 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP168 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP169 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP170 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP171 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP172 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP173 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP174 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP175 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP176 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP177 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP178 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP179 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP180 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP181 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP182 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP183 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP184 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP185 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP186 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP187 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP188 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP189 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP190 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP191 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP192 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP193 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP194 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP195 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP196 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP197 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP198 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP199 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP200 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP201 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP202 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP203 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP204 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP205 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP206 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP207 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP208 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP209 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP210 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN7 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN8 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN9 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN10 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN11 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN12 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN13 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN14 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN15 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN16 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN17 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN18 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN19 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN20 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN21 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN22 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN23 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN24 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN25 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN26 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN27 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN28 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN29 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN30 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN31 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN32 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN33 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN34 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN35 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN36 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN37 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN38 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN39 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN40 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN41 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN42 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN43 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN44 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN45 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN46 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN47 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN48 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN49 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN50 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN51 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN52 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN53 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN54 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN55 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN56 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN57 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN58 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN59 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN60 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN61 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN62 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN63 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN64 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN65 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN66 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN67 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN68 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN69 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN70 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN71 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN72 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN73 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN74 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN75 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN76 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN77 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN78 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN79 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN80 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN81 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN82 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN83 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN84 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_15

.SUBCKT decoder_stage_5 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y[12] y[13] y[14] y[15] y[16] y[17] y[18] y[19] y[20] y[21] y[22] y[23] y[24] y[25] y[26] y[27] y[28] y[29] y[30] y[31] y[32] y[33] y[34] y[35] y[36] y[37] y[38] y[39] y[40] y[41] y[42] y[43] y[44] y[45] y[46] y[47] y[48] y[49] y[50] y[51] y[52] y[53] y[54] y[55] y[56] y[57] y[58] y[59] y[60] y[61] y[62] y[63] y[64] y[65] y[66] y[67] y[68] y[69] y[70] y[71] y[72] y[73] y[74] y[75] y[76] y[77] y[78] y[79] y[80] y[81] y[82] y[83] y[84] y[85] y[86] y[87] y[88] y[89] y[90] y[91] y[92] y[93] y[94] y[95] y[96] y[97] y[98] y[99] y[100] y[101] y[102] y[103] y[104] y[105] y[106] y[107] y[108] y[109] y[110] y[111] y[112] y[113] y[114] y[115] y[116] y[117] y[118] y[119] y[120] y[121] y[122] y[123] y[124] y[125] y[126] y[127] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] y_b[12] y_b[13] y_b[14] y_b[15] y_b[16] y_b[17] y_b[18] y_b[19] y_b[20] y_b[21] y_b[22] y_b[23] y_b[24] y_b[25] y_b[26] y_b[27] y_b[28] y_b[29] y_b[30] y_b[31] y_b[32] y_b[33] y_b[34] y_b[35] y_b[36] y_b[37] y_b[38] y_b[39] y_b[40] y_b[41] y_b[42] y_b[43] y_b[44] y_b[45] y_b[46] y_b[47] y_b[48] y_b[49] y_b[50] y_b[51] y_b[52] y_b[53] y_b[54] y_b[55] y_b[56] y_b[57] y_b[58] y_b[59] y_b[60] y_b[61] y_b[62] y_b[63] y_b[64] y_b[65] y_b[66] y_b[67] y_b[68] y_b[69] y_b[70] y_b[71] y_b[72] y_b[73] y_b[74] y_b[75] y_b[76] y_b[77] y_b[78] y_b[79] y_b[80] y_b[81] y_b[82] y_b[83] y_b[84] y_b[85] y_b[86] y_b[87] y_b[88] y_b[89] y_b[90] y_b[91] y_b[92] y_b[93] y_b[94] y_b[95] y_b[96] y_b[97] y_b[98] y_b[99] y_b[100] y_b[101] y_b[102] y_b[103] y_b[104] y_b[105] y_b[106] y_b[107] y_b[108] y_b[109] y_b[110] y_b[111] y_b[112] y_b[113] y_b[114] y_b[115] y_b[116] y_b[117] y_b[118] y_b[119] y_b[120] y_b[121] y_b[122] y_b[123] y_b[124] y_b[125] y_b[126] y_b[127] predecode_0_0 predecode_0_1 predecode_0_2 predecode_0_3 predecode_0_4 predecode_0_5 predecode_0_6 predecode_0_7 predecode_0_8 predecode_0_9 predecode_0_10 predecode_0_11 predecode_0_12 predecode_0_13 predecode_0_14 predecode_0_15 predecode_1_0 predecode_1_1 predecode_1_2 predecode_1_3 predecode_1_4 predecode_1_5 predecode_1_6 predecode_1_7

  Xgate_0_0_0 vdd predecode_0_0 predecode_1_0 x_0[0] y_b_noconn_0_0_0 vss and2_1
  Xgate_0_1_0 vdd predecode_0_1 predecode_1_0 x_0[1] y_b_noconn_0_1_0 vss and2_1
  Xgate_0_2_0 vdd predecode_0_2 predecode_1_0 x_0[2] y_b_noconn_0_2_0 vss and2_1
  Xgate_0_3_0 vdd predecode_0_3 predecode_1_0 x_0[3] y_b_noconn_0_3_0 vss and2_1
  Xgate_0_4_0 vdd predecode_0_4 predecode_1_0 x_0[4] y_b_noconn_0_4_0 vss and2_1
  Xgate_0_5_0 vdd predecode_0_5 predecode_1_0 x_0[5] y_b_noconn_0_5_0 vss and2_1
  Xgate_0_6_0 vdd predecode_0_6 predecode_1_0 x_0[6] y_b_noconn_0_6_0 vss and2_1
  Xgate_0_7_0 vdd predecode_0_7 predecode_1_0 x_0[7] y_b_noconn_0_7_0 vss and2_1
  Xgate_0_8_0 vdd predecode_0_8 predecode_1_0 x_0[8] y_b_noconn_0_8_0 vss and2_1
  Xgate_0_9_0 vdd predecode_0_9 predecode_1_0 x_0[9] y_b_noconn_0_9_0 vss and2_1
  Xgate_0_10_0 vdd predecode_0_10 predecode_1_0 x_0[10] y_b_noconn_0_10_0 vss and2_1
  Xgate_0_11_0 vdd predecode_0_11 predecode_1_0 x_0[11] y_b_noconn_0_11_0 vss and2_1
  Xgate_0_12_0 vdd predecode_0_12 predecode_1_0 x_0[12] y_b_noconn_0_12_0 vss and2_1
  Xgate_0_13_0 vdd predecode_0_13 predecode_1_0 x_0[13] y_b_noconn_0_13_0 vss and2_1
  Xgate_0_14_0 vdd predecode_0_14 predecode_1_0 x_0[14] y_b_noconn_0_14_0 vss and2_1
  Xgate_0_15_0 vdd predecode_0_15 predecode_1_0 x_0[15] y_b_noconn_0_15_0 vss and2_1
  Xgate_0_16_0 vdd predecode_0_0 predecode_1_1 x_0[16] y_b_noconn_0_16_0 vss and2_1
  Xgate_0_17_0 vdd predecode_0_1 predecode_1_1 x_0[17] y_b_noconn_0_17_0 vss and2_1
  Xgate_0_18_0 vdd predecode_0_2 predecode_1_1 x_0[18] y_b_noconn_0_18_0 vss and2_1
  Xgate_0_19_0 vdd predecode_0_3 predecode_1_1 x_0[19] y_b_noconn_0_19_0 vss and2_1
  Xgate_0_20_0 vdd predecode_0_4 predecode_1_1 x_0[20] y_b_noconn_0_20_0 vss and2_1
  Xgate_0_21_0 vdd predecode_0_5 predecode_1_1 x_0[21] y_b_noconn_0_21_0 vss and2_1
  Xgate_0_22_0 vdd predecode_0_6 predecode_1_1 x_0[22] y_b_noconn_0_22_0 vss and2_1
  Xgate_0_23_0 vdd predecode_0_7 predecode_1_1 x_0[23] y_b_noconn_0_23_0 vss and2_1
  Xgate_0_24_0 vdd predecode_0_8 predecode_1_1 x_0[24] y_b_noconn_0_24_0 vss and2_1
  Xgate_0_25_0 vdd predecode_0_9 predecode_1_1 x_0[25] y_b_noconn_0_25_0 vss and2_1
  Xgate_0_26_0 vdd predecode_0_10 predecode_1_1 x_0[26] y_b_noconn_0_26_0 vss and2_1
  Xgate_0_27_0 vdd predecode_0_11 predecode_1_1 x_0[27] y_b_noconn_0_27_0 vss and2_1
  Xgate_0_28_0 vdd predecode_0_12 predecode_1_1 x_0[28] y_b_noconn_0_28_0 vss and2_1
  Xgate_0_29_0 vdd predecode_0_13 predecode_1_1 x_0[29] y_b_noconn_0_29_0 vss and2_1
  Xgate_0_30_0 vdd predecode_0_14 predecode_1_1 x_0[30] y_b_noconn_0_30_0 vss and2_1
  Xgate_0_31_0 vdd predecode_0_15 predecode_1_1 x_0[31] y_b_noconn_0_31_0 vss and2_1
  Xgate_0_32_0 vdd predecode_0_0 predecode_1_2 x_0[32] y_b_noconn_0_32_0 vss and2_1
  Xgate_0_33_0 vdd predecode_0_1 predecode_1_2 x_0[33] y_b_noconn_0_33_0 vss and2_1
  Xgate_0_34_0 vdd predecode_0_2 predecode_1_2 x_0[34] y_b_noconn_0_34_0 vss and2_1
  Xgate_0_35_0 vdd predecode_0_3 predecode_1_2 x_0[35] y_b_noconn_0_35_0 vss and2_1
  Xgate_0_36_0 vdd predecode_0_4 predecode_1_2 x_0[36] y_b_noconn_0_36_0 vss and2_1
  Xgate_0_37_0 vdd predecode_0_5 predecode_1_2 x_0[37] y_b_noconn_0_37_0 vss and2_1
  Xgate_0_38_0 vdd predecode_0_6 predecode_1_2 x_0[38] y_b_noconn_0_38_0 vss and2_1
  Xgate_0_39_0 vdd predecode_0_7 predecode_1_2 x_0[39] y_b_noconn_0_39_0 vss and2_1
  Xgate_0_40_0 vdd predecode_0_8 predecode_1_2 x_0[40] y_b_noconn_0_40_0 vss and2_1
  Xgate_0_41_0 vdd predecode_0_9 predecode_1_2 x_0[41] y_b_noconn_0_41_0 vss and2_1
  Xgate_0_42_0 vdd predecode_0_10 predecode_1_2 x_0[42] y_b_noconn_0_42_0 vss and2_1
  Xgate_0_43_0 vdd predecode_0_11 predecode_1_2 x_0[43] y_b_noconn_0_43_0 vss and2_1
  Xgate_0_44_0 vdd predecode_0_12 predecode_1_2 x_0[44] y_b_noconn_0_44_0 vss and2_1
  Xgate_0_45_0 vdd predecode_0_13 predecode_1_2 x_0[45] y_b_noconn_0_45_0 vss and2_1
  Xgate_0_46_0 vdd predecode_0_14 predecode_1_2 x_0[46] y_b_noconn_0_46_0 vss and2_1
  Xgate_0_47_0 vdd predecode_0_15 predecode_1_2 x_0[47] y_b_noconn_0_47_0 vss and2_1
  Xgate_0_48_0 vdd predecode_0_0 predecode_1_3 x_0[48] y_b_noconn_0_48_0 vss and2_1
  Xgate_0_49_0 vdd predecode_0_1 predecode_1_3 x_0[49] y_b_noconn_0_49_0 vss and2_1
  Xgate_0_50_0 vdd predecode_0_2 predecode_1_3 x_0[50] y_b_noconn_0_50_0 vss and2_1
  Xgate_0_51_0 vdd predecode_0_3 predecode_1_3 x_0[51] y_b_noconn_0_51_0 vss and2_1
  Xgate_0_52_0 vdd predecode_0_4 predecode_1_3 x_0[52] y_b_noconn_0_52_0 vss and2_1
  Xgate_0_53_0 vdd predecode_0_5 predecode_1_3 x_0[53] y_b_noconn_0_53_0 vss and2_1
  Xgate_0_54_0 vdd predecode_0_6 predecode_1_3 x_0[54] y_b_noconn_0_54_0 vss and2_1
  Xgate_0_55_0 vdd predecode_0_7 predecode_1_3 x_0[55] y_b_noconn_0_55_0 vss and2_1
  Xgate_0_56_0 vdd predecode_0_8 predecode_1_3 x_0[56] y_b_noconn_0_56_0 vss and2_1
  Xgate_0_57_0 vdd predecode_0_9 predecode_1_3 x_0[57] y_b_noconn_0_57_0 vss and2_1
  Xgate_0_58_0 vdd predecode_0_10 predecode_1_3 x_0[58] y_b_noconn_0_58_0 vss and2_1
  Xgate_0_59_0 vdd predecode_0_11 predecode_1_3 x_0[59] y_b_noconn_0_59_0 vss and2_1
  Xgate_0_60_0 vdd predecode_0_12 predecode_1_3 x_0[60] y_b_noconn_0_60_0 vss and2_1
  Xgate_0_61_0 vdd predecode_0_13 predecode_1_3 x_0[61] y_b_noconn_0_61_0 vss and2_1
  Xgate_0_62_0 vdd predecode_0_14 predecode_1_3 x_0[62] y_b_noconn_0_62_0 vss and2_1
  Xgate_0_63_0 vdd predecode_0_15 predecode_1_3 x_0[63] y_b_noconn_0_63_0 vss and2_1
  Xgate_0_64_0 vdd predecode_0_0 predecode_1_4 x_0[64] y_b_noconn_0_64_0 vss and2_1
  Xgate_0_65_0 vdd predecode_0_1 predecode_1_4 x_0[65] y_b_noconn_0_65_0 vss and2_1
  Xgate_0_66_0 vdd predecode_0_2 predecode_1_4 x_0[66] y_b_noconn_0_66_0 vss and2_1
  Xgate_0_67_0 vdd predecode_0_3 predecode_1_4 x_0[67] y_b_noconn_0_67_0 vss and2_1
  Xgate_0_68_0 vdd predecode_0_4 predecode_1_4 x_0[68] y_b_noconn_0_68_0 vss and2_1
  Xgate_0_69_0 vdd predecode_0_5 predecode_1_4 x_0[69] y_b_noconn_0_69_0 vss and2_1
  Xgate_0_70_0 vdd predecode_0_6 predecode_1_4 x_0[70] y_b_noconn_0_70_0 vss and2_1
  Xgate_0_71_0 vdd predecode_0_7 predecode_1_4 x_0[71] y_b_noconn_0_71_0 vss and2_1
  Xgate_0_72_0 vdd predecode_0_8 predecode_1_4 x_0[72] y_b_noconn_0_72_0 vss and2_1
  Xgate_0_73_0 vdd predecode_0_9 predecode_1_4 x_0[73] y_b_noconn_0_73_0 vss and2_1
  Xgate_0_74_0 vdd predecode_0_10 predecode_1_4 x_0[74] y_b_noconn_0_74_0 vss and2_1
  Xgate_0_75_0 vdd predecode_0_11 predecode_1_4 x_0[75] y_b_noconn_0_75_0 vss and2_1
  Xgate_0_76_0 vdd predecode_0_12 predecode_1_4 x_0[76] y_b_noconn_0_76_0 vss and2_1
  Xgate_0_77_0 vdd predecode_0_13 predecode_1_4 x_0[77] y_b_noconn_0_77_0 vss and2_1
  Xgate_0_78_0 vdd predecode_0_14 predecode_1_4 x_0[78] y_b_noconn_0_78_0 vss and2_1
  Xgate_0_79_0 vdd predecode_0_15 predecode_1_4 x_0[79] y_b_noconn_0_79_0 vss and2_1
  Xgate_0_80_0 vdd predecode_0_0 predecode_1_5 x_0[80] y_b_noconn_0_80_0 vss and2_1
  Xgate_0_81_0 vdd predecode_0_1 predecode_1_5 x_0[81] y_b_noconn_0_81_0 vss and2_1
  Xgate_0_82_0 vdd predecode_0_2 predecode_1_5 x_0[82] y_b_noconn_0_82_0 vss and2_1
  Xgate_0_83_0 vdd predecode_0_3 predecode_1_5 x_0[83] y_b_noconn_0_83_0 vss and2_1
  Xgate_0_84_0 vdd predecode_0_4 predecode_1_5 x_0[84] y_b_noconn_0_84_0 vss and2_1
  Xgate_0_85_0 vdd predecode_0_5 predecode_1_5 x_0[85] y_b_noconn_0_85_0 vss and2_1
  Xgate_0_86_0 vdd predecode_0_6 predecode_1_5 x_0[86] y_b_noconn_0_86_0 vss and2_1
  Xgate_0_87_0 vdd predecode_0_7 predecode_1_5 x_0[87] y_b_noconn_0_87_0 vss and2_1
  Xgate_0_88_0 vdd predecode_0_8 predecode_1_5 x_0[88] y_b_noconn_0_88_0 vss and2_1
  Xgate_0_89_0 vdd predecode_0_9 predecode_1_5 x_0[89] y_b_noconn_0_89_0 vss and2_1
  Xgate_0_90_0 vdd predecode_0_10 predecode_1_5 x_0[90] y_b_noconn_0_90_0 vss and2_1
  Xgate_0_91_0 vdd predecode_0_11 predecode_1_5 x_0[91] y_b_noconn_0_91_0 vss and2_1
  Xgate_0_92_0 vdd predecode_0_12 predecode_1_5 x_0[92] y_b_noconn_0_92_0 vss and2_1
  Xgate_0_93_0 vdd predecode_0_13 predecode_1_5 x_0[93] y_b_noconn_0_93_0 vss and2_1
  Xgate_0_94_0 vdd predecode_0_14 predecode_1_5 x_0[94] y_b_noconn_0_94_0 vss and2_1
  Xgate_0_95_0 vdd predecode_0_15 predecode_1_5 x_0[95] y_b_noconn_0_95_0 vss and2_1
  Xgate_0_96_0 vdd predecode_0_0 predecode_1_6 x_0[96] y_b_noconn_0_96_0 vss and2_1
  Xgate_0_97_0 vdd predecode_0_1 predecode_1_6 x_0[97] y_b_noconn_0_97_0 vss and2_1
  Xgate_0_98_0 vdd predecode_0_2 predecode_1_6 x_0[98] y_b_noconn_0_98_0 vss and2_1
  Xgate_0_99_0 vdd predecode_0_3 predecode_1_6 x_0[99] y_b_noconn_0_99_0 vss and2_1
  Xgate_0_100_0 vdd predecode_0_4 predecode_1_6 x_0[100] y_b_noconn_0_100_0 vss and2_1
  Xgate_0_101_0 vdd predecode_0_5 predecode_1_6 x_0[101] y_b_noconn_0_101_0 vss and2_1
  Xgate_0_102_0 vdd predecode_0_6 predecode_1_6 x_0[102] y_b_noconn_0_102_0 vss and2_1
  Xgate_0_103_0 vdd predecode_0_7 predecode_1_6 x_0[103] y_b_noconn_0_103_0 vss and2_1
  Xgate_0_104_0 vdd predecode_0_8 predecode_1_6 x_0[104] y_b_noconn_0_104_0 vss and2_1
  Xgate_0_105_0 vdd predecode_0_9 predecode_1_6 x_0[105] y_b_noconn_0_105_0 vss and2_1
  Xgate_0_106_0 vdd predecode_0_10 predecode_1_6 x_0[106] y_b_noconn_0_106_0 vss and2_1
  Xgate_0_107_0 vdd predecode_0_11 predecode_1_6 x_0[107] y_b_noconn_0_107_0 vss and2_1
  Xgate_0_108_0 vdd predecode_0_12 predecode_1_6 x_0[108] y_b_noconn_0_108_0 vss and2_1
  Xgate_0_109_0 vdd predecode_0_13 predecode_1_6 x_0[109] y_b_noconn_0_109_0 vss and2_1
  Xgate_0_110_0 vdd predecode_0_14 predecode_1_6 x_0[110] y_b_noconn_0_110_0 vss and2_1
  Xgate_0_111_0 vdd predecode_0_15 predecode_1_6 x_0[111] y_b_noconn_0_111_0 vss and2_1
  Xgate_0_112_0 vdd predecode_0_0 predecode_1_7 x_0[112] y_b_noconn_0_112_0 vss and2_1
  Xgate_0_113_0 vdd predecode_0_1 predecode_1_7 x_0[113] y_b_noconn_0_113_0 vss and2_1
  Xgate_0_114_0 vdd predecode_0_2 predecode_1_7 x_0[114] y_b_noconn_0_114_0 vss and2_1
  Xgate_0_115_0 vdd predecode_0_3 predecode_1_7 x_0[115] y_b_noconn_0_115_0 vss and2_1
  Xgate_0_116_0 vdd predecode_0_4 predecode_1_7 x_0[116] y_b_noconn_0_116_0 vss and2_1
  Xgate_0_117_0 vdd predecode_0_5 predecode_1_7 x_0[117] y_b_noconn_0_117_0 vss and2_1
  Xgate_0_118_0 vdd predecode_0_6 predecode_1_7 x_0[118] y_b_noconn_0_118_0 vss and2_1
  Xgate_0_119_0 vdd predecode_0_7 predecode_1_7 x_0[119] y_b_noconn_0_119_0 vss and2_1
  Xgate_0_120_0 vdd predecode_0_8 predecode_1_7 x_0[120] y_b_noconn_0_120_0 vss and2_1
  Xgate_0_121_0 vdd predecode_0_9 predecode_1_7 x_0[121] y_b_noconn_0_121_0 vss and2_1
  Xgate_0_122_0 vdd predecode_0_10 predecode_1_7 x_0[122] y_b_noconn_0_122_0 vss and2_1
  Xgate_0_123_0 vdd predecode_0_11 predecode_1_7 x_0[123] y_b_noconn_0_123_0 vss and2_1
  Xgate_0_124_0 vdd predecode_0_12 predecode_1_7 x_0[124] y_b_noconn_0_124_0 vss and2_1
  Xgate_0_125_0 vdd predecode_0_13 predecode_1_7 x_0[125] y_b_noconn_0_125_0 vss and2_1
  Xgate_0_126_0 vdd predecode_0_14 predecode_1_7 x_0[126] y_b_noconn_0_126_0 vss and2_1
  Xgate_0_127_0 vdd predecode_0_15 predecode_1_7 x_0[127] y_b_noconn_0_127_0 vss and2_1
  Xgate_1_0_0 vdd vss x_0[0] x_1[0] multi_finger_inv_10
  Xgate_1_1_0 vdd vss x_0[1] x_1[1] multi_finger_inv_10
  Xgate_1_2_0 vdd vss x_0[2] x_1[2] multi_finger_inv_10
  Xgate_1_3_0 vdd vss x_0[3] x_1[3] multi_finger_inv_10
  Xgate_1_4_0 vdd vss x_0[4] x_1[4] multi_finger_inv_10
  Xgate_1_5_0 vdd vss x_0[5] x_1[5] multi_finger_inv_10
  Xgate_1_6_0 vdd vss x_0[6] x_1[6] multi_finger_inv_10
  Xgate_1_7_0 vdd vss x_0[7] x_1[7] multi_finger_inv_10
  Xgate_1_8_0 vdd vss x_0[8] x_1[8] multi_finger_inv_10
  Xgate_1_9_0 vdd vss x_0[9] x_1[9] multi_finger_inv_10
  Xgate_1_10_0 vdd vss x_0[10] x_1[10] multi_finger_inv_10
  Xgate_1_11_0 vdd vss x_0[11] x_1[11] multi_finger_inv_10
  Xgate_1_12_0 vdd vss x_0[12] x_1[12] multi_finger_inv_10
  Xgate_1_13_0 vdd vss x_0[13] x_1[13] multi_finger_inv_10
  Xgate_1_14_0 vdd vss x_0[14] x_1[14] multi_finger_inv_10
  Xgate_1_15_0 vdd vss x_0[15] x_1[15] multi_finger_inv_10
  Xgate_1_16_0 vdd vss x_0[16] x_1[16] multi_finger_inv_10
  Xgate_1_17_0 vdd vss x_0[17] x_1[17] multi_finger_inv_10
  Xgate_1_18_0 vdd vss x_0[18] x_1[18] multi_finger_inv_10
  Xgate_1_19_0 vdd vss x_0[19] x_1[19] multi_finger_inv_10
  Xgate_1_20_0 vdd vss x_0[20] x_1[20] multi_finger_inv_10
  Xgate_1_21_0 vdd vss x_0[21] x_1[21] multi_finger_inv_10
  Xgate_1_22_0 vdd vss x_0[22] x_1[22] multi_finger_inv_10
  Xgate_1_23_0 vdd vss x_0[23] x_1[23] multi_finger_inv_10
  Xgate_1_24_0 vdd vss x_0[24] x_1[24] multi_finger_inv_10
  Xgate_1_25_0 vdd vss x_0[25] x_1[25] multi_finger_inv_10
  Xgate_1_26_0 vdd vss x_0[26] x_1[26] multi_finger_inv_10
  Xgate_1_27_0 vdd vss x_0[27] x_1[27] multi_finger_inv_10
  Xgate_1_28_0 vdd vss x_0[28] x_1[28] multi_finger_inv_10
  Xgate_1_29_0 vdd vss x_0[29] x_1[29] multi_finger_inv_10
  Xgate_1_30_0 vdd vss x_0[30] x_1[30] multi_finger_inv_10
  Xgate_1_31_0 vdd vss x_0[31] x_1[31] multi_finger_inv_10
  Xgate_1_32_0 vdd vss x_0[32] x_1[32] multi_finger_inv_10
  Xgate_1_33_0 vdd vss x_0[33] x_1[33] multi_finger_inv_10
  Xgate_1_34_0 vdd vss x_0[34] x_1[34] multi_finger_inv_10
  Xgate_1_35_0 vdd vss x_0[35] x_1[35] multi_finger_inv_10
  Xgate_1_36_0 vdd vss x_0[36] x_1[36] multi_finger_inv_10
  Xgate_1_37_0 vdd vss x_0[37] x_1[37] multi_finger_inv_10
  Xgate_1_38_0 vdd vss x_0[38] x_1[38] multi_finger_inv_10
  Xgate_1_39_0 vdd vss x_0[39] x_1[39] multi_finger_inv_10
  Xgate_1_40_0 vdd vss x_0[40] x_1[40] multi_finger_inv_10
  Xgate_1_41_0 vdd vss x_0[41] x_1[41] multi_finger_inv_10
  Xgate_1_42_0 vdd vss x_0[42] x_1[42] multi_finger_inv_10
  Xgate_1_43_0 vdd vss x_0[43] x_1[43] multi_finger_inv_10
  Xgate_1_44_0 vdd vss x_0[44] x_1[44] multi_finger_inv_10
  Xgate_1_45_0 vdd vss x_0[45] x_1[45] multi_finger_inv_10
  Xgate_1_46_0 vdd vss x_0[46] x_1[46] multi_finger_inv_10
  Xgate_1_47_0 vdd vss x_0[47] x_1[47] multi_finger_inv_10
  Xgate_1_48_0 vdd vss x_0[48] x_1[48] multi_finger_inv_10
  Xgate_1_49_0 vdd vss x_0[49] x_1[49] multi_finger_inv_10
  Xgate_1_50_0 vdd vss x_0[50] x_1[50] multi_finger_inv_10
  Xgate_1_51_0 vdd vss x_0[51] x_1[51] multi_finger_inv_10
  Xgate_1_52_0 vdd vss x_0[52] x_1[52] multi_finger_inv_10
  Xgate_1_53_0 vdd vss x_0[53] x_1[53] multi_finger_inv_10
  Xgate_1_54_0 vdd vss x_0[54] x_1[54] multi_finger_inv_10
  Xgate_1_55_0 vdd vss x_0[55] x_1[55] multi_finger_inv_10
  Xgate_1_56_0 vdd vss x_0[56] x_1[56] multi_finger_inv_10
  Xgate_1_57_0 vdd vss x_0[57] x_1[57] multi_finger_inv_10
  Xgate_1_58_0 vdd vss x_0[58] x_1[58] multi_finger_inv_10
  Xgate_1_59_0 vdd vss x_0[59] x_1[59] multi_finger_inv_10
  Xgate_1_60_0 vdd vss x_0[60] x_1[60] multi_finger_inv_10
  Xgate_1_61_0 vdd vss x_0[61] x_1[61] multi_finger_inv_10
  Xgate_1_62_0 vdd vss x_0[62] x_1[62] multi_finger_inv_10
  Xgate_1_63_0 vdd vss x_0[63] x_1[63] multi_finger_inv_10
  Xgate_1_64_0 vdd vss x_0[64] x_1[64] multi_finger_inv_10
  Xgate_1_65_0 vdd vss x_0[65] x_1[65] multi_finger_inv_10
  Xgate_1_66_0 vdd vss x_0[66] x_1[66] multi_finger_inv_10
  Xgate_1_67_0 vdd vss x_0[67] x_1[67] multi_finger_inv_10
  Xgate_1_68_0 vdd vss x_0[68] x_1[68] multi_finger_inv_10
  Xgate_1_69_0 vdd vss x_0[69] x_1[69] multi_finger_inv_10
  Xgate_1_70_0 vdd vss x_0[70] x_1[70] multi_finger_inv_10
  Xgate_1_71_0 vdd vss x_0[71] x_1[71] multi_finger_inv_10
  Xgate_1_72_0 vdd vss x_0[72] x_1[72] multi_finger_inv_10
  Xgate_1_73_0 vdd vss x_0[73] x_1[73] multi_finger_inv_10
  Xgate_1_74_0 vdd vss x_0[74] x_1[74] multi_finger_inv_10
  Xgate_1_75_0 vdd vss x_0[75] x_1[75] multi_finger_inv_10
  Xgate_1_76_0 vdd vss x_0[76] x_1[76] multi_finger_inv_10
  Xgate_1_77_0 vdd vss x_0[77] x_1[77] multi_finger_inv_10
  Xgate_1_78_0 vdd vss x_0[78] x_1[78] multi_finger_inv_10
  Xgate_1_79_0 vdd vss x_0[79] x_1[79] multi_finger_inv_10
  Xgate_1_80_0 vdd vss x_0[80] x_1[80] multi_finger_inv_10
  Xgate_1_81_0 vdd vss x_0[81] x_1[81] multi_finger_inv_10
  Xgate_1_82_0 vdd vss x_0[82] x_1[82] multi_finger_inv_10
  Xgate_1_83_0 vdd vss x_0[83] x_1[83] multi_finger_inv_10
  Xgate_1_84_0 vdd vss x_0[84] x_1[84] multi_finger_inv_10
  Xgate_1_85_0 vdd vss x_0[85] x_1[85] multi_finger_inv_10
  Xgate_1_86_0 vdd vss x_0[86] x_1[86] multi_finger_inv_10
  Xgate_1_87_0 vdd vss x_0[87] x_1[87] multi_finger_inv_10
  Xgate_1_88_0 vdd vss x_0[88] x_1[88] multi_finger_inv_10
  Xgate_1_89_0 vdd vss x_0[89] x_1[89] multi_finger_inv_10
  Xgate_1_90_0 vdd vss x_0[90] x_1[90] multi_finger_inv_10
  Xgate_1_91_0 vdd vss x_0[91] x_1[91] multi_finger_inv_10
  Xgate_1_92_0 vdd vss x_0[92] x_1[92] multi_finger_inv_10
  Xgate_1_93_0 vdd vss x_0[93] x_1[93] multi_finger_inv_10
  Xgate_1_94_0 vdd vss x_0[94] x_1[94] multi_finger_inv_10
  Xgate_1_95_0 vdd vss x_0[95] x_1[95] multi_finger_inv_10
  Xgate_1_96_0 vdd vss x_0[96] x_1[96] multi_finger_inv_10
  Xgate_1_97_0 vdd vss x_0[97] x_1[97] multi_finger_inv_10
  Xgate_1_98_0 vdd vss x_0[98] x_1[98] multi_finger_inv_10
  Xgate_1_99_0 vdd vss x_0[99] x_1[99] multi_finger_inv_10
  Xgate_1_100_0 vdd vss x_0[100] x_1[100] multi_finger_inv_10
  Xgate_1_101_0 vdd vss x_0[101] x_1[101] multi_finger_inv_10
  Xgate_1_102_0 vdd vss x_0[102] x_1[102] multi_finger_inv_10
  Xgate_1_103_0 vdd vss x_0[103] x_1[103] multi_finger_inv_10
  Xgate_1_104_0 vdd vss x_0[104] x_1[104] multi_finger_inv_10
  Xgate_1_105_0 vdd vss x_0[105] x_1[105] multi_finger_inv_10
  Xgate_1_106_0 vdd vss x_0[106] x_1[106] multi_finger_inv_10
  Xgate_1_107_0 vdd vss x_0[107] x_1[107] multi_finger_inv_10
  Xgate_1_108_0 vdd vss x_0[108] x_1[108] multi_finger_inv_10
  Xgate_1_109_0 vdd vss x_0[109] x_1[109] multi_finger_inv_10
  Xgate_1_110_0 vdd vss x_0[110] x_1[110] multi_finger_inv_10
  Xgate_1_111_0 vdd vss x_0[111] x_1[111] multi_finger_inv_10
  Xgate_1_112_0 vdd vss x_0[112] x_1[112] multi_finger_inv_10
  Xgate_1_113_0 vdd vss x_0[113] x_1[113] multi_finger_inv_10
  Xgate_1_114_0 vdd vss x_0[114] x_1[114] multi_finger_inv_10
  Xgate_1_115_0 vdd vss x_0[115] x_1[115] multi_finger_inv_10
  Xgate_1_116_0 vdd vss x_0[116] x_1[116] multi_finger_inv_10
  Xgate_1_117_0 vdd vss x_0[117] x_1[117] multi_finger_inv_10
  Xgate_1_118_0 vdd vss x_0[118] x_1[118] multi_finger_inv_10
  Xgate_1_119_0 vdd vss x_0[119] x_1[119] multi_finger_inv_10
  Xgate_1_120_0 vdd vss x_0[120] x_1[120] multi_finger_inv_10
  Xgate_1_121_0 vdd vss x_0[121] x_1[121] multi_finger_inv_10
  Xgate_1_122_0 vdd vss x_0[122] x_1[122] multi_finger_inv_10
  Xgate_1_123_0 vdd vss x_0[123] x_1[123] multi_finger_inv_10
  Xgate_1_124_0 vdd vss x_0[124] x_1[124] multi_finger_inv_10
  Xgate_1_125_0 vdd vss x_0[125] x_1[125] multi_finger_inv_10
  Xgate_1_126_0 vdd vss x_0[126] x_1[126] multi_finger_inv_10
  Xgate_1_127_0 vdd vss x_0[127] x_1[127] multi_finger_inv_10
  Xgate_2_0_0 vdd vss x_1[0] x_2[0] multi_finger_inv_11
  Xgate_2_1_0 vdd vss x_1[1] x_2[1] multi_finger_inv_11
  Xgate_2_2_0 vdd vss x_1[2] x_2[2] multi_finger_inv_11
  Xgate_2_3_0 vdd vss x_1[3] x_2[3] multi_finger_inv_11
  Xgate_2_4_0 vdd vss x_1[4] x_2[4] multi_finger_inv_11
  Xgate_2_5_0 vdd vss x_1[5] x_2[5] multi_finger_inv_11
  Xgate_2_6_0 vdd vss x_1[6] x_2[6] multi_finger_inv_11
  Xgate_2_7_0 vdd vss x_1[7] x_2[7] multi_finger_inv_11
  Xgate_2_8_0 vdd vss x_1[8] x_2[8] multi_finger_inv_11
  Xgate_2_9_0 vdd vss x_1[9] x_2[9] multi_finger_inv_11
  Xgate_2_10_0 vdd vss x_1[10] x_2[10] multi_finger_inv_11
  Xgate_2_11_0 vdd vss x_1[11] x_2[11] multi_finger_inv_11
  Xgate_2_12_0 vdd vss x_1[12] x_2[12] multi_finger_inv_11
  Xgate_2_13_0 vdd vss x_1[13] x_2[13] multi_finger_inv_11
  Xgate_2_14_0 vdd vss x_1[14] x_2[14] multi_finger_inv_11
  Xgate_2_15_0 vdd vss x_1[15] x_2[15] multi_finger_inv_11
  Xgate_2_16_0 vdd vss x_1[16] x_2[16] multi_finger_inv_11
  Xgate_2_17_0 vdd vss x_1[17] x_2[17] multi_finger_inv_11
  Xgate_2_18_0 vdd vss x_1[18] x_2[18] multi_finger_inv_11
  Xgate_2_19_0 vdd vss x_1[19] x_2[19] multi_finger_inv_11
  Xgate_2_20_0 vdd vss x_1[20] x_2[20] multi_finger_inv_11
  Xgate_2_21_0 vdd vss x_1[21] x_2[21] multi_finger_inv_11
  Xgate_2_22_0 vdd vss x_1[22] x_2[22] multi_finger_inv_11
  Xgate_2_23_0 vdd vss x_1[23] x_2[23] multi_finger_inv_11
  Xgate_2_24_0 vdd vss x_1[24] x_2[24] multi_finger_inv_11
  Xgate_2_25_0 vdd vss x_1[25] x_2[25] multi_finger_inv_11
  Xgate_2_26_0 vdd vss x_1[26] x_2[26] multi_finger_inv_11
  Xgate_2_27_0 vdd vss x_1[27] x_2[27] multi_finger_inv_11
  Xgate_2_28_0 vdd vss x_1[28] x_2[28] multi_finger_inv_11
  Xgate_2_29_0 vdd vss x_1[29] x_2[29] multi_finger_inv_11
  Xgate_2_30_0 vdd vss x_1[30] x_2[30] multi_finger_inv_11
  Xgate_2_31_0 vdd vss x_1[31] x_2[31] multi_finger_inv_11
  Xgate_2_32_0 vdd vss x_1[32] x_2[32] multi_finger_inv_11
  Xgate_2_33_0 vdd vss x_1[33] x_2[33] multi_finger_inv_11
  Xgate_2_34_0 vdd vss x_1[34] x_2[34] multi_finger_inv_11
  Xgate_2_35_0 vdd vss x_1[35] x_2[35] multi_finger_inv_11
  Xgate_2_36_0 vdd vss x_1[36] x_2[36] multi_finger_inv_11
  Xgate_2_37_0 vdd vss x_1[37] x_2[37] multi_finger_inv_11
  Xgate_2_38_0 vdd vss x_1[38] x_2[38] multi_finger_inv_11
  Xgate_2_39_0 vdd vss x_1[39] x_2[39] multi_finger_inv_11
  Xgate_2_40_0 vdd vss x_1[40] x_2[40] multi_finger_inv_11
  Xgate_2_41_0 vdd vss x_1[41] x_2[41] multi_finger_inv_11
  Xgate_2_42_0 vdd vss x_1[42] x_2[42] multi_finger_inv_11
  Xgate_2_43_0 vdd vss x_1[43] x_2[43] multi_finger_inv_11
  Xgate_2_44_0 vdd vss x_1[44] x_2[44] multi_finger_inv_11
  Xgate_2_45_0 vdd vss x_1[45] x_2[45] multi_finger_inv_11
  Xgate_2_46_0 vdd vss x_1[46] x_2[46] multi_finger_inv_11
  Xgate_2_47_0 vdd vss x_1[47] x_2[47] multi_finger_inv_11
  Xgate_2_48_0 vdd vss x_1[48] x_2[48] multi_finger_inv_11
  Xgate_2_49_0 vdd vss x_1[49] x_2[49] multi_finger_inv_11
  Xgate_2_50_0 vdd vss x_1[50] x_2[50] multi_finger_inv_11
  Xgate_2_51_0 vdd vss x_1[51] x_2[51] multi_finger_inv_11
  Xgate_2_52_0 vdd vss x_1[52] x_2[52] multi_finger_inv_11
  Xgate_2_53_0 vdd vss x_1[53] x_2[53] multi_finger_inv_11
  Xgate_2_54_0 vdd vss x_1[54] x_2[54] multi_finger_inv_11
  Xgate_2_55_0 vdd vss x_1[55] x_2[55] multi_finger_inv_11
  Xgate_2_56_0 vdd vss x_1[56] x_2[56] multi_finger_inv_11
  Xgate_2_57_0 vdd vss x_1[57] x_2[57] multi_finger_inv_11
  Xgate_2_58_0 vdd vss x_1[58] x_2[58] multi_finger_inv_11
  Xgate_2_59_0 vdd vss x_1[59] x_2[59] multi_finger_inv_11
  Xgate_2_60_0 vdd vss x_1[60] x_2[60] multi_finger_inv_11
  Xgate_2_61_0 vdd vss x_1[61] x_2[61] multi_finger_inv_11
  Xgate_2_62_0 vdd vss x_1[62] x_2[62] multi_finger_inv_11
  Xgate_2_63_0 vdd vss x_1[63] x_2[63] multi_finger_inv_11
  Xgate_2_64_0 vdd vss x_1[64] x_2[64] multi_finger_inv_11
  Xgate_2_65_0 vdd vss x_1[65] x_2[65] multi_finger_inv_11
  Xgate_2_66_0 vdd vss x_1[66] x_2[66] multi_finger_inv_11
  Xgate_2_67_0 vdd vss x_1[67] x_2[67] multi_finger_inv_11
  Xgate_2_68_0 vdd vss x_1[68] x_2[68] multi_finger_inv_11
  Xgate_2_69_0 vdd vss x_1[69] x_2[69] multi_finger_inv_11
  Xgate_2_70_0 vdd vss x_1[70] x_2[70] multi_finger_inv_11
  Xgate_2_71_0 vdd vss x_1[71] x_2[71] multi_finger_inv_11
  Xgate_2_72_0 vdd vss x_1[72] x_2[72] multi_finger_inv_11
  Xgate_2_73_0 vdd vss x_1[73] x_2[73] multi_finger_inv_11
  Xgate_2_74_0 vdd vss x_1[74] x_2[74] multi_finger_inv_11
  Xgate_2_75_0 vdd vss x_1[75] x_2[75] multi_finger_inv_11
  Xgate_2_76_0 vdd vss x_1[76] x_2[76] multi_finger_inv_11
  Xgate_2_77_0 vdd vss x_1[77] x_2[77] multi_finger_inv_11
  Xgate_2_78_0 vdd vss x_1[78] x_2[78] multi_finger_inv_11
  Xgate_2_79_0 vdd vss x_1[79] x_2[79] multi_finger_inv_11
  Xgate_2_80_0 vdd vss x_1[80] x_2[80] multi_finger_inv_11
  Xgate_2_81_0 vdd vss x_1[81] x_2[81] multi_finger_inv_11
  Xgate_2_82_0 vdd vss x_1[82] x_2[82] multi_finger_inv_11
  Xgate_2_83_0 vdd vss x_1[83] x_2[83] multi_finger_inv_11
  Xgate_2_84_0 vdd vss x_1[84] x_2[84] multi_finger_inv_11
  Xgate_2_85_0 vdd vss x_1[85] x_2[85] multi_finger_inv_11
  Xgate_2_86_0 vdd vss x_1[86] x_2[86] multi_finger_inv_11
  Xgate_2_87_0 vdd vss x_1[87] x_2[87] multi_finger_inv_11
  Xgate_2_88_0 vdd vss x_1[88] x_2[88] multi_finger_inv_11
  Xgate_2_89_0 vdd vss x_1[89] x_2[89] multi_finger_inv_11
  Xgate_2_90_0 vdd vss x_1[90] x_2[90] multi_finger_inv_11
  Xgate_2_91_0 vdd vss x_1[91] x_2[91] multi_finger_inv_11
  Xgate_2_92_0 vdd vss x_1[92] x_2[92] multi_finger_inv_11
  Xgate_2_93_0 vdd vss x_1[93] x_2[93] multi_finger_inv_11
  Xgate_2_94_0 vdd vss x_1[94] x_2[94] multi_finger_inv_11
  Xgate_2_95_0 vdd vss x_1[95] x_2[95] multi_finger_inv_11
  Xgate_2_96_0 vdd vss x_1[96] x_2[96] multi_finger_inv_11
  Xgate_2_97_0 vdd vss x_1[97] x_2[97] multi_finger_inv_11
  Xgate_2_98_0 vdd vss x_1[98] x_2[98] multi_finger_inv_11
  Xgate_2_99_0 vdd vss x_1[99] x_2[99] multi_finger_inv_11
  Xgate_2_100_0 vdd vss x_1[100] x_2[100] multi_finger_inv_11
  Xgate_2_101_0 vdd vss x_1[101] x_2[101] multi_finger_inv_11
  Xgate_2_102_0 vdd vss x_1[102] x_2[102] multi_finger_inv_11
  Xgate_2_103_0 vdd vss x_1[103] x_2[103] multi_finger_inv_11
  Xgate_2_104_0 vdd vss x_1[104] x_2[104] multi_finger_inv_11
  Xgate_2_105_0 vdd vss x_1[105] x_2[105] multi_finger_inv_11
  Xgate_2_106_0 vdd vss x_1[106] x_2[106] multi_finger_inv_11
  Xgate_2_107_0 vdd vss x_1[107] x_2[107] multi_finger_inv_11
  Xgate_2_108_0 vdd vss x_1[108] x_2[108] multi_finger_inv_11
  Xgate_2_109_0 vdd vss x_1[109] x_2[109] multi_finger_inv_11
  Xgate_2_110_0 vdd vss x_1[110] x_2[110] multi_finger_inv_11
  Xgate_2_111_0 vdd vss x_1[111] x_2[111] multi_finger_inv_11
  Xgate_2_112_0 vdd vss x_1[112] x_2[112] multi_finger_inv_11
  Xgate_2_113_0 vdd vss x_1[113] x_2[113] multi_finger_inv_11
  Xgate_2_114_0 vdd vss x_1[114] x_2[114] multi_finger_inv_11
  Xgate_2_115_0 vdd vss x_1[115] x_2[115] multi_finger_inv_11
  Xgate_2_116_0 vdd vss x_1[116] x_2[116] multi_finger_inv_11
  Xgate_2_117_0 vdd vss x_1[117] x_2[117] multi_finger_inv_11
  Xgate_2_118_0 vdd vss x_1[118] x_2[118] multi_finger_inv_11
  Xgate_2_119_0 vdd vss x_1[119] x_2[119] multi_finger_inv_11
  Xgate_2_120_0 vdd vss x_1[120] x_2[120] multi_finger_inv_11
  Xgate_2_121_0 vdd vss x_1[121] x_2[121] multi_finger_inv_11
  Xgate_2_122_0 vdd vss x_1[122] x_2[122] multi_finger_inv_11
  Xgate_2_123_0 vdd vss x_1[123] x_2[123] multi_finger_inv_11
  Xgate_2_124_0 vdd vss x_1[124] x_2[124] multi_finger_inv_11
  Xgate_2_125_0 vdd vss x_1[125] x_2[125] multi_finger_inv_11
  Xgate_2_126_0 vdd vss x_1[126] x_2[126] multi_finger_inv_11
  Xgate_2_127_0 vdd vss x_1[127] x_2[127] multi_finger_inv_11
  Xgate_3_0_0 vdd vss x_2[0] x_3[0] multi_finger_inv_12
  Xgate_3_1_0 vdd vss x_2[1] x_3[1] multi_finger_inv_12
  Xgate_3_2_0 vdd vss x_2[2] x_3[2] multi_finger_inv_12
  Xgate_3_3_0 vdd vss x_2[3] x_3[3] multi_finger_inv_12
  Xgate_3_4_0 vdd vss x_2[4] x_3[4] multi_finger_inv_12
  Xgate_3_5_0 vdd vss x_2[5] x_3[5] multi_finger_inv_12
  Xgate_3_6_0 vdd vss x_2[6] x_3[6] multi_finger_inv_12
  Xgate_3_7_0 vdd vss x_2[7] x_3[7] multi_finger_inv_12
  Xgate_3_8_0 vdd vss x_2[8] x_3[8] multi_finger_inv_12
  Xgate_3_9_0 vdd vss x_2[9] x_3[9] multi_finger_inv_12
  Xgate_3_10_0 vdd vss x_2[10] x_3[10] multi_finger_inv_12
  Xgate_3_11_0 vdd vss x_2[11] x_3[11] multi_finger_inv_12
  Xgate_3_12_0 vdd vss x_2[12] x_3[12] multi_finger_inv_12
  Xgate_3_13_0 vdd vss x_2[13] x_3[13] multi_finger_inv_12
  Xgate_3_14_0 vdd vss x_2[14] x_3[14] multi_finger_inv_12
  Xgate_3_15_0 vdd vss x_2[15] x_3[15] multi_finger_inv_12
  Xgate_3_16_0 vdd vss x_2[16] x_3[16] multi_finger_inv_12
  Xgate_3_17_0 vdd vss x_2[17] x_3[17] multi_finger_inv_12
  Xgate_3_18_0 vdd vss x_2[18] x_3[18] multi_finger_inv_12
  Xgate_3_19_0 vdd vss x_2[19] x_3[19] multi_finger_inv_12
  Xgate_3_20_0 vdd vss x_2[20] x_3[20] multi_finger_inv_12
  Xgate_3_21_0 vdd vss x_2[21] x_3[21] multi_finger_inv_12
  Xgate_3_22_0 vdd vss x_2[22] x_3[22] multi_finger_inv_12
  Xgate_3_23_0 vdd vss x_2[23] x_3[23] multi_finger_inv_12
  Xgate_3_24_0 vdd vss x_2[24] x_3[24] multi_finger_inv_12
  Xgate_3_25_0 vdd vss x_2[25] x_3[25] multi_finger_inv_12
  Xgate_3_26_0 vdd vss x_2[26] x_3[26] multi_finger_inv_12
  Xgate_3_27_0 vdd vss x_2[27] x_3[27] multi_finger_inv_12
  Xgate_3_28_0 vdd vss x_2[28] x_3[28] multi_finger_inv_12
  Xgate_3_29_0 vdd vss x_2[29] x_3[29] multi_finger_inv_12
  Xgate_3_30_0 vdd vss x_2[30] x_3[30] multi_finger_inv_12
  Xgate_3_31_0 vdd vss x_2[31] x_3[31] multi_finger_inv_12
  Xgate_3_32_0 vdd vss x_2[32] x_3[32] multi_finger_inv_12
  Xgate_3_33_0 vdd vss x_2[33] x_3[33] multi_finger_inv_12
  Xgate_3_34_0 vdd vss x_2[34] x_3[34] multi_finger_inv_12
  Xgate_3_35_0 vdd vss x_2[35] x_3[35] multi_finger_inv_12
  Xgate_3_36_0 vdd vss x_2[36] x_3[36] multi_finger_inv_12
  Xgate_3_37_0 vdd vss x_2[37] x_3[37] multi_finger_inv_12
  Xgate_3_38_0 vdd vss x_2[38] x_3[38] multi_finger_inv_12
  Xgate_3_39_0 vdd vss x_2[39] x_3[39] multi_finger_inv_12
  Xgate_3_40_0 vdd vss x_2[40] x_3[40] multi_finger_inv_12
  Xgate_3_41_0 vdd vss x_2[41] x_3[41] multi_finger_inv_12
  Xgate_3_42_0 vdd vss x_2[42] x_3[42] multi_finger_inv_12
  Xgate_3_43_0 vdd vss x_2[43] x_3[43] multi_finger_inv_12
  Xgate_3_44_0 vdd vss x_2[44] x_3[44] multi_finger_inv_12
  Xgate_3_45_0 vdd vss x_2[45] x_3[45] multi_finger_inv_12
  Xgate_3_46_0 vdd vss x_2[46] x_3[46] multi_finger_inv_12
  Xgate_3_47_0 vdd vss x_2[47] x_3[47] multi_finger_inv_12
  Xgate_3_48_0 vdd vss x_2[48] x_3[48] multi_finger_inv_12
  Xgate_3_49_0 vdd vss x_2[49] x_3[49] multi_finger_inv_12
  Xgate_3_50_0 vdd vss x_2[50] x_3[50] multi_finger_inv_12
  Xgate_3_51_0 vdd vss x_2[51] x_3[51] multi_finger_inv_12
  Xgate_3_52_0 vdd vss x_2[52] x_3[52] multi_finger_inv_12
  Xgate_3_53_0 vdd vss x_2[53] x_3[53] multi_finger_inv_12
  Xgate_3_54_0 vdd vss x_2[54] x_3[54] multi_finger_inv_12
  Xgate_3_55_0 vdd vss x_2[55] x_3[55] multi_finger_inv_12
  Xgate_3_56_0 vdd vss x_2[56] x_3[56] multi_finger_inv_12
  Xgate_3_57_0 vdd vss x_2[57] x_3[57] multi_finger_inv_12
  Xgate_3_58_0 vdd vss x_2[58] x_3[58] multi_finger_inv_12
  Xgate_3_59_0 vdd vss x_2[59] x_3[59] multi_finger_inv_12
  Xgate_3_60_0 vdd vss x_2[60] x_3[60] multi_finger_inv_12
  Xgate_3_61_0 vdd vss x_2[61] x_3[61] multi_finger_inv_12
  Xgate_3_62_0 vdd vss x_2[62] x_3[62] multi_finger_inv_12
  Xgate_3_63_0 vdd vss x_2[63] x_3[63] multi_finger_inv_12
  Xgate_3_64_0 vdd vss x_2[64] x_3[64] multi_finger_inv_12
  Xgate_3_65_0 vdd vss x_2[65] x_3[65] multi_finger_inv_12
  Xgate_3_66_0 vdd vss x_2[66] x_3[66] multi_finger_inv_12
  Xgate_3_67_0 vdd vss x_2[67] x_3[67] multi_finger_inv_12
  Xgate_3_68_0 vdd vss x_2[68] x_3[68] multi_finger_inv_12
  Xgate_3_69_0 vdd vss x_2[69] x_3[69] multi_finger_inv_12
  Xgate_3_70_0 vdd vss x_2[70] x_3[70] multi_finger_inv_12
  Xgate_3_71_0 vdd vss x_2[71] x_3[71] multi_finger_inv_12
  Xgate_3_72_0 vdd vss x_2[72] x_3[72] multi_finger_inv_12
  Xgate_3_73_0 vdd vss x_2[73] x_3[73] multi_finger_inv_12
  Xgate_3_74_0 vdd vss x_2[74] x_3[74] multi_finger_inv_12
  Xgate_3_75_0 vdd vss x_2[75] x_3[75] multi_finger_inv_12
  Xgate_3_76_0 vdd vss x_2[76] x_3[76] multi_finger_inv_12
  Xgate_3_77_0 vdd vss x_2[77] x_3[77] multi_finger_inv_12
  Xgate_3_78_0 vdd vss x_2[78] x_3[78] multi_finger_inv_12
  Xgate_3_79_0 vdd vss x_2[79] x_3[79] multi_finger_inv_12
  Xgate_3_80_0 vdd vss x_2[80] x_3[80] multi_finger_inv_12
  Xgate_3_81_0 vdd vss x_2[81] x_3[81] multi_finger_inv_12
  Xgate_3_82_0 vdd vss x_2[82] x_3[82] multi_finger_inv_12
  Xgate_3_83_0 vdd vss x_2[83] x_3[83] multi_finger_inv_12
  Xgate_3_84_0 vdd vss x_2[84] x_3[84] multi_finger_inv_12
  Xgate_3_85_0 vdd vss x_2[85] x_3[85] multi_finger_inv_12
  Xgate_3_86_0 vdd vss x_2[86] x_3[86] multi_finger_inv_12
  Xgate_3_87_0 vdd vss x_2[87] x_3[87] multi_finger_inv_12
  Xgate_3_88_0 vdd vss x_2[88] x_3[88] multi_finger_inv_12
  Xgate_3_89_0 vdd vss x_2[89] x_3[89] multi_finger_inv_12
  Xgate_3_90_0 vdd vss x_2[90] x_3[90] multi_finger_inv_12
  Xgate_3_91_0 vdd vss x_2[91] x_3[91] multi_finger_inv_12
  Xgate_3_92_0 vdd vss x_2[92] x_3[92] multi_finger_inv_12
  Xgate_3_93_0 vdd vss x_2[93] x_3[93] multi_finger_inv_12
  Xgate_3_94_0 vdd vss x_2[94] x_3[94] multi_finger_inv_12
  Xgate_3_95_0 vdd vss x_2[95] x_3[95] multi_finger_inv_12
  Xgate_3_96_0 vdd vss x_2[96] x_3[96] multi_finger_inv_12
  Xgate_3_97_0 vdd vss x_2[97] x_3[97] multi_finger_inv_12
  Xgate_3_98_0 vdd vss x_2[98] x_3[98] multi_finger_inv_12
  Xgate_3_99_0 vdd vss x_2[99] x_3[99] multi_finger_inv_12
  Xgate_3_100_0 vdd vss x_2[100] x_3[100] multi_finger_inv_12
  Xgate_3_101_0 vdd vss x_2[101] x_3[101] multi_finger_inv_12
  Xgate_3_102_0 vdd vss x_2[102] x_3[102] multi_finger_inv_12
  Xgate_3_103_0 vdd vss x_2[103] x_3[103] multi_finger_inv_12
  Xgate_3_104_0 vdd vss x_2[104] x_3[104] multi_finger_inv_12
  Xgate_3_105_0 vdd vss x_2[105] x_3[105] multi_finger_inv_12
  Xgate_3_106_0 vdd vss x_2[106] x_3[106] multi_finger_inv_12
  Xgate_3_107_0 vdd vss x_2[107] x_3[107] multi_finger_inv_12
  Xgate_3_108_0 vdd vss x_2[108] x_3[108] multi_finger_inv_12
  Xgate_3_109_0 vdd vss x_2[109] x_3[109] multi_finger_inv_12
  Xgate_3_110_0 vdd vss x_2[110] x_3[110] multi_finger_inv_12
  Xgate_3_111_0 vdd vss x_2[111] x_3[111] multi_finger_inv_12
  Xgate_3_112_0 vdd vss x_2[112] x_3[112] multi_finger_inv_12
  Xgate_3_113_0 vdd vss x_2[113] x_3[113] multi_finger_inv_12
  Xgate_3_114_0 vdd vss x_2[114] x_3[114] multi_finger_inv_12
  Xgate_3_115_0 vdd vss x_2[115] x_3[115] multi_finger_inv_12
  Xgate_3_116_0 vdd vss x_2[116] x_3[116] multi_finger_inv_12
  Xgate_3_117_0 vdd vss x_2[117] x_3[117] multi_finger_inv_12
  Xgate_3_118_0 vdd vss x_2[118] x_3[118] multi_finger_inv_12
  Xgate_3_119_0 vdd vss x_2[119] x_3[119] multi_finger_inv_12
  Xgate_3_120_0 vdd vss x_2[120] x_3[120] multi_finger_inv_12
  Xgate_3_121_0 vdd vss x_2[121] x_3[121] multi_finger_inv_12
  Xgate_3_122_0 vdd vss x_2[122] x_3[122] multi_finger_inv_12
  Xgate_3_123_0 vdd vss x_2[123] x_3[123] multi_finger_inv_12
  Xgate_3_124_0 vdd vss x_2[124] x_3[124] multi_finger_inv_12
  Xgate_3_125_0 vdd vss x_2[125] x_3[125] multi_finger_inv_12
  Xgate_3_126_0 vdd vss x_2[126] x_3[126] multi_finger_inv_12
  Xgate_3_127_0 vdd vss x_2[127] x_3[127] multi_finger_inv_12
  Xgate_4_0_0 vdd vss x_3[0] x_4[0] multi_finger_inv_13
  Xgate_4_1_0 vdd vss x_3[1] x_4[1] multi_finger_inv_13
  Xgate_4_2_0 vdd vss x_3[2] x_4[2] multi_finger_inv_13
  Xgate_4_3_0 vdd vss x_3[3] x_4[3] multi_finger_inv_13
  Xgate_4_4_0 vdd vss x_3[4] x_4[4] multi_finger_inv_13
  Xgate_4_5_0 vdd vss x_3[5] x_4[5] multi_finger_inv_13
  Xgate_4_6_0 vdd vss x_3[6] x_4[6] multi_finger_inv_13
  Xgate_4_7_0 vdd vss x_3[7] x_4[7] multi_finger_inv_13
  Xgate_4_8_0 vdd vss x_3[8] x_4[8] multi_finger_inv_13
  Xgate_4_9_0 vdd vss x_3[9] x_4[9] multi_finger_inv_13
  Xgate_4_10_0 vdd vss x_3[10] x_4[10] multi_finger_inv_13
  Xgate_4_11_0 vdd vss x_3[11] x_4[11] multi_finger_inv_13
  Xgate_4_12_0 vdd vss x_3[12] x_4[12] multi_finger_inv_13
  Xgate_4_13_0 vdd vss x_3[13] x_4[13] multi_finger_inv_13
  Xgate_4_14_0 vdd vss x_3[14] x_4[14] multi_finger_inv_13
  Xgate_4_15_0 vdd vss x_3[15] x_4[15] multi_finger_inv_13
  Xgate_4_16_0 vdd vss x_3[16] x_4[16] multi_finger_inv_13
  Xgate_4_17_0 vdd vss x_3[17] x_4[17] multi_finger_inv_13
  Xgate_4_18_0 vdd vss x_3[18] x_4[18] multi_finger_inv_13
  Xgate_4_19_0 vdd vss x_3[19] x_4[19] multi_finger_inv_13
  Xgate_4_20_0 vdd vss x_3[20] x_4[20] multi_finger_inv_13
  Xgate_4_21_0 vdd vss x_3[21] x_4[21] multi_finger_inv_13
  Xgate_4_22_0 vdd vss x_3[22] x_4[22] multi_finger_inv_13
  Xgate_4_23_0 vdd vss x_3[23] x_4[23] multi_finger_inv_13
  Xgate_4_24_0 vdd vss x_3[24] x_4[24] multi_finger_inv_13
  Xgate_4_25_0 vdd vss x_3[25] x_4[25] multi_finger_inv_13
  Xgate_4_26_0 vdd vss x_3[26] x_4[26] multi_finger_inv_13
  Xgate_4_27_0 vdd vss x_3[27] x_4[27] multi_finger_inv_13
  Xgate_4_28_0 vdd vss x_3[28] x_4[28] multi_finger_inv_13
  Xgate_4_29_0 vdd vss x_3[29] x_4[29] multi_finger_inv_13
  Xgate_4_30_0 vdd vss x_3[30] x_4[30] multi_finger_inv_13
  Xgate_4_31_0 vdd vss x_3[31] x_4[31] multi_finger_inv_13
  Xgate_4_32_0 vdd vss x_3[32] x_4[32] multi_finger_inv_13
  Xgate_4_33_0 vdd vss x_3[33] x_4[33] multi_finger_inv_13
  Xgate_4_34_0 vdd vss x_3[34] x_4[34] multi_finger_inv_13
  Xgate_4_35_0 vdd vss x_3[35] x_4[35] multi_finger_inv_13
  Xgate_4_36_0 vdd vss x_3[36] x_4[36] multi_finger_inv_13
  Xgate_4_37_0 vdd vss x_3[37] x_4[37] multi_finger_inv_13
  Xgate_4_38_0 vdd vss x_3[38] x_4[38] multi_finger_inv_13
  Xgate_4_39_0 vdd vss x_3[39] x_4[39] multi_finger_inv_13
  Xgate_4_40_0 vdd vss x_3[40] x_4[40] multi_finger_inv_13
  Xgate_4_41_0 vdd vss x_3[41] x_4[41] multi_finger_inv_13
  Xgate_4_42_0 vdd vss x_3[42] x_4[42] multi_finger_inv_13
  Xgate_4_43_0 vdd vss x_3[43] x_4[43] multi_finger_inv_13
  Xgate_4_44_0 vdd vss x_3[44] x_4[44] multi_finger_inv_13
  Xgate_4_45_0 vdd vss x_3[45] x_4[45] multi_finger_inv_13
  Xgate_4_46_0 vdd vss x_3[46] x_4[46] multi_finger_inv_13
  Xgate_4_47_0 vdd vss x_3[47] x_4[47] multi_finger_inv_13
  Xgate_4_48_0 vdd vss x_3[48] x_4[48] multi_finger_inv_13
  Xgate_4_49_0 vdd vss x_3[49] x_4[49] multi_finger_inv_13
  Xgate_4_50_0 vdd vss x_3[50] x_4[50] multi_finger_inv_13
  Xgate_4_51_0 vdd vss x_3[51] x_4[51] multi_finger_inv_13
  Xgate_4_52_0 vdd vss x_3[52] x_4[52] multi_finger_inv_13
  Xgate_4_53_0 vdd vss x_3[53] x_4[53] multi_finger_inv_13
  Xgate_4_54_0 vdd vss x_3[54] x_4[54] multi_finger_inv_13
  Xgate_4_55_0 vdd vss x_3[55] x_4[55] multi_finger_inv_13
  Xgate_4_56_0 vdd vss x_3[56] x_4[56] multi_finger_inv_13
  Xgate_4_57_0 vdd vss x_3[57] x_4[57] multi_finger_inv_13
  Xgate_4_58_0 vdd vss x_3[58] x_4[58] multi_finger_inv_13
  Xgate_4_59_0 vdd vss x_3[59] x_4[59] multi_finger_inv_13
  Xgate_4_60_0 vdd vss x_3[60] x_4[60] multi_finger_inv_13
  Xgate_4_61_0 vdd vss x_3[61] x_4[61] multi_finger_inv_13
  Xgate_4_62_0 vdd vss x_3[62] x_4[62] multi_finger_inv_13
  Xgate_4_63_0 vdd vss x_3[63] x_4[63] multi_finger_inv_13
  Xgate_4_64_0 vdd vss x_3[64] x_4[64] multi_finger_inv_13
  Xgate_4_65_0 vdd vss x_3[65] x_4[65] multi_finger_inv_13
  Xgate_4_66_0 vdd vss x_3[66] x_4[66] multi_finger_inv_13
  Xgate_4_67_0 vdd vss x_3[67] x_4[67] multi_finger_inv_13
  Xgate_4_68_0 vdd vss x_3[68] x_4[68] multi_finger_inv_13
  Xgate_4_69_0 vdd vss x_3[69] x_4[69] multi_finger_inv_13
  Xgate_4_70_0 vdd vss x_3[70] x_4[70] multi_finger_inv_13
  Xgate_4_71_0 vdd vss x_3[71] x_4[71] multi_finger_inv_13
  Xgate_4_72_0 vdd vss x_3[72] x_4[72] multi_finger_inv_13
  Xgate_4_73_0 vdd vss x_3[73] x_4[73] multi_finger_inv_13
  Xgate_4_74_0 vdd vss x_3[74] x_4[74] multi_finger_inv_13
  Xgate_4_75_0 vdd vss x_3[75] x_4[75] multi_finger_inv_13
  Xgate_4_76_0 vdd vss x_3[76] x_4[76] multi_finger_inv_13
  Xgate_4_77_0 vdd vss x_3[77] x_4[77] multi_finger_inv_13
  Xgate_4_78_0 vdd vss x_3[78] x_4[78] multi_finger_inv_13
  Xgate_4_79_0 vdd vss x_3[79] x_4[79] multi_finger_inv_13
  Xgate_4_80_0 vdd vss x_3[80] x_4[80] multi_finger_inv_13
  Xgate_4_81_0 vdd vss x_3[81] x_4[81] multi_finger_inv_13
  Xgate_4_82_0 vdd vss x_3[82] x_4[82] multi_finger_inv_13
  Xgate_4_83_0 vdd vss x_3[83] x_4[83] multi_finger_inv_13
  Xgate_4_84_0 vdd vss x_3[84] x_4[84] multi_finger_inv_13
  Xgate_4_85_0 vdd vss x_3[85] x_4[85] multi_finger_inv_13
  Xgate_4_86_0 vdd vss x_3[86] x_4[86] multi_finger_inv_13
  Xgate_4_87_0 vdd vss x_3[87] x_4[87] multi_finger_inv_13
  Xgate_4_88_0 vdd vss x_3[88] x_4[88] multi_finger_inv_13
  Xgate_4_89_0 vdd vss x_3[89] x_4[89] multi_finger_inv_13
  Xgate_4_90_0 vdd vss x_3[90] x_4[90] multi_finger_inv_13
  Xgate_4_91_0 vdd vss x_3[91] x_4[91] multi_finger_inv_13
  Xgate_4_92_0 vdd vss x_3[92] x_4[92] multi_finger_inv_13
  Xgate_4_93_0 vdd vss x_3[93] x_4[93] multi_finger_inv_13
  Xgate_4_94_0 vdd vss x_3[94] x_4[94] multi_finger_inv_13
  Xgate_4_95_0 vdd vss x_3[95] x_4[95] multi_finger_inv_13
  Xgate_4_96_0 vdd vss x_3[96] x_4[96] multi_finger_inv_13
  Xgate_4_97_0 vdd vss x_3[97] x_4[97] multi_finger_inv_13
  Xgate_4_98_0 vdd vss x_3[98] x_4[98] multi_finger_inv_13
  Xgate_4_99_0 vdd vss x_3[99] x_4[99] multi_finger_inv_13
  Xgate_4_100_0 vdd vss x_3[100] x_4[100] multi_finger_inv_13
  Xgate_4_101_0 vdd vss x_3[101] x_4[101] multi_finger_inv_13
  Xgate_4_102_0 vdd vss x_3[102] x_4[102] multi_finger_inv_13
  Xgate_4_103_0 vdd vss x_3[103] x_4[103] multi_finger_inv_13
  Xgate_4_104_0 vdd vss x_3[104] x_4[104] multi_finger_inv_13
  Xgate_4_105_0 vdd vss x_3[105] x_4[105] multi_finger_inv_13
  Xgate_4_106_0 vdd vss x_3[106] x_4[106] multi_finger_inv_13
  Xgate_4_107_0 vdd vss x_3[107] x_4[107] multi_finger_inv_13
  Xgate_4_108_0 vdd vss x_3[108] x_4[108] multi_finger_inv_13
  Xgate_4_109_0 vdd vss x_3[109] x_4[109] multi_finger_inv_13
  Xgate_4_110_0 vdd vss x_3[110] x_4[110] multi_finger_inv_13
  Xgate_4_111_0 vdd vss x_3[111] x_4[111] multi_finger_inv_13
  Xgate_4_112_0 vdd vss x_3[112] x_4[112] multi_finger_inv_13
  Xgate_4_113_0 vdd vss x_3[113] x_4[113] multi_finger_inv_13
  Xgate_4_114_0 vdd vss x_3[114] x_4[114] multi_finger_inv_13
  Xgate_4_115_0 vdd vss x_3[115] x_4[115] multi_finger_inv_13
  Xgate_4_116_0 vdd vss x_3[116] x_4[116] multi_finger_inv_13
  Xgate_4_117_0 vdd vss x_3[117] x_4[117] multi_finger_inv_13
  Xgate_4_118_0 vdd vss x_3[118] x_4[118] multi_finger_inv_13
  Xgate_4_119_0 vdd vss x_3[119] x_4[119] multi_finger_inv_13
  Xgate_4_120_0 vdd vss x_3[120] x_4[120] multi_finger_inv_13
  Xgate_4_121_0 vdd vss x_3[121] x_4[121] multi_finger_inv_13
  Xgate_4_122_0 vdd vss x_3[122] x_4[122] multi_finger_inv_13
  Xgate_4_123_0 vdd vss x_3[123] x_4[123] multi_finger_inv_13
  Xgate_4_124_0 vdd vss x_3[124] x_4[124] multi_finger_inv_13
  Xgate_4_125_0 vdd vss x_3[125] x_4[125] multi_finger_inv_13
  Xgate_4_126_0 vdd vss x_3[126] x_4[126] multi_finger_inv_13
  Xgate_4_127_0 vdd vss x_3[127] x_4[127] multi_finger_inv_13
  Xgate_5_0_0 vdd vss x_4[0] y_b[0] multi_finger_inv_14
  Xgate_5_1_0 vdd vss x_4[1] y_b[1] multi_finger_inv_14
  Xgate_5_2_0 vdd vss x_4[2] y_b[2] multi_finger_inv_14
  Xgate_5_3_0 vdd vss x_4[3] y_b[3] multi_finger_inv_14
  Xgate_5_4_0 vdd vss x_4[4] y_b[4] multi_finger_inv_14
  Xgate_5_5_0 vdd vss x_4[5] y_b[5] multi_finger_inv_14
  Xgate_5_6_0 vdd vss x_4[6] y_b[6] multi_finger_inv_14
  Xgate_5_7_0 vdd vss x_4[7] y_b[7] multi_finger_inv_14
  Xgate_5_8_0 vdd vss x_4[8] y_b[8] multi_finger_inv_14
  Xgate_5_9_0 vdd vss x_4[9] y_b[9] multi_finger_inv_14
  Xgate_5_10_0 vdd vss x_4[10] y_b[10] multi_finger_inv_14
  Xgate_5_11_0 vdd vss x_4[11] y_b[11] multi_finger_inv_14
  Xgate_5_12_0 vdd vss x_4[12] y_b[12] multi_finger_inv_14
  Xgate_5_13_0 vdd vss x_4[13] y_b[13] multi_finger_inv_14
  Xgate_5_14_0 vdd vss x_4[14] y_b[14] multi_finger_inv_14
  Xgate_5_15_0 vdd vss x_4[15] y_b[15] multi_finger_inv_14
  Xgate_5_16_0 vdd vss x_4[16] y_b[16] multi_finger_inv_14
  Xgate_5_17_0 vdd vss x_4[17] y_b[17] multi_finger_inv_14
  Xgate_5_18_0 vdd vss x_4[18] y_b[18] multi_finger_inv_14
  Xgate_5_19_0 vdd vss x_4[19] y_b[19] multi_finger_inv_14
  Xgate_5_20_0 vdd vss x_4[20] y_b[20] multi_finger_inv_14
  Xgate_5_21_0 vdd vss x_4[21] y_b[21] multi_finger_inv_14
  Xgate_5_22_0 vdd vss x_4[22] y_b[22] multi_finger_inv_14
  Xgate_5_23_0 vdd vss x_4[23] y_b[23] multi_finger_inv_14
  Xgate_5_24_0 vdd vss x_4[24] y_b[24] multi_finger_inv_14
  Xgate_5_25_0 vdd vss x_4[25] y_b[25] multi_finger_inv_14
  Xgate_5_26_0 vdd vss x_4[26] y_b[26] multi_finger_inv_14
  Xgate_5_27_0 vdd vss x_4[27] y_b[27] multi_finger_inv_14
  Xgate_5_28_0 vdd vss x_4[28] y_b[28] multi_finger_inv_14
  Xgate_5_29_0 vdd vss x_4[29] y_b[29] multi_finger_inv_14
  Xgate_5_30_0 vdd vss x_4[30] y_b[30] multi_finger_inv_14
  Xgate_5_31_0 vdd vss x_4[31] y_b[31] multi_finger_inv_14
  Xgate_5_32_0 vdd vss x_4[32] y_b[32] multi_finger_inv_14
  Xgate_5_33_0 vdd vss x_4[33] y_b[33] multi_finger_inv_14
  Xgate_5_34_0 vdd vss x_4[34] y_b[34] multi_finger_inv_14
  Xgate_5_35_0 vdd vss x_4[35] y_b[35] multi_finger_inv_14
  Xgate_5_36_0 vdd vss x_4[36] y_b[36] multi_finger_inv_14
  Xgate_5_37_0 vdd vss x_4[37] y_b[37] multi_finger_inv_14
  Xgate_5_38_0 vdd vss x_4[38] y_b[38] multi_finger_inv_14
  Xgate_5_39_0 vdd vss x_4[39] y_b[39] multi_finger_inv_14
  Xgate_5_40_0 vdd vss x_4[40] y_b[40] multi_finger_inv_14
  Xgate_5_41_0 vdd vss x_4[41] y_b[41] multi_finger_inv_14
  Xgate_5_42_0 vdd vss x_4[42] y_b[42] multi_finger_inv_14
  Xgate_5_43_0 vdd vss x_4[43] y_b[43] multi_finger_inv_14
  Xgate_5_44_0 vdd vss x_4[44] y_b[44] multi_finger_inv_14
  Xgate_5_45_0 vdd vss x_4[45] y_b[45] multi_finger_inv_14
  Xgate_5_46_0 vdd vss x_4[46] y_b[46] multi_finger_inv_14
  Xgate_5_47_0 vdd vss x_4[47] y_b[47] multi_finger_inv_14
  Xgate_5_48_0 vdd vss x_4[48] y_b[48] multi_finger_inv_14
  Xgate_5_49_0 vdd vss x_4[49] y_b[49] multi_finger_inv_14
  Xgate_5_50_0 vdd vss x_4[50] y_b[50] multi_finger_inv_14
  Xgate_5_51_0 vdd vss x_4[51] y_b[51] multi_finger_inv_14
  Xgate_5_52_0 vdd vss x_4[52] y_b[52] multi_finger_inv_14
  Xgate_5_53_0 vdd vss x_4[53] y_b[53] multi_finger_inv_14
  Xgate_5_54_0 vdd vss x_4[54] y_b[54] multi_finger_inv_14
  Xgate_5_55_0 vdd vss x_4[55] y_b[55] multi_finger_inv_14
  Xgate_5_56_0 vdd vss x_4[56] y_b[56] multi_finger_inv_14
  Xgate_5_57_0 vdd vss x_4[57] y_b[57] multi_finger_inv_14
  Xgate_5_58_0 vdd vss x_4[58] y_b[58] multi_finger_inv_14
  Xgate_5_59_0 vdd vss x_4[59] y_b[59] multi_finger_inv_14
  Xgate_5_60_0 vdd vss x_4[60] y_b[60] multi_finger_inv_14
  Xgate_5_61_0 vdd vss x_4[61] y_b[61] multi_finger_inv_14
  Xgate_5_62_0 vdd vss x_4[62] y_b[62] multi_finger_inv_14
  Xgate_5_63_0 vdd vss x_4[63] y_b[63] multi_finger_inv_14
  Xgate_5_64_0 vdd vss x_4[64] y_b[64] multi_finger_inv_14
  Xgate_5_65_0 vdd vss x_4[65] y_b[65] multi_finger_inv_14
  Xgate_5_66_0 vdd vss x_4[66] y_b[66] multi_finger_inv_14
  Xgate_5_67_0 vdd vss x_4[67] y_b[67] multi_finger_inv_14
  Xgate_5_68_0 vdd vss x_4[68] y_b[68] multi_finger_inv_14
  Xgate_5_69_0 vdd vss x_4[69] y_b[69] multi_finger_inv_14
  Xgate_5_70_0 vdd vss x_4[70] y_b[70] multi_finger_inv_14
  Xgate_5_71_0 vdd vss x_4[71] y_b[71] multi_finger_inv_14
  Xgate_5_72_0 vdd vss x_4[72] y_b[72] multi_finger_inv_14
  Xgate_5_73_0 vdd vss x_4[73] y_b[73] multi_finger_inv_14
  Xgate_5_74_0 vdd vss x_4[74] y_b[74] multi_finger_inv_14
  Xgate_5_75_0 vdd vss x_4[75] y_b[75] multi_finger_inv_14
  Xgate_5_76_0 vdd vss x_4[76] y_b[76] multi_finger_inv_14
  Xgate_5_77_0 vdd vss x_4[77] y_b[77] multi_finger_inv_14
  Xgate_5_78_0 vdd vss x_4[78] y_b[78] multi_finger_inv_14
  Xgate_5_79_0 vdd vss x_4[79] y_b[79] multi_finger_inv_14
  Xgate_5_80_0 vdd vss x_4[80] y_b[80] multi_finger_inv_14
  Xgate_5_81_0 vdd vss x_4[81] y_b[81] multi_finger_inv_14
  Xgate_5_82_0 vdd vss x_4[82] y_b[82] multi_finger_inv_14
  Xgate_5_83_0 vdd vss x_4[83] y_b[83] multi_finger_inv_14
  Xgate_5_84_0 vdd vss x_4[84] y_b[84] multi_finger_inv_14
  Xgate_5_85_0 vdd vss x_4[85] y_b[85] multi_finger_inv_14
  Xgate_5_86_0 vdd vss x_4[86] y_b[86] multi_finger_inv_14
  Xgate_5_87_0 vdd vss x_4[87] y_b[87] multi_finger_inv_14
  Xgate_5_88_0 vdd vss x_4[88] y_b[88] multi_finger_inv_14
  Xgate_5_89_0 vdd vss x_4[89] y_b[89] multi_finger_inv_14
  Xgate_5_90_0 vdd vss x_4[90] y_b[90] multi_finger_inv_14
  Xgate_5_91_0 vdd vss x_4[91] y_b[91] multi_finger_inv_14
  Xgate_5_92_0 vdd vss x_4[92] y_b[92] multi_finger_inv_14
  Xgate_5_93_0 vdd vss x_4[93] y_b[93] multi_finger_inv_14
  Xgate_5_94_0 vdd vss x_4[94] y_b[94] multi_finger_inv_14
  Xgate_5_95_0 vdd vss x_4[95] y_b[95] multi_finger_inv_14
  Xgate_5_96_0 vdd vss x_4[96] y_b[96] multi_finger_inv_14
  Xgate_5_97_0 vdd vss x_4[97] y_b[97] multi_finger_inv_14
  Xgate_5_98_0 vdd vss x_4[98] y_b[98] multi_finger_inv_14
  Xgate_5_99_0 vdd vss x_4[99] y_b[99] multi_finger_inv_14
  Xgate_5_100_0 vdd vss x_4[100] y_b[100] multi_finger_inv_14
  Xgate_5_101_0 vdd vss x_4[101] y_b[101] multi_finger_inv_14
  Xgate_5_102_0 vdd vss x_4[102] y_b[102] multi_finger_inv_14
  Xgate_5_103_0 vdd vss x_4[103] y_b[103] multi_finger_inv_14
  Xgate_5_104_0 vdd vss x_4[104] y_b[104] multi_finger_inv_14
  Xgate_5_105_0 vdd vss x_4[105] y_b[105] multi_finger_inv_14
  Xgate_5_106_0 vdd vss x_4[106] y_b[106] multi_finger_inv_14
  Xgate_5_107_0 vdd vss x_4[107] y_b[107] multi_finger_inv_14
  Xgate_5_108_0 vdd vss x_4[108] y_b[108] multi_finger_inv_14
  Xgate_5_109_0 vdd vss x_4[109] y_b[109] multi_finger_inv_14
  Xgate_5_110_0 vdd vss x_4[110] y_b[110] multi_finger_inv_14
  Xgate_5_111_0 vdd vss x_4[111] y_b[111] multi_finger_inv_14
  Xgate_5_112_0 vdd vss x_4[112] y_b[112] multi_finger_inv_14
  Xgate_5_113_0 vdd vss x_4[113] y_b[113] multi_finger_inv_14
  Xgate_5_114_0 vdd vss x_4[114] y_b[114] multi_finger_inv_14
  Xgate_5_115_0 vdd vss x_4[115] y_b[115] multi_finger_inv_14
  Xgate_5_116_0 vdd vss x_4[116] y_b[116] multi_finger_inv_14
  Xgate_5_117_0 vdd vss x_4[117] y_b[117] multi_finger_inv_14
  Xgate_5_118_0 vdd vss x_4[118] y_b[118] multi_finger_inv_14
  Xgate_5_119_0 vdd vss x_4[119] y_b[119] multi_finger_inv_14
  Xgate_5_120_0 vdd vss x_4[120] y_b[120] multi_finger_inv_14
  Xgate_5_121_0 vdd vss x_4[121] y_b[121] multi_finger_inv_14
  Xgate_5_122_0 vdd vss x_4[122] y_b[122] multi_finger_inv_14
  Xgate_5_123_0 vdd vss x_4[123] y_b[123] multi_finger_inv_14
  Xgate_5_124_0 vdd vss x_4[124] y_b[124] multi_finger_inv_14
  Xgate_5_125_0 vdd vss x_4[125] y_b[125] multi_finger_inv_14
  Xgate_5_126_0 vdd vss x_4[126] y_b[126] multi_finger_inv_14
  Xgate_5_127_0 vdd vss x_4[127] y_b[127] multi_finger_inv_14
  Xgate_6_0_0 vdd vss y_b[0] y[0] multi_finger_inv_15
  Xgate_6_1_0 vdd vss y_b[1] y[1] multi_finger_inv_15
  Xgate_6_2_0 vdd vss y_b[2] y[2] multi_finger_inv_15
  Xgate_6_3_0 vdd vss y_b[3] y[3] multi_finger_inv_15
  Xgate_6_4_0 vdd vss y_b[4] y[4] multi_finger_inv_15
  Xgate_6_5_0 vdd vss y_b[5] y[5] multi_finger_inv_15
  Xgate_6_6_0 vdd vss y_b[6] y[6] multi_finger_inv_15
  Xgate_6_7_0 vdd vss y_b[7] y[7] multi_finger_inv_15
  Xgate_6_8_0 vdd vss y_b[8] y[8] multi_finger_inv_15
  Xgate_6_9_0 vdd vss y_b[9] y[9] multi_finger_inv_15
  Xgate_6_10_0 vdd vss y_b[10] y[10] multi_finger_inv_15
  Xgate_6_11_0 vdd vss y_b[11] y[11] multi_finger_inv_15
  Xgate_6_12_0 vdd vss y_b[12] y[12] multi_finger_inv_15
  Xgate_6_13_0 vdd vss y_b[13] y[13] multi_finger_inv_15
  Xgate_6_14_0 vdd vss y_b[14] y[14] multi_finger_inv_15
  Xgate_6_15_0 vdd vss y_b[15] y[15] multi_finger_inv_15
  Xgate_6_16_0 vdd vss y_b[16] y[16] multi_finger_inv_15
  Xgate_6_17_0 vdd vss y_b[17] y[17] multi_finger_inv_15
  Xgate_6_18_0 vdd vss y_b[18] y[18] multi_finger_inv_15
  Xgate_6_19_0 vdd vss y_b[19] y[19] multi_finger_inv_15
  Xgate_6_20_0 vdd vss y_b[20] y[20] multi_finger_inv_15
  Xgate_6_21_0 vdd vss y_b[21] y[21] multi_finger_inv_15
  Xgate_6_22_0 vdd vss y_b[22] y[22] multi_finger_inv_15
  Xgate_6_23_0 vdd vss y_b[23] y[23] multi_finger_inv_15
  Xgate_6_24_0 vdd vss y_b[24] y[24] multi_finger_inv_15
  Xgate_6_25_0 vdd vss y_b[25] y[25] multi_finger_inv_15
  Xgate_6_26_0 vdd vss y_b[26] y[26] multi_finger_inv_15
  Xgate_6_27_0 vdd vss y_b[27] y[27] multi_finger_inv_15
  Xgate_6_28_0 vdd vss y_b[28] y[28] multi_finger_inv_15
  Xgate_6_29_0 vdd vss y_b[29] y[29] multi_finger_inv_15
  Xgate_6_30_0 vdd vss y_b[30] y[30] multi_finger_inv_15
  Xgate_6_31_0 vdd vss y_b[31] y[31] multi_finger_inv_15
  Xgate_6_32_0 vdd vss y_b[32] y[32] multi_finger_inv_15
  Xgate_6_33_0 vdd vss y_b[33] y[33] multi_finger_inv_15
  Xgate_6_34_0 vdd vss y_b[34] y[34] multi_finger_inv_15
  Xgate_6_35_0 vdd vss y_b[35] y[35] multi_finger_inv_15
  Xgate_6_36_0 vdd vss y_b[36] y[36] multi_finger_inv_15
  Xgate_6_37_0 vdd vss y_b[37] y[37] multi_finger_inv_15
  Xgate_6_38_0 vdd vss y_b[38] y[38] multi_finger_inv_15
  Xgate_6_39_0 vdd vss y_b[39] y[39] multi_finger_inv_15
  Xgate_6_40_0 vdd vss y_b[40] y[40] multi_finger_inv_15
  Xgate_6_41_0 vdd vss y_b[41] y[41] multi_finger_inv_15
  Xgate_6_42_0 vdd vss y_b[42] y[42] multi_finger_inv_15
  Xgate_6_43_0 vdd vss y_b[43] y[43] multi_finger_inv_15
  Xgate_6_44_0 vdd vss y_b[44] y[44] multi_finger_inv_15
  Xgate_6_45_0 vdd vss y_b[45] y[45] multi_finger_inv_15
  Xgate_6_46_0 vdd vss y_b[46] y[46] multi_finger_inv_15
  Xgate_6_47_0 vdd vss y_b[47] y[47] multi_finger_inv_15
  Xgate_6_48_0 vdd vss y_b[48] y[48] multi_finger_inv_15
  Xgate_6_49_0 vdd vss y_b[49] y[49] multi_finger_inv_15
  Xgate_6_50_0 vdd vss y_b[50] y[50] multi_finger_inv_15
  Xgate_6_51_0 vdd vss y_b[51] y[51] multi_finger_inv_15
  Xgate_6_52_0 vdd vss y_b[52] y[52] multi_finger_inv_15
  Xgate_6_53_0 vdd vss y_b[53] y[53] multi_finger_inv_15
  Xgate_6_54_0 vdd vss y_b[54] y[54] multi_finger_inv_15
  Xgate_6_55_0 vdd vss y_b[55] y[55] multi_finger_inv_15
  Xgate_6_56_0 vdd vss y_b[56] y[56] multi_finger_inv_15
  Xgate_6_57_0 vdd vss y_b[57] y[57] multi_finger_inv_15
  Xgate_6_58_0 vdd vss y_b[58] y[58] multi_finger_inv_15
  Xgate_6_59_0 vdd vss y_b[59] y[59] multi_finger_inv_15
  Xgate_6_60_0 vdd vss y_b[60] y[60] multi_finger_inv_15
  Xgate_6_61_0 vdd vss y_b[61] y[61] multi_finger_inv_15
  Xgate_6_62_0 vdd vss y_b[62] y[62] multi_finger_inv_15
  Xgate_6_63_0 vdd vss y_b[63] y[63] multi_finger_inv_15
  Xgate_6_64_0 vdd vss y_b[64] y[64] multi_finger_inv_15
  Xgate_6_65_0 vdd vss y_b[65] y[65] multi_finger_inv_15
  Xgate_6_66_0 vdd vss y_b[66] y[66] multi_finger_inv_15
  Xgate_6_67_0 vdd vss y_b[67] y[67] multi_finger_inv_15
  Xgate_6_68_0 vdd vss y_b[68] y[68] multi_finger_inv_15
  Xgate_6_69_0 vdd vss y_b[69] y[69] multi_finger_inv_15
  Xgate_6_70_0 vdd vss y_b[70] y[70] multi_finger_inv_15
  Xgate_6_71_0 vdd vss y_b[71] y[71] multi_finger_inv_15
  Xgate_6_72_0 vdd vss y_b[72] y[72] multi_finger_inv_15
  Xgate_6_73_0 vdd vss y_b[73] y[73] multi_finger_inv_15
  Xgate_6_74_0 vdd vss y_b[74] y[74] multi_finger_inv_15
  Xgate_6_75_0 vdd vss y_b[75] y[75] multi_finger_inv_15
  Xgate_6_76_0 vdd vss y_b[76] y[76] multi_finger_inv_15
  Xgate_6_77_0 vdd vss y_b[77] y[77] multi_finger_inv_15
  Xgate_6_78_0 vdd vss y_b[78] y[78] multi_finger_inv_15
  Xgate_6_79_0 vdd vss y_b[79] y[79] multi_finger_inv_15
  Xgate_6_80_0 vdd vss y_b[80] y[80] multi_finger_inv_15
  Xgate_6_81_0 vdd vss y_b[81] y[81] multi_finger_inv_15
  Xgate_6_82_0 vdd vss y_b[82] y[82] multi_finger_inv_15
  Xgate_6_83_0 vdd vss y_b[83] y[83] multi_finger_inv_15
  Xgate_6_84_0 vdd vss y_b[84] y[84] multi_finger_inv_15
  Xgate_6_85_0 vdd vss y_b[85] y[85] multi_finger_inv_15
  Xgate_6_86_0 vdd vss y_b[86] y[86] multi_finger_inv_15
  Xgate_6_87_0 vdd vss y_b[87] y[87] multi_finger_inv_15
  Xgate_6_88_0 vdd vss y_b[88] y[88] multi_finger_inv_15
  Xgate_6_89_0 vdd vss y_b[89] y[89] multi_finger_inv_15
  Xgate_6_90_0 vdd vss y_b[90] y[90] multi_finger_inv_15
  Xgate_6_91_0 vdd vss y_b[91] y[91] multi_finger_inv_15
  Xgate_6_92_0 vdd vss y_b[92] y[92] multi_finger_inv_15
  Xgate_6_93_0 vdd vss y_b[93] y[93] multi_finger_inv_15
  Xgate_6_94_0 vdd vss y_b[94] y[94] multi_finger_inv_15
  Xgate_6_95_0 vdd vss y_b[95] y[95] multi_finger_inv_15
  Xgate_6_96_0 vdd vss y_b[96] y[96] multi_finger_inv_15
  Xgate_6_97_0 vdd vss y_b[97] y[97] multi_finger_inv_15
  Xgate_6_98_0 vdd vss y_b[98] y[98] multi_finger_inv_15
  Xgate_6_99_0 vdd vss y_b[99] y[99] multi_finger_inv_15
  Xgate_6_100_0 vdd vss y_b[100] y[100] multi_finger_inv_15
  Xgate_6_101_0 vdd vss y_b[101] y[101] multi_finger_inv_15
  Xgate_6_102_0 vdd vss y_b[102] y[102] multi_finger_inv_15
  Xgate_6_103_0 vdd vss y_b[103] y[103] multi_finger_inv_15
  Xgate_6_104_0 vdd vss y_b[104] y[104] multi_finger_inv_15
  Xgate_6_105_0 vdd vss y_b[105] y[105] multi_finger_inv_15
  Xgate_6_106_0 vdd vss y_b[106] y[106] multi_finger_inv_15
  Xgate_6_107_0 vdd vss y_b[107] y[107] multi_finger_inv_15
  Xgate_6_108_0 vdd vss y_b[108] y[108] multi_finger_inv_15
  Xgate_6_109_0 vdd vss y_b[109] y[109] multi_finger_inv_15
  Xgate_6_110_0 vdd vss y_b[110] y[110] multi_finger_inv_15
  Xgate_6_111_0 vdd vss y_b[111] y[111] multi_finger_inv_15
  Xgate_6_112_0 vdd vss y_b[112] y[112] multi_finger_inv_15
  Xgate_6_113_0 vdd vss y_b[113] y[113] multi_finger_inv_15
  Xgate_6_114_0 vdd vss y_b[114] y[114] multi_finger_inv_15
  Xgate_6_115_0 vdd vss y_b[115] y[115] multi_finger_inv_15
  Xgate_6_116_0 vdd vss y_b[116] y[116] multi_finger_inv_15
  Xgate_6_117_0 vdd vss y_b[117] y[117] multi_finger_inv_15
  Xgate_6_118_0 vdd vss y_b[118] y[118] multi_finger_inv_15
  Xgate_6_119_0 vdd vss y_b[119] y[119] multi_finger_inv_15
  Xgate_6_120_0 vdd vss y_b[120] y[120] multi_finger_inv_15
  Xgate_6_121_0 vdd vss y_b[121] y[121] multi_finger_inv_15
  Xgate_6_122_0 vdd vss y_b[122] y[122] multi_finger_inv_15
  Xgate_6_123_0 vdd vss y_b[123] y[123] multi_finger_inv_15
  Xgate_6_124_0 vdd vss y_b[124] y[124] multi_finger_inv_15
  Xgate_6_125_0 vdd vss y_b[125] y[125] multi_finger_inv_15
  Xgate_6_126_0 vdd vss y_b[126] y[126] multi_finger_inv_15
  Xgate_6_127_0 vdd vss y_b[127] y[127] multi_finger_inv_15

.ENDS decoder_stage_5

.SUBCKT nand2_1 vdd vss a b y

  Xn1 x a vss vss mos_w2000_l150_m1_nf1_id0
  Xn2 y b x vss mos_w2000_l150_m1_nf1_id0
  Xp1 y a vdd vdd mos_w2500_l150_m1_nf1_id1
  Xp2 y b vdd vdd mos_w2500_l150_m1_nf1_id1

.ENDS nand2_1

.SUBCKT multi_finger_inv_16 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_16

.SUBCKT multi_finger_inv_17 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_17

.SUBCKT multi_finger_inv_18 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_18

.SUBCKT multi_finger_inv_19 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP19 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP20 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP21 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP22 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP23 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP24 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP25 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP26 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP27 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN7 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN8 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN9 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN10 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_19

.SUBCKT multi_finger_inv_20 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP19 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP20 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP21 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP22 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP23 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP24 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP25 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP26 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP27 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP28 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP29 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP30 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP31 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP32 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP33 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP34 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP35 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP36 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP37 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP38 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP39 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP40 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP41 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP42 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP43 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP44 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP45 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP46 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP47 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP48 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP49 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP50 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP51 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP52 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP53 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP54 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP55 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP56 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP57 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP58 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP59 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP60 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP61 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP62 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP63 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP64 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP65 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP66 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP67 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP68 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP69 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP70 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP71 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP72 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP73 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN7 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN8 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN9 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN10 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN11 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN12 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN13 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN14 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN15 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN16 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN17 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN18 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN19 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN20 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN21 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN22 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN23 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN24 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN25 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN26 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN27 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN28 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_20

.SUBCKT decoder_stage_6 vdd vss y[0] y[1] y[2] y[3] y_b[0] y_b[1] y_b[2] y_b[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1

  Xgate_0_0_0 vdd vss predecode_0_0 predecode_1_0 x_0[0] nand2_1
  Xgate_0_1_0 vdd vss predecode_0_1 predecode_1_0 x_0[1] nand2_1
  Xgate_0_2_0 vdd vss predecode_0_0 predecode_1_1 x_0[2] nand2_1
  Xgate_0_3_0 vdd vss predecode_0_1 predecode_1_1 x_0[3] nand2_1
  Xgate_1_0_0 vdd vss x_0[0] x_1[0] multi_finger_inv_16
  Xgate_1_1_0 vdd vss x_0[1] x_1[1] multi_finger_inv_16
  Xgate_1_2_0 vdd vss x_0[2] x_1[2] multi_finger_inv_16
  Xgate_1_3_0 vdd vss x_0[3] x_1[3] multi_finger_inv_16
  Xgate_2_0_0 vdd vss x_1[0] x_2[0] multi_finger_inv_17
  Xgate_2_0_1 vdd vss x_1[0] x_2[0] multi_finger_inv_17
  Xgate_2_0_2 vdd vss x_1[0] x_2[0] multi_finger_inv_17
  Xgate_2_1_0 vdd vss x_1[1] x_2[1] multi_finger_inv_17
  Xgate_2_1_1 vdd vss x_1[1] x_2[1] multi_finger_inv_17
  Xgate_2_1_2 vdd vss x_1[1] x_2[1] multi_finger_inv_17
  Xgate_2_2_0 vdd vss x_1[2] x_2[2] multi_finger_inv_17
  Xgate_2_2_1 vdd vss x_1[2] x_2[2] multi_finger_inv_17
  Xgate_2_2_2 vdd vss x_1[2] x_2[2] multi_finger_inv_17
  Xgate_2_3_0 vdd vss x_1[3] x_2[3] multi_finger_inv_17
  Xgate_2_3_1 vdd vss x_1[3] x_2[3] multi_finger_inv_17
  Xgate_2_3_2 vdd vss x_1[3] x_2[3] multi_finger_inv_17
  Xgate_3_0_0 vdd vss x_2[0] x_3[0] multi_finger_inv_18
  Xgate_3_0_1 vdd vss x_2[0] x_3[0] multi_finger_inv_18
  Xgate_3_0_2 vdd vss x_2[0] x_3[0] multi_finger_inv_18
  Xgate_3_0_3 vdd vss x_2[0] x_3[0] multi_finger_inv_18
  Xgate_3_0_4 vdd vss x_2[0] x_3[0] multi_finger_inv_18
  Xgate_3_0_5 vdd vss x_2[0] x_3[0] multi_finger_inv_18
  Xgate_3_1_0 vdd vss x_2[1] x_3[1] multi_finger_inv_18
  Xgate_3_1_1 vdd vss x_2[1] x_3[1] multi_finger_inv_18
  Xgate_3_1_2 vdd vss x_2[1] x_3[1] multi_finger_inv_18
  Xgate_3_1_3 vdd vss x_2[1] x_3[1] multi_finger_inv_18
  Xgate_3_1_4 vdd vss x_2[1] x_3[1] multi_finger_inv_18
  Xgate_3_1_5 vdd vss x_2[1] x_3[1] multi_finger_inv_18
  Xgate_3_2_0 vdd vss x_2[2] x_3[2] multi_finger_inv_18
  Xgate_3_2_1 vdd vss x_2[2] x_3[2] multi_finger_inv_18
  Xgate_3_2_2 vdd vss x_2[2] x_3[2] multi_finger_inv_18
  Xgate_3_2_3 vdd vss x_2[2] x_3[2] multi_finger_inv_18
  Xgate_3_2_4 vdd vss x_2[2] x_3[2] multi_finger_inv_18
  Xgate_3_2_5 vdd vss x_2[2] x_3[2] multi_finger_inv_18
  Xgate_3_3_0 vdd vss x_2[3] x_3[3] multi_finger_inv_18
  Xgate_3_3_1 vdd vss x_2[3] x_3[3] multi_finger_inv_18
  Xgate_3_3_2 vdd vss x_2[3] x_3[3] multi_finger_inv_18
  Xgate_3_3_3 vdd vss x_2[3] x_3[3] multi_finger_inv_18
  Xgate_3_3_4 vdd vss x_2[3] x_3[3] multi_finger_inv_18
  Xgate_3_3_5 vdd vss x_2[3] x_3[3] multi_finger_inv_18
  Xgate_4_0_0 vdd vss x_3[0] y_b[0] multi_finger_inv_19
  Xgate_4_0_1 vdd vss x_3[0] y_b[0] multi_finger_inv_19
  Xgate_4_0_2 vdd vss x_3[0] y_b[0] multi_finger_inv_19
  Xgate_4_0_3 vdd vss x_3[0] y_b[0] multi_finger_inv_19
  Xgate_4_0_4 vdd vss x_3[0] y_b[0] multi_finger_inv_19
  Xgate_4_0_5 vdd vss x_3[0] y_b[0] multi_finger_inv_19
  Xgate_4_1_0 vdd vss x_3[1] y_b[1] multi_finger_inv_19
  Xgate_4_1_1 vdd vss x_3[1] y_b[1] multi_finger_inv_19
  Xgate_4_1_2 vdd vss x_3[1] y_b[1] multi_finger_inv_19
  Xgate_4_1_3 vdd vss x_3[1] y_b[1] multi_finger_inv_19
  Xgate_4_1_4 vdd vss x_3[1] y_b[1] multi_finger_inv_19
  Xgate_4_1_5 vdd vss x_3[1] y_b[1] multi_finger_inv_19
  Xgate_4_2_0 vdd vss x_3[2] y_b[2] multi_finger_inv_19
  Xgate_4_2_1 vdd vss x_3[2] y_b[2] multi_finger_inv_19
  Xgate_4_2_2 vdd vss x_3[2] y_b[2] multi_finger_inv_19
  Xgate_4_2_3 vdd vss x_3[2] y_b[2] multi_finger_inv_19
  Xgate_4_2_4 vdd vss x_3[2] y_b[2] multi_finger_inv_19
  Xgate_4_2_5 vdd vss x_3[2] y_b[2] multi_finger_inv_19
  Xgate_4_3_0 vdd vss x_3[3] y_b[3] multi_finger_inv_19
  Xgate_4_3_1 vdd vss x_3[3] y_b[3] multi_finger_inv_19
  Xgate_4_3_2 vdd vss x_3[3] y_b[3] multi_finger_inv_19
  Xgate_4_3_3 vdd vss x_3[3] y_b[3] multi_finger_inv_19
  Xgate_4_3_4 vdd vss x_3[3] y_b[3] multi_finger_inv_19
  Xgate_4_3_5 vdd vss x_3[3] y_b[3] multi_finger_inv_19
  Xgate_5_0_0 vdd vss y_b[0] y[0] multi_finger_inv_20
  Xgate_5_0_1 vdd vss y_b[0] y[0] multi_finger_inv_20
  Xgate_5_0_2 vdd vss y_b[0] y[0] multi_finger_inv_20
  Xgate_5_0_3 vdd vss y_b[0] y[0] multi_finger_inv_20
  Xgate_5_0_4 vdd vss y_b[0] y[0] multi_finger_inv_20
  Xgate_5_0_5 vdd vss y_b[0] y[0] multi_finger_inv_20
  Xgate_5_1_0 vdd vss y_b[1] y[1] multi_finger_inv_20
  Xgate_5_1_1 vdd vss y_b[1] y[1] multi_finger_inv_20
  Xgate_5_1_2 vdd vss y_b[1] y[1] multi_finger_inv_20
  Xgate_5_1_3 vdd vss y_b[1] y[1] multi_finger_inv_20
  Xgate_5_1_4 vdd vss y_b[1] y[1] multi_finger_inv_20
  Xgate_5_1_5 vdd vss y_b[1] y[1] multi_finger_inv_20
  Xgate_5_2_0 vdd vss y_b[2] y[2] multi_finger_inv_20
  Xgate_5_2_1 vdd vss y_b[2] y[2] multi_finger_inv_20
  Xgate_5_2_2 vdd vss y_b[2] y[2] multi_finger_inv_20
  Xgate_5_2_3 vdd vss y_b[2] y[2] multi_finger_inv_20
  Xgate_5_2_4 vdd vss y_b[2] y[2] multi_finger_inv_20
  Xgate_5_2_5 vdd vss y_b[2] y[2] multi_finger_inv_20
  Xgate_5_3_0 vdd vss y_b[3] y[3] multi_finger_inv_20
  Xgate_5_3_1 vdd vss y_b[3] y[3] multi_finger_inv_20
  Xgate_5_3_2 vdd vss y_b[3] y[3] multi_finger_inv_20
  Xgate_5_3_3 vdd vss y_b[3] y[3] multi_finger_inv_20
  Xgate_5_3_4 vdd vss y_b[3] y[3] multi_finger_inv_20
  Xgate_5_3_5 vdd vss y_b[3] y[3] multi_finger_inv_20

.ENDS decoder_stage_6

.SUBCKT decoder_1 vdd vss y[0] y[1] y[2] y[3] y_b[0] y_b[1] y_b[2] y_b[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1

  X0 vdd vss y[0] y[1] y[2] y[3] y_b[0] y_b[1] y_b[2] y_b[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 decoder_stage_6

.ENDS decoder_1

.SUBCKT sram_sp_hstrap_wrapper BR VDD VSS BL VNB VPB

  X0 BR VDD VSS BL VNB VPB sram_sp_hstrap

.ENDS sram_sp_hstrap_wrapper

.SUBCKT sram_sp_cell BL BR VDD VSS WL VNB VPB

  X0 QB WL BR VNB sky130_fd_pr__special_nfet_pass l=0.150 nf=1 w=0.140

  X1 Q QB VSS VNB sky130_fd_pr__special_nfet_latch l=0.150 nf=1 w=0.210

  X2 BL WL Q VNB sky130_fd_pr__special_nfet_pass l=0.150 nf=1 w=0.140

  X3 Q WL Q VPB sky130_fd_pr__special_pfet_pass l=0.025 nf=1 w=0.140

  X4 QB WL QB VPB sky130_fd_pr__special_pfet_pass l=0.025 nf=1 w=0.140

  X5 VDD Q QB VPB sky130_fd_pr__special_pfet_pass l=0.150 nf=1 w=0.140

  X6 Q QB VDD VPB sky130_fd_pr__special_pfet_pass l=0.150 nf=1 w=0.140

  X7 VSS Q QB VNB sky130_fd_pr__special_nfet_latch l=0.150 nf=1 w=0.210


.ENDS sram_sp_cell

.SUBCKT sram_sp_cell_wrapper BL BR VDD VSS WL VNB VPB

  X0 BL BR VDD VSS WL VNB VPB sram_sp_cell

.ENDS sram_sp_cell_wrapper

.SUBCKT sram_sp_colend BR VDD VSS BL VNB VPB

  X0 BR VNB BR VNB sky130_fd_pr__special_nfet_pass l=0.140 nf=1 w=0.140


.ENDS sram_sp_colend

.SUBCKT sram_sp_colend_wrapper BR VDD VSS BL VNB VPB

  X0 BR VDD VSS BL VNB VPB sram_sp_colend

.ENDS sram_sp_colend_wrapper

.SUBCKT sram_sp_horiz_wlstrap_p2 VSS VNB

  X0 VSS VSS VSS VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.420


.ENDS sram_sp_horiz_wlstrap_p2

.SUBCKT sram_sp_horiz_wlstrap_p2_wrapper VSS VNB

  X0 VSS VNB sram_sp_horiz_wlstrap_p2

.ENDS sram_sp_horiz_wlstrap_p2_wrapper

.SUBCKT sp_cell_array vdd vss dummy_bl dummy_br bl[0] bl[1] bl[2] bl[3] bl[4] bl[5] bl[6] bl[7] bl[8] bl[9] bl[10] bl[11] bl[12] bl[13] bl[14] bl[15] bl[16] bl[17] bl[18] bl[19] bl[20] bl[21] bl[22] bl[23] bl[24] bl[25] bl[26] bl[27] bl[28] bl[29] bl[30] bl[31] bl[32] bl[33] bl[34] bl[35] bl[36] bl[37] bl[38] bl[39] bl[40] bl[41] bl[42] bl[43] bl[44] bl[45] bl[46] bl[47] bl[48] bl[49] bl[50] bl[51] bl[52] bl[53] bl[54] bl[55] bl[56] bl[57] bl[58] bl[59] bl[60] bl[61] bl[62] bl[63] bl[64] bl[65] bl[66] bl[67] bl[68] bl[69] bl[70] bl[71] bl[72] bl[73] bl[74] bl[75] bl[76] bl[77] bl[78] bl[79] bl[80] bl[81] bl[82] bl[83] bl[84] bl[85] bl[86] bl[87] bl[88] bl[89] bl[90] bl[91] bl[92] bl[93] bl[94] bl[95] bl[96] bl[97] bl[98] bl[99] bl[100] bl[101] bl[102] bl[103] bl[104] bl[105] bl[106] bl[107] bl[108] bl[109] bl[110] bl[111] bl[112] bl[113] bl[114] bl[115] bl[116] bl[117] bl[118] bl[119] bl[120] bl[121] bl[122] bl[123] bl[124] bl[125] bl[126] bl[127] bl[128] bl[129] bl[130] bl[131] bl[132] bl[133] bl[134] bl[135] bl[136] bl[137] bl[138] bl[139] bl[140] bl[141] bl[142] bl[143] bl[144] bl[145] bl[146] bl[147] bl[148] bl[149] bl[150] bl[151] bl[152] bl[153] bl[154] bl[155] bl[156] bl[157] bl[158] bl[159] bl[160] bl[161] bl[162] bl[163] bl[164] bl[165] bl[166] bl[167] bl[168] bl[169] bl[170] bl[171] bl[172] bl[173] bl[174] bl[175] bl[176] bl[177] bl[178] bl[179] bl[180] bl[181] bl[182] bl[183] bl[184] bl[185] bl[186] bl[187] bl[188] bl[189] bl[190] bl[191] bl[192] bl[193] bl[194] bl[195] bl[196] bl[197] bl[198] bl[199] bl[200] bl[201] bl[202] bl[203] bl[204] bl[205] bl[206] bl[207] bl[208] bl[209] bl[210] bl[211] bl[212] bl[213] bl[214] bl[215] bl[216] bl[217] bl[218] bl[219] bl[220] bl[221] bl[222] bl[223] bl[224] bl[225] bl[226] bl[227] bl[228] bl[229] bl[230] bl[231] bl[232] bl[233] bl[234] bl[235] bl[236] bl[237] bl[238] bl[239] bl[240] bl[241] bl[242] bl[243] bl[244] bl[245] bl[246] bl[247] bl[248] bl[249] bl[250] bl[251] bl[252] bl[253] bl[254] bl[255] br[0] br[1] br[2] br[3] br[4] br[5] br[6] br[7] br[8] br[9] br[10] br[11] br[12] br[13] br[14] br[15] br[16] br[17] br[18] br[19] br[20] br[21] br[22] br[23] br[24] br[25] br[26] br[27] br[28] br[29] br[30] br[31] br[32] br[33] br[34] br[35] br[36] br[37] br[38] br[39] br[40] br[41] br[42] br[43] br[44] br[45] br[46] br[47] br[48] br[49] br[50] br[51] br[52] br[53] br[54] br[55] br[56] br[57] br[58] br[59] br[60] br[61] br[62] br[63] br[64] br[65] br[66] br[67] br[68] br[69] br[70] br[71] br[72] br[73] br[74] br[75] br[76] br[77] br[78] br[79] br[80] br[81] br[82] br[83] br[84] br[85] br[86] br[87] br[88] br[89] br[90] br[91] br[92] br[93] br[94] br[95] br[96] br[97] br[98] br[99] br[100] br[101] br[102] br[103] br[104] br[105] br[106] br[107] br[108] br[109] br[110] br[111] br[112] br[113] br[114] br[115] br[116] br[117] br[118] br[119] br[120] br[121] br[122] br[123] br[124] br[125] br[126] br[127] br[128] br[129] br[130] br[131] br[132] br[133] br[134] br[135] br[136] br[137] br[138] br[139] br[140] br[141] br[142] br[143] br[144] br[145] br[146] br[147] br[148] br[149] br[150] br[151] br[152] br[153] br[154] br[155] br[156] br[157] br[158] br[159] br[160] br[161] br[162] br[163] br[164] br[165] br[166] br[167] br[168] br[169] br[170] br[171] br[172] br[173] br[174] br[175] br[176] br[177] br[178] br[179] br[180] br[181] br[182] br[183] br[184] br[185] br[186] br[187] br[188] br[189] br[190] br[191] br[192] br[193] br[194] br[195] br[196] br[197] br[198] br[199] br[200] br[201] br[202] br[203] br[204] br[205] br[206] br[207] br[208] br[209] br[210] br[211] br[212] br[213] br[214] br[215] br[216] br[217] br[218] br[219] br[220] br[221] br[222] br[223] br[224] br[225] br[226] br[227] br[228] br[229] br[230] br[231] br[232] br[233] br[234] br[235] br[236] br[237] br[238] br[239] br[240] br[241] br[242] br[243] br[244] br[245] br[246] br[247] br[248] br[249] br[250] br[251] br[252] br[253] br[254] br[255] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127]

  Xcell_0_0 bl[0] br[0] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_1 bl[1] br[1] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_2 bl[2] br[2] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_3 bl[3] br[3] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_4 bl[4] br[4] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_5 bl[5] br[5] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_6 bl[6] br[6] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_7 bl[7] br[7] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_8 bl[8] br[8] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_9 bl[9] br[9] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_10 bl[10] br[10] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_11 bl[11] br[11] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_12 bl[12] br[12] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_13 bl[13] br[13] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_14 bl[14] br[14] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_15 bl[15] br[15] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_16 bl[16] br[16] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_17 bl[17] br[17] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_18 bl[18] br[18] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_19 bl[19] br[19] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_20 bl[20] br[20] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_21 bl[21] br[21] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_22 bl[22] br[22] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_23 bl[23] br[23] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_24 bl[24] br[24] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_25 bl[25] br[25] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_26 bl[26] br[26] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_27 bl[27] br[27] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_28 bl[28] br[28] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_29 bl[29] br[29] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_30 bl[30] br[30] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_31 bl[31] br[31] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_32 bl[32] br[32] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_33 bl[33] br[33] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_34 bl[34] br[34] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_35 bl[35] br[35] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_36 bl[36] br[36] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_37 bl[37] br[37] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_38 bl[38] br[38] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_39 bl[39] br[39] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_40 bl[40] br[40] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_41 bl[41] br[41] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_42 bl[42] br[42] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_43 bl[43] br[43] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_44 bl[44] br[44] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_45 bl[45] br[45] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_46 bl[46] br[46] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_47 bl[47] br[47] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_48 bl[48] br[48] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_49 bl[49] br[49] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_50 bl[50] br[50] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_51 bl[51] br[51] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_52 bl[52] br[52] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_53 bl[53] br[53] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_54 bl[54] br[54] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_55 bl[55] br[55] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_56 bl[56] br[56] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_57 bl[57] br[57] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_58 bl[58] br[58] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_59 bl[59] br[59] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_60 bl[60] br[60] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_61 bl[61] br[61] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_62 bl[62] br[62] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_63 bl[63] br[63] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_64 bl[64] br[64] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_65 bl[65] br[65] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_66 bl[66] br[66] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_67 bl[67] br[67] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_68 bl[68] br[68] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_69 bl[69] br[69] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_70 bl[70] br[70] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_71 bl[71] br[71] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_72 bl[72] br[72] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_73 bl[73] br[73] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_74 bl[74] br[74] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_75 bl[75] br[75] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_76 bl[76] br[76] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_77 bl[77] br[77] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_78 bl[78] br[78] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_79 bl[79] br[79] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_80 bl[80] br[80] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_81 bl[81] br[81] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_82 bl[82] br[82] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_83 bl[83] br[83] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_84 bl[84] br[84] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_85 bl[85] br[85] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_86 bl[86] br[86] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_87 bl[87] br[87] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_88 bl[88] br[88] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_89 bl[89] br[89] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_90 bl[90] br[90] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_91 bl[91] br[91] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_92 bl[92] br[92] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_93 bl[93] br[93] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_94 bl[94] br[94] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_95 bl[95] br[95] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_96 bl[96] br[96] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_97 bl[97] br[97] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_98 bl[98] br[98] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_99 bl[99] br[99] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_100 bl[100] br[100] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_101 bl[101] br[101] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_102 bl[102] br[102] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_103 bl[103] br[103] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_104 bl[104] br[104] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_105 bl[105] br[105] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_106 bl[106] br[106] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_107 bl[107] br[107] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_108 bl[108] br[108] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_109 bl[109] br[109] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_110 bl[110] br[110] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_111 bl[111] br[111] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_112 bl[112] br[112] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_113 bl[113] br[113] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_114 bl[114] br[114] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_115 bl[115] br[115] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_116 bl[116] br[116] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_117 bl[117] br[117] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_118 bl[118] br[118] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_119 bl[119] br[119] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_120 bl[120] br[120] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_121 bl[121] br[121] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_122 bl[122] br[122] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_123 bl[123] br[123] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_124 bl[124] br[124] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_125 bl[125] br[125] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_126 bl[126] br[126] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_127 bl[127] br[127] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_128 bl[128] br[128] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_129 bl[129] br[129] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_130 bl[130] br[130] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_131 bl[131] br[131] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_132 bl[132] br[132] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_133 bl[133] br[133] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_134 bl[134] br[134] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_135 bl[135] br[135] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_136 bl[136] br[136] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_137 bl[137] br[137] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_138 bl[138] br[138] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_139 bl[139] br[139] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_140 bl[140] br[140] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_141 bl[141] br[141] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_142 bl[142] br[142] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_143 bl[143] br[143] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_144 bl[144] br[144] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_145 bl[145] br[145] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_146 bl[146] br[146] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_147 bl[147] br[147] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_148 bl[148] br[148] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_149 bl[149] br[149] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_150 bl[150] br[150] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_151 bl[151] br[151] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_152 bl[152] br[152] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_153 bl[153] br[153] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_154 bl[154] br[154] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_155 bl[155] br[155] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_156 bl[156] br[156] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_157 bl[157] br[157] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_158 bl[158] br[158] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_159 bl[159] br[159] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_160 bl[160] br[160] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_161 bl[161] br[161] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_162 bl[162] br[162] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_163 bl[163] br[163] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_164 bl[164] br[164] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_165 bl[165] br[165] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_166 bl[166] br[166] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_167 bl[167] br[167] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_168 bl[168] br[168] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_169 bl[169] br[169] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_170 bl[170] br[170] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_171 bl[171] br[171] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_172 bl[172] br[172] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_173 bl[173] br[173] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_174 bl[174] br[174] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_175 bl[175] br[175] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_176 bl[176] br[176] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_177 bl[177] br[177] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_178 bl[178] br[178] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_179 bl[179] br[179] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_180 bl[180] br[180] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_181 bl[181] br[181] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_182 bl[182] br[182] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_183 bl[183] br[183] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_184 bl[184] br[184] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_185 bl[185] br[185] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_186 bl[186] br[186] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_187 bl[187] br[187] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_188 bl[188] br[188] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_189 bl[189] br[189] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_190 bl[190] br[190] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_191 bl[191] br[191] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_192 bl[192] br[192] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_193 bl[193] br[193] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_194 bl[194] br[194] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_195 bl[195] br[195] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_196 bl[196] br[196] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_197 bl[197] br[197] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_198 bl[198] br[198] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_199 bl[199] br[199] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_200 bl[200] br[200] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_201 bl[201] br[201] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_202 bl[202] br[202] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_203 bl[203] br[203] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_204 bl[204] br[204] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_205 bl[205] br[205] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_206 bl[206] br[206] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_207 bl[207] br[207] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_208 bl[208] br[208] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_209 bl[209] br[209] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_210 bl[210] br[210] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_211 bl[211] br[211] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_212 bl[212] br[212] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_213 bl[213] br[213] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_214 bl[214] br[214] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_215 bl[215] br[215] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_216 bl[216] br[216] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_217 bl[217] br[217] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_218 bl[218] br[218] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_219 bl[219] br[219] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_220 bl[220] br[220] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_221 bl[221] br[221] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_222 bl[222] br[222] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_223 bl[223] br[223] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_224 bl[224] br[224] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_225 bl[225] br[225] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_226 bl[226] br[226] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_227 bl[227] br[227] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_228 bl[228] br[228] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_229 bl[229] br[229] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_230 bl[230] br[230] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_231 bl[231] br[231] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_232 bl[232] br[232] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_233 bl[233] br[233] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_234 bl[234] br[234] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_235 bl[235] br[235] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_236 bl[236] br[236] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_237 bl[237] br[237] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_238 bl[238] br[238] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_239 bl[239] br[239] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_240 bl[240] br[240] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_241 bl[241] br[241] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_242 bl[242] br[242] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_243 bl[243] br[243] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_244 bl[244] br[244] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_245 bl[245] br[245] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_246 bl[246] br[246] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_247 bl[247] br[247] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_248 bl[248] br[248] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_249 bl[249] br[249] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_250 bl[250] br[250] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_251 bl[251] br[251] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_252 bl[252] br[252] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_253 bl[253] br[253] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_254 bl[254] br[254] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_255 bl[255] br[255] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_1_0 bl[0] br[0] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_1 bl[1] br[1] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_2 bl[2] br[2] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_3 bl[3] br[3] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_4 bl[4] br[4] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_5 bl[5] br[5] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_6 bl[6] br[6] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_7 bl[7] br[7] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_8 bl[8] br[8] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_9 bl[9] br[9] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_10 bl[10] br[10] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_11 bl[11] br[11] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_12 bl[12] br[12] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_13 bl[13] br[13] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_14 bl[14] br[14] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_15 bl[15] br[15] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_16 bl[16] br[16] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_17 bl[17] br[17] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_18 bl[18] br[18] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_19 bl[19] br[19] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_20 bl[20] br[20] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_21 bl[21] br[21] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_22 bl[22] br[22] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_23 bl[23] br[23] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_24 bl[24] br[24] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_25 bl[25] br[25] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_26 bl[26] br[26] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_27 bl[27] br[27] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_28 bl[28] br[28] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_29 bl[29] br[29] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_30 bl[30] br[30] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_31 bl[31] br[31] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_32 bl[32] br[32] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_33 bl[33] br[33] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_34 bl[34] br[34] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_35 bl[35] br[35] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_36 bl[36] br[36] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_37 bl[37] br[37] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_38 bl[38] br[38] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_39 bl[39] br[39] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_40 bl[40] br[40] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_41 bl[41] br[41] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_42 bl[42] br[42] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_43 bl[43] br[43] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_44 bl[44] br[44] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_45 bl[45] br[45] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_46 bl[46] br[46] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_47 bl[47] br[47] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_48 bl[48] br[48] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_49 bl[49] br[49] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_50 bl[50] br[50] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_51 bl[51] br[51] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_52 bl[52] br[52] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_53 bl[53] br[53] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_54 bl[54] br[54] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_55 bl[55] br[55] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_56 bl[56] br[56] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_57 bl[57] br[57] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_58 bl[58] br[58] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_59 bl[59] br[59] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_60 bl[60] br[60] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_61 bl[61] br[61] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_62 bl[62] br[62] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_63 bl[63] br[63] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_64 bl[64] br[64] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_65 bl[65] br[65] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_66 bl[66] br[66] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_67 bl[67] br[67] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_68 bl[68] br[68] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_69 bl[69] br[69] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_70 bl[70] br[70] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_71 bl[71] br[71] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_72 bl[72] br[72] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_73 bl[73] br[73] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_74 bl[74] br[74] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_75 bl[75] br[75] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_76 bl[76] br[76] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_77 bl[77] br[77] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_78 bl[78] br[78] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_79 bl[79] br[79] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_80 bl[80] br[80] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_81 bl[81] br[81] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_82 bl[82] br[82] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_83 bl[83] br[83] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_84 bl[84] br[84] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_85 bl[85] br[85] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_86 bl[86] br[86] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_87 bl[87] br[87] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_88 bl[88] br[88] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_89 bl[89] br[89] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_90 bl[90] br[90] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_91 bl[91] br[91] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_92 bl[92] br[92] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_93 bl[93] br[93] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_94 bl[94] br[94] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_95 bl[95] br[95] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_96 bl[96] br[96] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_97 bl[97] br[97] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_98 bl[98] br[98] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_99 bl[99] br[99] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_100 bl[100] br[100] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_101 bl[101] br[101] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_102 bl[102] br[102] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_103 bl[103] br[103] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_104 bl[104] br[104] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_105 bl[105] br[105] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_106 bl[106] br[106] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_107 bl[107] br[107] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_108 bl[108] br[108] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_109 bl[109] br[109] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_110 bl[110] br[110] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_111 bl[111] br[111] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_112 bl[112] br[112] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_113 bl[113] br[113] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_114 bl[114] br[114] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_115 bl[115] br[115] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_116 bl[116] br[116] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_117 bl[117] br[117] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_118 bl[118] br[118] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_119 bl[119] br[119] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_120 bl[120] br[120] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_121 bl[121] br[121] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_122 bl[122] br[122] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_123 bl[123] br[123] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_124 bl[124] br[124] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_125 bl[125] br[125] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_126 bl[126] br[126] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_127 bl[127] br[127] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_128 bl[128] br[128] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_129 bl[129] br[129] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_130 bl[130] br[130] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_131 bl[131] br[131] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_132 bl[132] br[132] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_133 bl[133] br[133] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_134 bl[134] br[134] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_135 bl[135] br[135] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_136 bl[136] br[136] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_137 bl[137] br[137] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_138 bl[138] br[138] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_139 bl[139] br[139] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_140 bl[140] br[140] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_141 bl[141] br[141] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_142 bl[142] br[142] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_143 bl[143] br[143] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_144 bl[144] br[144] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_145 bl[145] br[145] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_146 bl[146] br[146] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_147 bl[147] br[147] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_148 bl[148] br[148] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_149 bl[149] br[149] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_150 bl[150] br[150] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_151 bl[151] br[151] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_152 bl[152] br[152] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_153 bl[153] br[153] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_154 bl[154] br[154] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_155 bl[155] br[155] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_156 bl[156] br[156] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_157 bl[157] br[157] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_158 bl[158] br[158] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_159 bl[159] br[159] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_160 bl[160] br[160] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_161 bl[161] br[161] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_162 bl[162] br[162] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_163 bl[163] br[163] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_164 bl[164] br[164] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_165 bl[165] br[165] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_166 bl[166] br[166] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_167 bl[167] br[167] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_168 bl[168] br[168] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_169 bl[169] br[169] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_170 bl[170] br[170] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_171 bl[171] br[171] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_172 bl[172] br[172] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_173 bl[173] br[173] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_174 bl[174] br[174] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_175 bl[175] br[175] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_176 bl[176] br[176] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_177 bl[177] br[177] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_178 bl[178] br[178] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_179 bl[179] br[179] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_180 bl[180] br[180] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_181 bl[181] br[181] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_182 bl[182] br[182] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_183 bl[183] br[183] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_184 bl[184] br[184] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_185 bl[185] br[185] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_186 bl[186] br[186] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_187 bl[187] br[187] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_188 bl[188] br[188] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_189 bl[189] br[189] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_190 bl[190] br[190] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_191 bl[191] br[191] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_192 bl[192] br[192] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_193 bl[193] br[193] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_194 bl[194] br[194] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_195 bl[195] br[195] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_196 bl[196] br[196] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_197 bl[197] br[197] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_198 bl[198] br[198] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_199 bl[199] br[199] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_200 bl[200] br[200] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_201 bl[201] br[201] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_202 bl[202] br[202] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_203 bl[203] br[203] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_204 bl[204] br[204] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_205 bl[205] br[205] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_206 bl[206] br[206] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_207 bl[207] br[207] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_208 bl[208] br[208] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_209 bl[209] br[209] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_210 bl[210] br[210] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_211 bl[211] br[211] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_212 bl[212] br[212] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_213 bl[213] br[213] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_214 bl[214] br[214] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_215 bl[215] br[215] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_216 bl[216] br[216] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_217 bl[217] br[217] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_218 bl[218] br[218] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_219 bl[219] br[219] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_220 bl[220] br[220] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_221 bl[221] br[221] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_222 bl[222] br[222] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_223 bl[223] br[223] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_224 bl[224] br[224] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_225 bl[225] br[225] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_226 bl[226] br[226] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_227 bl[227] br[227] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_228 bl[228] br[228] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_229 bl[229] br[229] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_230 bl[230] br[230] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_231 bl[231] br[231] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_232 bl[232] br[232] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_233 bl[233] br[233] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_234 bl[234] br[234] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_235 bl[235] br[235] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_236 bl[236] br[236] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_237 bl[237] br[237] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_238 bl[238] br[238] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_239 bl[239] br[239] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_240 bl[240] br[240] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_241 bl[241] br[241] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_242 bl[242] br[242] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_243 bl[243] br[243] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_244 bl[244] br[244] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_245 bl[245] br[245] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_246 bl[246] br[246] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_247 bl[247] br[247] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_248 bl[248] br[248] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_249 bl[249] br[249] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_250 bl[250] br[250] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_251 bl[251] br[251] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_252 bl[252] br[252] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_253 bl[253] br[253] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_254 bl[254] br[254] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_255 bl[255] br[255] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_2_0 bl[0] br[0] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_1 bl[1] br[1] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_2 bl[2] br[2] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_3 bl[3] br[3] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_4 bl[4] br[4] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_5 bl[5] br[5] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_6 bl[6] br[6] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_7 bl[7] br[7] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_8 bl[8] br[8] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_9 bl[9] br[9] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_10 bl[10] br[10] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_11 bl[11] br[11] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_12 bl[12] br[12] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_13 bl[13] br[13] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_14 bl[14] br[14] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_15 bl[15] br[15] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_16 bl[16] br[16] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_17 bl[17] br[17] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_18 bl[18] br[18] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_19 bl[19] br[19] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_20 bl[20] br[20] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_21 bl[21] br[21] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_22 bl[22] br[22] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_23 bl[23] br[23] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_24 bl[24] br[24] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_25 bl[25] br[25] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_26 bl[26] br[26] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_27 bl[27] br[27] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_28 bl[28] br[28] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_29 bl[29] br[29] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_30 bl[30] br[30] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_31 bl[31] br[31] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_32 bl[32] br[32] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_33 bl[33] br[33] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_34 bl[34] br[34] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_35 bl[35] br[35] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_36 bl[36] br[36] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_37 bl[37] br[37] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_38 bl[38] br[38] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_39 bl[39] br[39] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_40 bl[40] br[40] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_41 bl[41] br[41] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_42 bl[42] br[42] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_43 bl[43] br[43] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_44 bl[44] br[44] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_45 bl[45] br[45] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_46 bl[46] br[46] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_47 bl[47] br[47] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_48 bl[48] br[48] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_49 bl[49] br[49] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_50 bl[50] br[50] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_51 bl[51] br[51] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_52 bl[52] br[52] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_53 bl[53] br[53] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_54 bl[54] br[54] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_55 bl[55] br[55] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_56 bl[56] br[56] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_57 bl[57] br[57] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_58 bl[58] br[58] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_59 bl[59] br[59] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_60 bl[60] br[60] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_61 bl[61] br[61] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_62 bl[62] br[62] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_63 bl[63] br[63] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_64 bl[64] br[64] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_65 bl[65] br[65] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_66 bl[66] br[66] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_67 bl[67] br[67] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_68 bl[68] br[68] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_69 bl[69] br[69] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_70 bl[70] br[70] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_71 bl[71] br[71] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_72 bl[72] br[72] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_73 bl[73] br[73] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_74 bl[74] br[74] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_75 bl[75] br[75] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_76 bl[76] br[76] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_77 bl[77] br[77] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_78 bl[78] br[78] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_79 bl[79] br[79] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_80 bl[80] br[80] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_81 bl[81] br[81] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_82 bl[82] br[82] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_83 bl[83] br[83] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_84 bl[84] br[84] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_85 bl[85] br[85] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_86 bl[86] br[86] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_87 bl[87] br[87] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_88 bl[88] br[88] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_89 bl[89] br[89] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_90 bl[90] br[90] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_91 bl[91] br[91] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_92 bl[92] br[92] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_93 bl[93] br[93] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_94 bl[94] br[94] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_95 bl[95] br[95] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_96 bl[96] br[96] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_97 bl[97] br[97] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_98 bl[98] br[98] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_99 bl[99] br[99] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_100 bl[100] br[100] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_101 bl[101] br[101] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_102 bl[102] br[102] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_103 bl[103] br[103] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_104 bl[104] br[104] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_105 bl[105] br[105] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_106 bl[106] br[106] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_107 bl[107] br[107] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_108 bl[108] br[108] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_109 bl[109] br[109] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_110 bl[110] br[110] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_111 bl[111] br[111] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_112 bl[112] br[112] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_113 bl[113] br[113] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_114 bl[114] br[114] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_115 bl[115] br[115] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_116 bl[116] br[116] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_117 bl[117] br[117] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_118 bl[118] br[118] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_119 bl[119] br[119] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_120 bl[120] br[120] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_121 bl[121] br[121] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_122 bl[122] br[122] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_123 bl[123] br[123] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_124 bl[124] br[124] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_125 bl[125] br[125] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_126 bl[126] br[126] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_127 bl[127] br[127] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_128 bl[128] br[128] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_129 bl[129] br[129] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_130 bl[130] br[130] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_131 bl[131] br[131] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_132 bl[132] br[132] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_133 bl[133] br[133] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_134 bl[134] br[134] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_135 bl[135] br[135] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_136 bl[136] br[136] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_137 bl[137] br[137] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_138 bl[138] br[138] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_139 bl[139] br[139] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_140 bl[140] br[140] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_141 bl[141] br[141] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_142 bl[142] br[142] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_143 bl[143] br[143] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_144 bl[144] br[144] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_145 bl[145] br[145] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_146 bl[146] br[146] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_147 bl[147] br[147] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_148 bl[148] br[148] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_149 bl[149] br[149] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_150 bl[150] br[150] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_151 bl[151] br[151] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_152 bl[152] br[152] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_153 bl[153] br[153] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_154 bl[154] br[154] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_155 bl[155] br[155] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_156 bl[156] br[156] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_157 bl[157] br[157] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_158 bl[158] br[158] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_159 bl[159] br[159] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_160 bl[160] br[160] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_161 bl[161] br[161] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_162 bl[162] br[162] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_163 bl[163] br[163] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_164 bl[164] br[164] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_165 bl[165] br[165] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_166 bl[166] br[166] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_167 bl[167] br[167] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_168 bl[168] br[168] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_169 bl[169] br[169] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_170 bl[170] br[170] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_171 bl[171] br[171] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_172 bl[172] br[172] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_173 bl[173] br[173] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_174 bl[174] br[174] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_175 bl[175] br[175] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_176 bl[176] br[176] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_177 bl[177] br[177] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_178 bl[178] br[178] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_179 bl[179] br[179] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_180 bl[180] br[180] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_181 bl[181] br[181] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_182 bl[182] br[182] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_183 bl[183] br[183] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_184 bl[184] br[184] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_185 bl[185] br[185] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_186 bl[186] br[186] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_187 bl[187] br[187] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_188 bl[188] br[188] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_189 bl[189] br[189] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_190 bl[190] br[190] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_191 bl[191] br[191] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_192 bl[192] br[192] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_193 bl[193] br[193] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_194 bl[194] br[194] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_195 bl[195] br[195] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_196 bl[196] br[196] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_197 bl[197] br[197] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_198 bl[198] br[198] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_199 bl[199] br[199] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_200 bl[200] br[200] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_201 bl[201] br[201] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_202 bl[202] br[202] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_203 bl[203] br[203] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_204 bl[204] br[204] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_205 bl[205] br[205] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_206 bl[206] br[206] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_207 bl[207] br[207] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_208 bl[208] br[208] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_209 bl[209] br[209] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_210 bl[210] br[210] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_211 bl[211] br[211] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_212 bl[212] br[212] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_213 bl[213] br[213] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_214 bl[214] br[214] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_215 bl[215] br[215] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_216 bl[216] br[216] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_217 bl[217] br[217] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_218 bl[218] br[218] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_219 bl[219] br[219] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_220 bl[220] br[220] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_221 bl[221] br[221] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_222 bl[222] br[222] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_223 bl[223] br[223] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_224 bl[224] br[224] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_225 bl[225] br[225] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_226 bl[226] br[226] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_227 bl[227] br[227] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_228 bl[228] br[228] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_229 bl[229] br[229] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_230 bl[230] br[230] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_231 bl[231] br[231] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_232 bl[232] br[232] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_233 bl[233] br[233] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_234 bl[234] br[234] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_235 bl[235] br[235] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_236 bl[236] br[236] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_237 bl[237] br[237] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_238 bl[238] br[238] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_239 bl[239] br[239] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_240 bl[240] br[240] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_241 bl[241] br[241] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_242 bl[242] br[242] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_243 bl[243] br[243] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_244 bl[244] br[244] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_245 bl[245] br[245] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_246 bl[246] br[246] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_247 bl[247] br[247] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_248 bl[248] br[248] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_249 bl[249] br[249] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_250 bl[250] br[250] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_251 bl[251] br[251] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_252 bl[252] br[252] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_253 bl[253] br[253] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_254 bl[254] br[254] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_255 bl[255] br[255] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_3_0 bl[0] br[0] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_1 bl[1] br[1] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_2 bl[2] br[2] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_3 bl[3] br[3] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_4 bl[4] br[4] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_5 bl[5] br[5] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_6 bl[6] br[6] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_7 bl[7] br[7] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_8 bl[8] br[8] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_9 bl[9] br[9] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_10 bl[10] br[10] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_11 bl[11] br[11] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_12 bl[12] br[12] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_13 bl[13] br[13] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_14 bl[14] br[14] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_15 bl[15] br[15] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_16 bl[16] br[16] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_17 bl[17] br[17] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_18 bl[18] br[18] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_19 bl[19] br[19] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_20 bl[20] br[20] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_21 bl[21] br[21] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_22 bl[22] br[22] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_23 bl[23] br[23] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_24 bl[24] br[24] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_25 bl[25] br[25] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_26 bl[26] br[26] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_27 bl[27] br[27] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_28 bl[28] br[28] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_29 bl[29] br[29] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_30 bl[30] br[30] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_31 bl[31] br[31] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_32 bl[32] br[32] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_33 bl[33] br[33] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_34 bl[34] br[34] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_35 bl[35] br[35] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_36 bl[36] br[36] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_37 bl[37] br[37] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_38 bl[38] br[38] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_39 bl[39] br[39] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_40 bl[40] br[40] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_41 bl[41] br[41] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_42 bl[42] br[42] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_43 bl[43] br[43] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_44 bl[44] br[44] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_45 bl[45] br[45] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_46 bl[46] br[46] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_47 bl[47] br[47] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_48 bl[48] br[48] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_49 bl[49] br[49] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_50 bl[50] br[50] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_51 bl[51] br[51] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_52 bl[52] br[52] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_53 bl[53] br[53] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_54 bl[54] br[54] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_55 bl[55] br[55] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_56 bl[56] br[56] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_57 bl[57] br[57] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_58 bl[58] br[58] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_59 bl[59] br[59] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_60 bl[60] br[60] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_61 bl[61] br[61] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_62 bl[62] br[62] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_63 bl[63] br[63] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_64 bl[64] br[64] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_65 bl[65] br[65] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_66 bl[66] br[66] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_67 bl[67] br[67] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_68 bl[68] br[68] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_69 bl[69] br[69] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_70 bl[70] br[70] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_71 bl[71] br[71] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_72 bl[72] br[72] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_73 bl[73] br[73] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_74 bl[74] br[74] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_75 bl[75] br[75] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_76 bl[76] br[76] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_77 bl[77] br[77] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_78 bl[78] br[78] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_79 bl[79] br[79] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_80 bl[80] br[80] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_81 bl[81] br[81] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_82 bl[82] br[82] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_83 bl[83] br[83] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_84 bl[84] br[84] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_85 bl[85] br[85] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_86 bl[86] br[86] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_87 bl[87] br[87] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_88 bl[88] br[88] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_89 bl[89] br[89] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_90 bl[90] br[90] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_91 bl[91] br[91] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_92 bl[92] br[92] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_93 bl[93] br[93] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_94 bl[94] br[94] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_95 bl[95] br[95] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_96 bl[96] br[96] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_97 bl[97] br[97] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_98 bl[98] br[98] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_99 bl[99] br[99] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_100 bl[100] br[100] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_101 bl[101] br[101] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_102 bl[102] br[102] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_103 bl[103] br[103] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_104 bl[104] br[104] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_105 bl[105] br[105] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_106 bl[106] br[106] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_107 bl[107] br[107] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_108 bl[108] br[108] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_109 bl[109] br[109] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_110 bl[110] br[110] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_111 bl[111] br[111] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_112 bl[112] br[112] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_113 bl[113] br[113] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_114 bl[114] br[114] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_115 bl[115] br[115] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_116 bl[116] br[116] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_117 bl[117] br[117] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_118 bl[118] br[118] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_119 bl[119] br[119] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_120 bl[120] br[120] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_121 bl[121] br[121] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_122 bl[122] br[122] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_123 bl[123] br[123] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_124 bl[124] br[124] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_125 bl[125] br[125] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_126 bl[126] br[126] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_127 bl[127] br[127] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_128 bl[128] br[128] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_129 bl[129] br[129] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_130 bl[130] br[130] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_131 bl[131] br[131] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_132 bl[132] br[132] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_133 bl[133] br[133] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_134 bl[134] br[134] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_135 bl[135] br[135] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_136 bl[136] br[136] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_137 bl[137] br[137] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_138 bl[138] br[138] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_139 bl[139] br[139] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_140 bl[140] br[140] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_141 bl[141] br[141] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_142 bl[142] br[142] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_143 bl[143] br[143] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_144 bl[144] br[144] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_145 bl[145] br[145] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_146 bl[146] br[146] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_147 bl[147] br[147] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_148 bl[148] br[148] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_149 bl[149] br[149] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_150 bl[150] br[150] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_151 bl[151] br[151] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_152 bl[152] br[152] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_153 bl[153] br[153] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_154 bl[154] br[154] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_155 bl[155] br[155] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_156 bl[156] br[156] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_157 bl[157] br[157] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_158 bl[158] br[158] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_159 bl[159] br[159] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_160 bl[160] br[160] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_161 bl[161] br[161] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_162 bl[162] br[162] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_163 bl[163] br[163] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_164 bl[164] br[164] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_165 bl[165] br[165] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_166 bl[166] br[166] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_167 bl[167] br[167] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_168 bl[168] br[168] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_169 bl[169] br[169] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_170 bl[170] br[170] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_171 bl[171] br[171] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_172 bl[172] br[172] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_173 bl[173] br[173] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_174 bl[174] br[174] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_175 bl[175] br[175] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_176 bl[176] br[176] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_177 bl[177] br[177] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_178 bl[178] br[178] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_179 bl[179] br[179] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_180 bl[180] br[180] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_181 bl[181] br[181] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_182 bl[182] br[182] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_183 bl[183] br[183] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_184 bl[184] br[184] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_185 bl[185] br[185] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_186 bl[186] br[186] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_187 bl[187] br[187] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_188 bl[188] br[188] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_189 bl[189] br[189] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_190 bl[190] br[190] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_191 bl[191] br[191] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_192 bl[192] br[192] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_193 bl[193] br[193] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_194 bl[194] br[194] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_195 bl[195] br[195] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_196 bl[196] br[196] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_197 bl[197] br[197] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_198 bl[198] br[198] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_199 bl[199] br[199] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_200 bl[200] br[200] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_201 bl[201] br[201] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_202 bl[202] br[202] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_203 bl[203] br[203] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_204 bl[204] br[204] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_205 bl[205] br[205] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_206 bl[206] br[206] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_207 bl[207] br[207] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_208 bl[208] br[208] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_209 bl[209] br[209] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_210 bl[210] br[210] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_211 bl[211] br[211] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_212 bl[212] br[212] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_213 bl[213] br[213] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_214 bl[214] br[214] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_215 bl[215] br[215] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_216 bl[216] br[216] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_217 bl[217] br[217] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_218 bl[218] br[218] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_219 bl[219] br[219] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_220 bl[220] br[220] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_221 bl[221] br[221] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_222 bl[222] br[222] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_223 bl[223] br[223] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_224 bl[224] br[224] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_225 bl[225] br[225] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_226 bl[226] br[226] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_227 bl[227] br[227] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_228 bl[228] br[228] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_229 bl[229] br[229] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_230 bl[230] br[230] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_231 bl[231] br[231] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_232 bl[232] br[232] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_233 bl[233] br[233] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_234 bl[234] br[234] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_235 bl[235] br[235] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_236 bl[236] br[236] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_237 bl[237] br[237] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_238 bl[238] br[238] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_239 bl[239] br[239] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_240 bl[240] br[240] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_241 bl[241] br[241] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_242 bl[242] br[242] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_243 bl[243] br[243] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_244 bl[244] br[244] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_245 bl[245] br[245] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_246 bl[246] br[246] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_247 bl[247] br[247] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_248 bl[248] br[248] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_249 bl[249] br[249] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_250 bl[250] br[250] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_251 bl[251] br[251] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_252 bl[252] br[252] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_253 bl[253] br[253] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_254 bl[254] br[254] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_255 bl[255] br[255] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_4_0 bl[0] br[0] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_1 bl[1] br[1] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_2 bl[2] br[2] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_3 bl[3] br[3] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_4 bl[4] br[4] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_5 bl[5] br[5] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_6 bl[6] br[6] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_7 bl[7] br[7] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_8 bl[8] br[8] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_9 bl[9] br[9] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_10 bl[10] br[10] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_11 bl[11] br[11] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_12 bl[12] br[12] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_13 bl[13] br[13] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_14 bl[14] br[14] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_15 bl[15] br[15] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_16 bl[16] br[16] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_17 bl[17] br[17] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_18 bl[18] br[18] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_19 bl[19] br[19] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_20 bl[20] br[20] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_21 bl[21] br[21] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_22 bl[22] br[22] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_23 bl[23] br[23] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_24 bl[24] br[24] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_25 bl[25] br[25] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_26 bl[26] br[26] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_27 bl[27] br[27] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_28 bl[28] br[28] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_29 bl[29] br[29] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_30 bl[30] br[30] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_31 bl[31] br[31] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_32 bl[32] br[32] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_33 bl[33] br[33] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_34 bl[34] br[34] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_35 bl[35] br[35] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_36 bl[36] br[36] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_37 bl[37] br[37] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_38 bl[38] br[38] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_39 bl[39] br[39] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_40 bl[40] br[40] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_41 bl[41] br[41] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_42 bl[42] br[42] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_43 bl[43] br[43] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_44 bl[44] br[44] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_45 bl[45] br[45] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_46 bl[46] br[46] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_47 bl[47] br[47] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_48 bl[48] br[48] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_49 bl[49] br[49] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_50 bl[50] br[50] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_51 bl[51] br[51] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_52 bl[52] br[52] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_53 bl[53] br[53] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_54 bl[54] br[54] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_55 bl[55] br[55] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_56 bl[56] br[56] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_57 bl[57] br[57] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_58 bl[58] br[58] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_59 bl[59] br[59] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_60 bl[60] br[60] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_61 bl[61] br[61] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_62 bl[62] br[62] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_63 bl[63] br[63] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_64 bl[64] br[64] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_65 bl[65] br[65] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_66 bl[66] br[66] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_67 bl[67] br[67] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_68 bl[68] br[68] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_69 bl[69] br[69] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_70 bl[70] br[70] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_71 bl[71] br[71] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_72 bl[72] br[72] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_73 bl[73] br[73] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_74 bl[74] br[74] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_75 bl[75] br[75] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_76 bl[76] br[76] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_77 bl[77] br[77] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_78 bl[78] br[78] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_79 bl[79] br[79] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_80 bl[80] br[80] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_81 bl[81] br[81] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_82 bl[82] br[82] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_83 bl[83] br[83] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_84 bl[84] br[84] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_85 bl[85] br[85] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_86 bl[86] br[86] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_87 bl[87] br[87] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_88 bl[88] br[88] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_89 bl[89] br[89] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_90 bl[90] br[90] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_91 bl[91] br[91] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_92 bl[92] br[92] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_93 bl[93] br[93] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_94 bl[94] br[94] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_95 bl[95] br[95] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_96 bl[96] br[96] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_97 bl[97] br[97] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_98 bl[98] br[98] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_99 bl[99] br[99] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_100 bl[100] br[100] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_101 bl[101] br[101] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_102 bl[102] br[102] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_103 bl[103] br[103] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_104 bl[104] br[104] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_105 bl[105] br[105] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_106 bl[106] br[106] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_107 bl[107] br[107] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_108 bl[108] br[108] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_109 bl[109] br[109] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_110 bl[110] br[110] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_111 bl[111] br[111] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_112 bl[112] br[112] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_113 bl[113] br[113] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_114 bl[114] br[114] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_115 bl[115] br[115] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_116 bl[116] br[116] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_117 bl[117] br[117] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_118 bl[118] br[118] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_119 bl[119] br[119] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_120 bl[120] br[120] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_121 bl[121] br[121] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_122 bl[122] br[122] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_123 bl[123] br[123] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_124 bl[124] br[124] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_125 bl[125] br[125] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_126 bl[126] br[126] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_127 bl[127] br[127] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_128 bl[128] br[128] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_129 bl[129] br[129] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_130 bl[130] br[130] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_131 bl[131] br[131] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_132 bl[132] br[132] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_133 bl[133] br[133] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_134 bl[134] br[134] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_135 bl[135] br[135] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_136 bl[136] br[136] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_137 bl[137] br[137] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_138 bl[138] br[138] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_139 bl[139] br[139] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_140 bl[140] br[140] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_141 bl[141] br[141] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_142 bl[142] br[142] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_143 bl[143] br[143] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_144 bl[144] br[144] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_145 bl[145] br[145] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_146 bl[146] br[146] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_147 bl[147] br[147] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_148 bl[148] br[148] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_149 bl[149] br[149] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_150 bl[150] br[150] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_151 bl[151] br[151] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_152 bl[152] br[152] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_153 bl[153] br[153] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_154 bl[154] br[154] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_155 bl[155] br[155] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_156 bl[156] br[156] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_157 bl[157] br[157] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_158 bl[158] br[158] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_159 bl[159] br[159] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_160 bl[160] br[160] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_161 bl[161] br[161] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_162 bl[162] br[162] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_163 bl[163] br[163] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_164 bl[164] br[164] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_165 bl[165] br[165] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_166 bl[166] br[166] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_167 bl[167] br[167] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_168 bl[168] br[168] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_169 bl[169] br[169] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_170 bl[170] br[170] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_171 bl[171] br[171] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_172 bl[172] br[172] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_173 bl[173] br[173] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_174 bl[174] br[174] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_175 bl[175] br[175] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_176 bl[176] br[176] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_177 bl[177] br[177] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_178 bl[178] br[178] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_179 bl[179] br[179] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_180 bl[180] br[180] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_181 bl[181] br[181] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_182 bl[182] br[182] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_183 bl[183] br[183] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_184 bl[184] br[184] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_185 bl[185] br[185] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_186 bl[186] br[186] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_187 bl[187] br[187] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_188 bl[188] br[188] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_189 bl[189] br[189] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_190 bl[190] br[190] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_191 bl[191] br[191] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_192 bl[192] br[192] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_193 bl[193] br[193] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_194 bl[194] br[194] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_195 bl[195] br[195] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_196 bl[196] br[196] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_197 bl[197] br[197] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_198 bl[198] br[198] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_199 bl[199] br[199] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_200 bl[200] br[200] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_201 bl[201] br[201] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_202 bl[202] br[202] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_203 bl[203] br[203] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_204 bl[204] br[204] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_205 bl[205] br[205] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_206 bl[206] br[206] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_207 bl[207] br[207] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_208 bl[208] br[208] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_209 bl[209] br[209] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_210 bl[210] br[210] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_211 bl[211] br[211] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_212 bl[212] br[212] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_213 bl[213] br[213] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_214 bl[214] br[214] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_215 bl[215] br[215] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_216 bl[216] br[216] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_217 bl[217] br[217] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_218 bl[218] br[218] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_219 bl[219] br[219] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_220 bl[220] br[220] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_221 bl[221] br[221] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_222 bl[222] br[222] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_223 bl[223] br[223] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_224 bl[224] br[224] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_225 bl[225] br[225] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_226 bl[226] br[226] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_227 bl[227] br[227] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_228 bl[228] br[228] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_229 bl[229] br[229] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_230 bl[230] br[230] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_231 bl[231] br[231] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_232 bl[232] br[232] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_233 bl[233] br[233] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_234 bl[234] br[234] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_235 bl[235] br[235] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_236 bl[236] br[236] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_237 bl[237] br[237] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_238 bl[238] br[238] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_239 bl[239] br[239] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_240 bl[240] br[240] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_241 bl[241] br[241] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_242 bl[242] br[242] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_243 bl[243] br[243] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_244 bl[244] br[244] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_245 bl[245] br[245] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_246 bl[246] br[246] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_247 bl[247] br[247] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_248 bl[248] br[248] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_249 bl[249] br[249] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_250 bl[250] br[250] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_251 bl[251] br[251] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_252 bl[252] br[252] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_253 bl[253] br[253] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_254 bl[254] br[254] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_255 bl[255] br[255] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_5_0 bl[0] br[0] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_1 bl[1] br[1] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_2 bl[2] br[2] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_3 bl[3] br[3] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_4 bl[4] br[4] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_5 bl[5] br[5] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_6 bl[6] br[6] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_7 bl[7] br[7] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_8 bl[8] br[8] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_9 bl[9] br[9] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_10 bl[10] br[10] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_11 bl[11] br[11] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_12 bl[12] br[12] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_13 bl[13] br[13] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_14 bl[14] br[14] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_15 bl[15] br[15] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_16 bl[16] br[16] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_17 bl[17] br[17] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_18 bl[18] br[18] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_19 bl[19] br[19] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_20 bl[20] br[20] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_21 bl[21] br[21] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_22 bl[22] br[22] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_23 bl[23] br[23] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_24 bl[24] br[24] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_25 bl[25] br[25] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_26 bl[26] br[26] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_27 bl[27] br[27] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_28 bl[28] br[28] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_29 bl[29] br[29] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_30 bl[30] br[30] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_31 bl[31] br[31] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_32 bl[32] br[32] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_33 bl[33] br[33] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_34 bl[34] br[34] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_35 bl[35] br[35] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_36 bl[36] br[36] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_37 bl[37] br[37] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_38 bl[38] br[38] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_39 bl[39] br[39] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_40 bl[40] br[40] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_41 bl[41] br[41] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_42 bl[42] br[42] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_43 bl[43] br[43] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_44 bl[44] br[44] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_45 bl[45] br[45] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_46 bl[46] br[46] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_47 bl[47] br[47] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_48 bl[48] br[48] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_49 bl[49] br[49] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_50 bl[50] br[50] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_51 bl[51] br[51] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_52 bl[52] br[52] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_53 bl[53] br[53] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_54 bl[54] br[54] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_55 bl[55] br[55] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_56 bl[56] br[56] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_57 bl[57] br[57] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_58 bl[58] br[58] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_59 bl[59] br[59] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_60 bl[60] br[60] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_61 bl[61] br[61] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_62 bl[62] br[62] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_63 bl[63] br[63] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_64 bl[64] br[64] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_65 bl[65] br[65] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_66 bl[66] br[66] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_67 bl[67] br[67] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_68 bl[68] br[68] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_69 bl[69] br[69] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_70 bl[70] br[70] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_71 bl[71] br[71] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_72 bl[72] br[72] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_73 bl[73] br[73] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_74 bl[74] br[74] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_75 bl[75] br[75] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_76 bl[76] br[76] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_77 bl[77] br[77] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_78 bl[78] br[78] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_79 bl[79] br[79] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_80 bl[80] br[80] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_81 bl[81] br[81] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_82 bl[82] br[82] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_83 bl[83] br[83] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_84 bl[84] br[84] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_85 bl[85] br[85] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_86 bl[86] br[86] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_87 bl[87] br[87] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_88 bl[88] br[88] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_89 bl[89] br[89] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_90 bl[90] br[90] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_91 bl[91] br[91] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_92 bl[92] br[92] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_93 bl[93] br[93] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_94 bl[94] br[94] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_95 bl[95] br[95] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_96 bl[96] br[96] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_97 bl[97] br[97] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_98 bl[98] br[98] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_99 bl[99] br[99] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_100 bl[100] br[100] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_101 bl[101] br[101] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_102 bl[102] br[102] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_103 bl[103] br[103] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_104 bl[104] br[104] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_105 bl[105] br[105] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_106 bl[106] br[106] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_107 bl[107] br[107] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_108 bl[108] br[108] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_109 bl[109] br[109] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_110 bl[110] br[110] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_111 bl[111] br[111] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_112 bl[112] br[112] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_113 bl[113] br[113] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_114 bl[114] br[114] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_115 bl[115] br[115] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_116 bl[116] br[116] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_117 bl[117] br[117] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_118 bl[118] br[118] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_119 bl[119] br[119] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_120 bl[120] br[120] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_121 bl[121] br[121] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_122 bl[122] br[122] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_123 bl[123] br[123] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_124 bl[124] br[124] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_125 bl[125] br[125] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_126 bl[126] br[126] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_127 bl[127] br[127] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_128 bl[128] br[128] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_129 bl[129] br[129] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_130 bl[130] br[130] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_131 bl[131] br[131] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_132 bl[132] br[132] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_133 bl[133] br[133] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_134 bl[134] br[134] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_135 bl[135] br[135] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_136 bl[136] br[136] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_137 bl[137] br[137] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_138 bl[138] br[138] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_139 bl[139] br[139] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_140 bl[140] br[140] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_141 bl[141] br[141] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_142 bl[142] br[142] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_143 bl[143] br[143] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_144 bl[144] br[144] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_145 bl[145] br[145] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_146 bl[146] br[146] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_147 bl[147] br[147] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_148 bl[148] br[148] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_149 bl[149] br[149] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_150 bl[150] br[150] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_151 bl[151] br[151] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_152 bl[152] br[152] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_153 bl[153] br[153] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_154 bl[154] br[154] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_155 bl[155] br[155] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_156 bl[156] br[156] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_157 bl[157] br[157] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_158 bl[158] br[158] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_159 bl[159] br[159] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_160 bl[160] br[160] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_161 bl[161] br[161] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_162 bl[162] br[162] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_163 bl[163] br[163] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_164 bl[164] br[164] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_165 bl[165] br[165] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_166 bl[166] br[166] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_167 bl[167] br[167] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_168 bl[168] br[168] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_169 bl[169] br[169] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_170 bl[170] br[170] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_171 bl[171] br[171] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_172 bl[172] br[172] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_173 bl[173] br[173] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_174 bl[174] br[174] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_175 bl[175] br[175] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_176 bl[176] br[176] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_177 bl[177] br[177] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_178 bl[178] br[178] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_179 bl[179] br[179] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_180 bl[180] br[180] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_181 bl[181] br[181] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_182 bl[182] br[182] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_183 bl[183] br[183] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_184 bl[184] br[184] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_185 bl[185] br[185] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_186 bl[186] br[186] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_187 bl[187] br[187] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_188 bl[188] br[188] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_189 bl[189] br[189] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_190 bl[190] br[190] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_191 bl[191] br[191] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_192 bl[192] br[192] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_193 bl[193] br[193] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_194 bl[194] br[194] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_195 bl[195] br[195] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_196 bl[196] br[196] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_197 bl[197] br[197] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_198 bl[198] br[198] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_199 bl[199] br[199] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_200 bl[200] br[200] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_201 bl[201] br[201] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_202 bl[202] br[202] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_203 bl[203] br[203] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_204 bl[204] br[204] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_205 bl[205] br[205] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_206 bl[206] br[206] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_207 bl[207] br[207] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_208 bl[208] br[208] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_209 bl[209] br[209] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_210 bl[210] br[210] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_211 bl[211] br[211] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_212 bl[212] br[212] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_213 bl[213] br[213] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_214 bl[214] br[214] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_215 bl[215] br[215] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_216 bl[216] br[216] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_217 bl[217] br[217] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_218 bl[218] br[218] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_219 bl[219] br[219] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_220 bl[220] br[220] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_221 bl[221] br[221] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_222 bl[222] br[222] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_223 bl[223] br[223] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_224 bl[224] br[224] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_225 bl[225] br[225] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_226 bl[226] br[226] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_227 bl[227] br[227] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_228 bl[228] br[228] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_229 bl[229] br[229] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_230 bl[230] br[230] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_231 bl[231] br[231] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_232 bl[232] br[232] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_233 bl[233] br[233] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_234 bl[234] br[234] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_235 bl[235] br[235] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_236 bl[236] br[236] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_237 bl[237] br[237] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_238 bl[238] br[238] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_239 bl[239] br[239] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_240 bl[240] br[240] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_241 bl[241] br[241] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_242 bl[242] br[242] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_243 bl[243] br[243] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_244 bl[244] br[244] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_245 bl[245] br[245] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_246 bl[246] br[246] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_247 bl[247] br[247] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_248 bl[248] br[248] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_249 bl[249] br[249] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_250 bl[250] br[250] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_251 bl[251] br[251] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_252 bl[252] br[252] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_253 bl[253] br[253] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_254 bl[254] br[254] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_255 bl[255] br[255] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_6_0 bl[0] br[0] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_1 bl[1] br[1] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_2 bl[2] br[2] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_3 bl[3] br[3] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_4 bl[4] br[4] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_5 bl[5] br[5] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_6 bl[6] br[6] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_7 bl[7] br[7] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_8 bl[8] br[8] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_9 bl[9] br[9] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_10 bl[10] br[10] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_11 bl[11] br[11] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_12 bl[12] br[12] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_13 bl[13] br[13] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_14 bl[14] br[14] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_15 bl[15] br[15] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_16 bl[16] br[16] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_17 bl[17] br[17] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_18 bl[18] br[18] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_19 bl[19] br[19] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_20 bl[20] br[20] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_21 bl[21] br[21] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_22 bl[22] br[22] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_23 bl[23] br[23] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_24 bl[24] br[24] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_25 bl[25] br[25] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_26 bl[26] br[26] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_27 bl[27] br[27] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_28 bl[28] br[28] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_29 bl[29] br[29] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_30 bl[30] br[30] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_31 bl[31] br[31] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_32 bl[32] br[32] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_33 bl[33] br[33] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_34 bl[34] br[34] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_35 bl[35] br[35] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_36 bl[36] br[36] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_37 bl[37] br[37] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_38 bl[38] br[38] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_39 bl[39] br[39] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_40 bl[40] br[40] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_41 bl[41] br[41] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_42 bl[42] br[42] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_43 bl[43] br[43] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_44 bl[44] br[44] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_45 bl[45] br[45] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_46 bl[46] br[46] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_47 bl[47] br[47] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_48 bl[48] br[48] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_49 bl[49] br[49] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_50 bl[50] br[50] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_51 bl[51] br[51] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_52 bl[52] br[52] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_53 bl[53] br[53] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_54 bl[54] br[54] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_55 bl[55] br[55] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_56 bl[56] br[56] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_57 bl[57] br[57] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_58 bl[58] br[58] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_59 bl[59] br[59] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_60 bl[60] br[60] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_61 bl[61] br[61] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_62 bl[62] br[62] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_63 bl[63] br[63] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_64 bl[64] br[64] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_65 bl[65] br[65] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_66 bl[66] br[66] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_67 bl[67] br[67] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_68 bl[68] br[68] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_69 bl[69] br[69] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_70 bl[70] br[70] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_71 bl[71] br[71] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_72 bl[72] br[72] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_73 bl[73] br[73] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_74 bl[74] br[74] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_75 bl[75] br[75] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_76 bl[76] br[76] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_77 bl[77] br[77] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_78 bl[78] br[78] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_79 bl[79] br[79] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_80 bl[80] br[80] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_81 bl[81] br[81] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_82 bl[82] br[82] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_83 bl[83] br[83] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_84 bl[84] br[84] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_85 bl[85] br[85] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_86 bl[86] br[86] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_87 bl[87] br[87] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_88 bl[88] br[88] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_89 bl[89] br[89] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_90 bl[90] br[90] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_91 bl[91] br[91] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_92 bl[92] br[92] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_93 bl[93] br[93] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_94 bl[94] br[94] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_95 bl[95] br[95] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_96 bl[96] br[96] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_97 bl[97] br[97] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_98 bl[98] br[98] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_99 bl[99] br[99] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_100 bl[100] br[100] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_101 bl[101] br[101] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_102 bl[102] br[102] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_103 bl[103] br[103] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_104 bl[104] br[104] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_105 bl[105] br[105] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_106 bl[106] br[106] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_107 bl[107] br[107] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_108 bl[108] br[108] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_109 bl[109] br[109] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_110 bl[110] br[110] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_111 bl[111] br[111] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_112 bl[112] br[112] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_113 bl[113] br[113] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_114 bl[114] br[114] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_115 bl[115] br[115] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_116 bl[116] br[116] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_117 bl[117] br[117] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_118 bl[118] br[118] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_119 bl[119] br[119] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_120 bl[120] br[120] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_121 bl[121] br[121] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_122 bl[122] br[122] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_123 bl[123] br[123] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_124 bl[124] br[124] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_125 bl[125] br[125] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_126 bl[126] br[126] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_127 bl[127] br[127] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_128 bl[128] br[128] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_129 bl[129] br[129] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_130 bl[130] br[130] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_131 bl[131] br[131] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_132 bl[132] br[132] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_133 bl[133] br[133] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_134 bl[134] br[134] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_135 bl[135] br[135] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_136 bl[136] br[136] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_137 bl[137] br[137] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_138 bl[138] br[138] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_139 bl[139] br[139] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_140 bl[140] br[140] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_141 bl[141] br[141] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_142 bl[142] br[142] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_143 bl[143] br[143] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_144 bl[144] br[144] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_145 bl[145] br[145] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_146 bl[146] br[146] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_147 bl[147] br[147] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_148 bl[148] br[148] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_149 bl[149] br[149] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_150 bl[150] br[150] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_151 bl[151] br[151] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_152 bl[152] br[152] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_153 bl[153] br[153] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_154 bl[154] br[154] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_155 bl[155] br[155] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_156 bl[156] br[156] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_157 bl[157] br[157] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_158 bl[158] br[158] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_159 bl[159] br[159] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_160 bl[160] br[160] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_161 bl[161] br[161] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_162 bl[162] br[162] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_163 bl[163] br[163] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_164 bl[164] br[164] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_165 bl[165] br[165] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_166 bl[166] br[166] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_167 bl[167] br[167] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_168 bl[168] br[168] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_169 bl[169] br[169] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_170 bl[170] br[170] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_171 bl[171] br[171] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_172 bl[172] br[172] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_173 bl[173] br[173] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_174 bl[174] br[174] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_175 bl[175] br[175] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_176 bl[176] br[176] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_177 bl[177] br[177] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_178 bl[178] br[178] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_179 bl[179] br[179] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_180 bl[180] br[180] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_181 bl[181] br[181] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_182 bl[182] br[182] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_183 bl[183] br[183] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_184 bl[184] br[184] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_185 bl[185] br[185] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_186 bl[186] br[186] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_187 bl[187] br[187] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_188 bl[188] br[188] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_189 bl[189] br[189] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_190 bl[190] br[190] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_191 bl[191] br[191] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_192 bl[192] br[192] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_193 bl[193] br[193] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_194 bl[194] br[194] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_195 bl[195] br[195] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_196 bl[196] br[196] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_197 bl[197] br[197] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_198 bl[198] br[198] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_199 bl[199] br[199] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_200 bl[200] br[200] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_201 bl[201] br[201] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_202 bl[202] br[202] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_203 bl[203] br[203] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_204 bl[204] br[204] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_205 bl[205] br[205] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_206 bl[206] br[206] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_207 bl[207] br[207] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_208 bl[208] br[208] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_209 bl[209] br[209] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_210 bl[210] br[210] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_211 bl[211] br[211] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_212 bl[212] br[212] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_213 bl[213] br[213] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_214 bl[214] br[214] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_215 bl[215] br[215] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_216 bl[216] br[216] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_217 bl[217] br[217] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_218 bl[218] br[218] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_219 bl[219] br[219] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_220 bl[220] br[220] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_221 bl[221] br[221] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_222 bl[222] br[222] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_223 bl[223] br[223] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_224 bl[224] br[224] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_225 bl[225] br[225] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_226 bl[226] br[226] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_227 bl[227] br[227] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_228 bl[228] br[228] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_229 bl[229] br[229] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_230 bl[230] br[230] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_231 bl[231] br[231] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_232 bl[232] br[232] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_233 bl[233] br[233] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_234 bl[234] br[234] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_235 bl[235] br[235] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_236 bl[236] br[236] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_237 bl[237] br[237] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_238 bl[238] br[238] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_239 bl[239] br[239] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_240 bl[240] br[240] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_241 bl[241] br[241] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_242 bl[242] br[242] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_243 bl[243] br[243] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_244 bl[244] br[244] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_245 bl[245] br[245] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_246 bl[246] br[246] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_247 bl[247] br[247] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_248 bl[248] br[248] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_249 bl[249] br[249] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_250 bl[250] br[250] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_251 bl[251] br[251] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_252 bl[252] br[252] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_253 bl[253] br[253] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_254 bl[254] br[254] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_255 bl[255] br[255] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_7_0 bl[0] br[0] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_1 bl[1] br[1] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_2 bl[2] br[2] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_3 bl[3] br[3] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_4 bl[4] br[4] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_5 bl[5] br[5] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_6 bl[6] br[6] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_7 bl[7] br[7] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_8 bl[8] br[8] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_9 bl[9] br[9] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_10 bl[10] br[10] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_11 bl[11] br[11] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_12 bl[12] br[12] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_13 bl[13] br[13] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_14 bl[14] br[14] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_15 bl[15] br[15] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_16 bl[16] br[16] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_17 bl[17] br[17] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_18 bl[18] br[18] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_19 bl[19] br[19] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_20 bl[20] br[20] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_21 bl[21] br[21] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_22 bl[22] br[22] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_23 bl[23] br[23] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_24 bl[24] br[24] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_25 bl[25] br[25] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_26 bl[26] br[26] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_27 bl[27] br[27] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_28 bl[28] br[28] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_29 bl[29] br[29] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_30 bl[30] br[30] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_31 bl[31] br[31] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_32 bl[32] br[32] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_33 bl[33] br[33] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_34 bl[34] br[34] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_35 bl[35] br[35] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_36 bl[36] br[36] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_37 bl[37] br[37] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_38 bl[38] br[38] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_39 bl[39] br[39] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_40 bl[40] br[40] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_41 bl[41] br[41] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_42 bl[42] br[42] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_43 bl[43] br[43] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_44 bl[44] br[44] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_45 bl[45] br[45] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_46 bl[46] br[46] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_47 bl[47] br[47] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_48 bl[48] br[48] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_49 bl[49] br[49] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_50 bl[50] br[50] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_51 bl[51] br[51] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_52 bl[52] br[52] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_53 bl[53] br[53] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_54 bl[54] br[54] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_55 bl[55] br[55] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_56 bl[56] br[56] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_57 bl[57] br[57] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_58 bl[58] br[58] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_59 bl[59] br[59] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_60 bl[60] br[60] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_61 bl[61] br[61] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_62 bl[62] br[62] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_63 bl[63] br[63] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_64 bl[64] br[64] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_65 bl[65] br[65] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_66 bl[66] br[66] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_67 bl[67] br[67] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_68 bl[68] br[68] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_69 bl[69] br[69] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_70 bl[70] br[70] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_71 bl[71] br[71] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_72 bl[72] br[72] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_73 bl[73] br[73] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_74 bl[74] br[74] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_75 bl[75] br[75] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_76 bl[76] br[76] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_77 bl[77] br[77] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_78 bl[78] br[78] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_79 bl[79] br[79] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_80 bl[80] br[80] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_81 bl[81] br[81] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_82 bl[82] br[82] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_83 bl[83] br[83] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_84 bl[84] br[84] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_85 bl[85] br[85] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_86 bl[86] br[86] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_87 bl[87] br[87] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_88 bl[88] br[88] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_89 bl[89] br[89] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_90 bl[90] br[90] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_91 bl[91] br[91] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_92 bl[92] br[92] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_93 bl[93] br[93] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_94 bl[94] br[94] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_95 bl[95] br[95] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_96 bl[96] br[96] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_97 bl[97] br[97] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_98 bl[98] br[98] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_99 bl[99] br[99] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_100 bl[100] br[100] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_101 bl[101] br[101] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_102 bl[102] br[102] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_103 bl[103] br[103] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_104 bl[104] br[104] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_105 bl[105] br[105] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_106 bl[106] br[106] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_107 bl[107] br[107] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_108 bl[108] br[108] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_109 bl[109] br[109] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_110 bl[110] br[110] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_111 bl[111] br[111] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_112 bl[112] br[112] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_113 bl[113] br[113] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_114 bl[114] br[114] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_115 bl[115] br[115] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_116 bl[116] br[116] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_117 bl[117] br[117] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_118 bl[118] br[118] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_119 bl[119] br[119] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_120 bl[120] br[120] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_121 bl[121] br[121] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_122 bl[122] br[122] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_123 bl[123] br[123] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_124 bl[124] br[124] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_125 bl[125] br[125] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_126 bl[126] br[126] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_127 bl[127] br[127] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_128 bl[128] br[128] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_129 bl[129] br[129] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_130 bl[130] br[130] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_131 bl[131] br[131] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_132 bl[132] br[132] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_133 bl[133] br[133] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_134 bl[134] br[134] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_135 bl[135] br[135] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_136 bl[136] br[136] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_137 bl[137] br[137] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_138 bl[138] br[138] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_139 bl[139] br[139] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_140 bl[140] br[140] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_141 bl[141] br[141] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_142 bl[142] br[142] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_143 bl[143] br[143] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_144 bl[144] br[144] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_145 bl[145] br[145] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_146 bl[146] br[146] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_147 bl[147] br[147] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_148 bl[148] br[148] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_149 bl[149] br[149] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_150 bl[150] br[150] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_151 bl[151] br[151] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_152 bl[152] br[152] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_153 bl[153] br[153] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_154 bl[154] br[154] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_155 bl[155] br[155] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_156 bl[156] br[156] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_157 bl[157] br[157] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_158 bl[158] br[158] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_159 bl[159] br[159] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_160 bl[160] br[160] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_161 bl[161] br[161] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_162 bl[162] br[162] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_163 bl[163] br[163] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_164 bl[164] br[164] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_165 bl[165] br[165] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_166 bl[166] br[166] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_167 bl[167] br[167] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_168 bl[168] br[168] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_169 bl[169] br[169] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_170 bl[170] br[170] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_171 bl[171] br[171] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_172 bl[172] br[172] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_173 bl[173] br[173] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_174 bl[174] br[174] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_175 bl[175] br[175] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_176 bl[176] br[176] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_177 bl[177] br[177] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_178 bl[178] br[178] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_179 bl[179] br[179] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_180 bl[180] br[180] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_181 bl[181] br[181] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_182 bl[182] br[182] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_183 bl[183] br[183] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_184 bl[184] br[184] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_185 bl[185] br[185] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_186 bl[186] br[186] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_187 bl[187] br[187] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_188 bl[188] br[188] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_189 bl[189] br[189] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_190 bl[190] br[190] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_191 bl[191] br[191] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_192 bl[192] br[192] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_193 bl[193] br[193] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_194 bl[194] br[194] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_195 bl[195] br[195] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_196 bl[196] br[196] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_197 bl[197] br[197] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_198 bl[198] br[198] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_199 bl[199] br[199] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_200 bl[200] br[200] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_201 bl[201] br[201] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_202 bl[202] br[202] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_203 bl[203] br[203] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_204 bl[204] br[204] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_205 bl[205] br[205] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_206 bl[206] br[206] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_207 bl[207] br[207] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_208 bl[208] br[208] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_209 bl[209] br[209] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_210 bl[210] br[210] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_211 bl[211] br[211] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_212 bl[212] br[212] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_213 bl[213] br[213] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_214 bl[214] br[214] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_215 bl[215] br[215] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_216 bl[216] br[216] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_217 bl[217] br[217] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_218 bl[218] br[218] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_219 bl[219] br[219] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_220 bl[220] br[220] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_221 bl[221] br[221] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_222 bl[222] br[222] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_223 bl[223] br[223] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_224 bl[224] br[224] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_225 bl[225] br[225] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_226 bl[226] br[226] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_227 bl[227] br[227] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_228 bl[228] br[228] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_229 bl[229] br[229] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_230 bl[230] br[230] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_231 bl[231] br[231] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_232 bl[232] br[232] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_233 bl[233] br[233] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_234 bl[234] br[234] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_235 bl[235] br[235] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_236 bl[236] br[236] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_237 bl[237] br[237] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_238 bl[238] br[238] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_239 bl[239] br[239] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_240 bl[240] br[240] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_241 bl[241] br[241] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_242 bl[242] br[242] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_243 bl[243] br[243] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_244 bl[244] br[244] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_245 bl[245] br[245] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_246 bl[246] br[246] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_247 bl[247] br[247] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_248 bl[248] br[248] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_249 bl[249] br[249] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_250 bl[250] br[250] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_251 bl[251] br[251] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_252 bl[252] br[252] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_253 bl[253] br[253] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_254 bl[254] br[254] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_255 bl[255] br[255] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_8_0 bl[0] br[0] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_1 bl[1] br[1] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_2 bl[2] br[2] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_3 bl[3] br[3] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_4 bl[4] br[4] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_5 bl[5] br[5] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_6 bl[6] br[6] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_7 bl[7] br[7] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_8 bl[8] br[8] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_9 bl[9] br[9] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_10 bl[10] br[10] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_11 bl[11] br[11] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_12 bl[12] br[12] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_13 bl[13] br[13] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_14 bl[14] br[14] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_15 bl[15] br[15] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_16 bl[16] br[16] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_17 bl[17] br[17] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_18 bl[18] br[18] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_19 bl[19] br[19] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_20 bl[20] br[20] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_21 bl[21] br[21] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_22 bl[22] br[22] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_23 bl[23] br[23] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_24 bl[24] br[24] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_25 bl[25] br[25] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_26 bl[26] br[26] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_27 bl[27] br[27] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_28 bl[28] br[28] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_29 bl[29] br[29] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_30 bl[30] br[30] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_31 bl[31] br[31] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_32 bl[32] br[32] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_33 bl[33] br[33] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_34 bl[34] br[34] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_35 bl[35] br[35] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_36 bl[36] br[36] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_37 bl[37] br[37] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_38 bl[38] br[38] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_39 bl[39] br[39] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_40 bl[40] br[40] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_41 bl[41] br[41] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_42 bl[42] br[42] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_43 bl[43] br[43] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_44 bl[44] br[44] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_45 bl[45] br[45] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_46 bl[46] br[46] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_47 bl[47] br[47] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_48 bl[48] br[48] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_49 bl[49] br[49] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_50 bl[50] br[50] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_51 bl[51] br[51] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_52 bl[52] br[52] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_53 bl[53] br[53] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_54 bl[54] br[54] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_55 bl[55] br[55] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_56 bl[56] br[56] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_57 bl[57] br[57] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_58 bl[58] br[58] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_59 bl[59] br[59] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_60 bl[60] br[60] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_61 bl[61] br[61] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_62 bl[62] br[62] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_63 bl[63] br[63] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_64 bl[64] br[64] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_65 bl[65] br[65] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_66 bl[66] br[66] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_67 bl[67] br[67] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_68 bl[68] br[68] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_69 bl[69] br[69] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_70 bl[70] br[70] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_71 bl[71] br[71] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_72 bl[72] br[72] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_73 bl[73] br[73] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_74 bl[74] br[74] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_75 bl[75] br[75] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_76 bl[76] br[76] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_77 bl[77] br[77] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_78 bl[78] br[78] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_79 bl[79] br[79] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_80 bl[80] br[80] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_81 bl[81] br[81] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_82 bl[82] br[82] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_83 bl[83] br[83] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_84 bl[84] br[84] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_85 bl[85] br[85] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_86 bl[86] br[86] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_87 bl[87] br[87] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_88 bl[88] br[88] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_89 bl[89] br[89] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_90 bl[90] br[90] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_91 bl[91] br[91] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_92 bl[92] br[92] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_93 bl[93] br[93] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_94 bl[94] br[94] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_95 bl[95] br[95] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_96 bl[96] br[96] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_97 bl[97] br[97] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_98 bl[98] br[98] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_99 bl[99] br[99] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_100 bl[100] br[100] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_101 bl[101] br[101] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_102 bl[102] br[102] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_103 bl[103] br[103] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_104 bl[104] br[104] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_105 bl[105] br[105] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_106 bl[106] br[106] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_107 bl[107] br[107] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_108 bl[108] br[108] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_109 bl[109] br[109] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_110 bl[110] br[110] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_111 bl[111] br[111] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_112 bl[112] br[112] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_113 bl[113] br[113] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_114 bl[114] br[114] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_115 bl[115] br[115] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_116 bl[116] br[116] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_117 bl[117] br[117] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_118 bl[118] br[118] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_119 bl[119] br[119] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_120 bl[120] br[120] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_121 bl[121] br[121] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_122 bl[122] br[122] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_123 bl[123] br[123] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_124 bl[124] br[124] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_125 bl[125] br[125] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_126 bl[126] br[126] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_127 bl[127] br[127] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_128 bl[128] br[128] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_129 bl[129] br[129] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_130 bl[130] br[130] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_131 bl[131] br[131] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_132 bl[132] br[132] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_133 bl[133] br[133] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_134 bl[134] br[134] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_135 bl[135] br[135] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_136 bl[136] br[136] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_137 bl[137] br[137] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_138 bl[138] br[138] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_139 bl[139] br[139] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_140 bl[140] br[140] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_141 bl[141] br[141] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_142 bl[142] br[142] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_143 bl[143] br[143] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_144 bl[144] br[144] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_145 bl[145] br[145] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_146 bl[146] br[146] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_147 bl[147] br[147] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_148 bl[148] br[148] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_149 bl[149] br[149] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_150 bl[150] br[150] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_151 bl[151] br[151] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_152 bl[152] br[152] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_153 bl[153] br[153] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_154 bl[154] br[154] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_155 bl[155] br[155] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_156 bl[156] br[156] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_157 bl[157] br[157] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_158 bl[158] br[158] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_159 bl[159] br[159] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_160 bl[160] br[160] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_161 bl[161] br[161] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_162 bl[162] br[162] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_163 bl[163] br[163] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_164 bl[164] br[164] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_165 bl[165] br[165] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_166 bl[166] br[166] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_167 bl[167] br[167] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_168 bl[168] br[168] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_169 bl[169] br[169] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_170 bl[170] br[170] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_171 bl[171] br[171] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_172 bl[172] br[172] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_173 bl[173] br[173] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_174 bl[174] br[174] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_175 bl[175] br[175] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_176 bl[176] br[176] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_177 bl[177] br[177] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_178 bl[178] br[178] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_179 bl[179] br[179] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_180 bl[180] br[180] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_181 bl[181] br[181] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_182 bl[182] br[182] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_183 bl[183] br[183] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_184 bl[184] br[184] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_185 bl[185] br[185] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_186 bl[186] br[186] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_187 bl[187] br[187] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_188 bl[188] br[188] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_189 bl[189] br[189] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_190 bl[190] br[190] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_191 bl[191] br[191] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_192 bl[192] br[192] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_193 bl[193] br[193] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_194 bl[194] br[194] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_195 bl[195] br[195] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_196 bl[196] br[196] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_197 bl[197] br[197] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_198 bl[198] br[198] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_199 bl[199] br[199] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_200 bl[200] br[200] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_201 bl[201] br[201] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_202 bl[202] br[202] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_203 bl[203] br[203] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_204 bl[204] br[204] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_205 bl[205] br[205] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_206 bl[206] br[206] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_207 bl[207] br[207] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_208 bl[208] br[208] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_209 bl[209] br[209] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_210 bl[210] br[210] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_211 bl[211] br[211] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_212 bl[212] br[212] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_213 bl[213] br[213] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_214 bl[214] br[214] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_215 bl[215] br[215] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_216 bl[216] br[216] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_217 bl[217] br[217] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_218 bl[218] br[218] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_219 bl[219] br[219] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_220 bl[220] br[220] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_221 bl[221] br[221] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_222 bl[222] br[222] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_223 bl[223] br[223] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_224 bl[224] br[224] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_225 bl[225] br[225] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_226 bl[226] br[226] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_227 bl[227] br[227] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_228 bl[228] br[228] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_229 bl[229] br[229] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_230 bl[230] br[230] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_231 bl[231] br[231] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_232 bl[232] br[232] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_233 bl[233] br[233] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_234 bl[234] br[234] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_235 bl[235] br[235] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_236 bl[236] br[236] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_237 bl[237] br[237] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_238 bl[238] br[238] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_239 bl[239] br[239] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_240 bl[240] br[240] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_241 bl[241] br[241] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_242 bl[242] br[242] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_243 bl[243] br[243] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_244 bl[244] br[244] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_245 bl[245] br[245] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_246 bl[246] br[246] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_247 bl[247] br[247] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_248 bl[248] br[248] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_249 bl[249] br[249] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_250 bl[250] br[250] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_251 bl[251] br[251] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_252 bl[252] br[252] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_253 bl[253] br[253] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_254 bl[254] br[254] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_255 bl[255] br[255] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_9_0 bl[0] br[0] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_1 bl[1] br[1] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_2 bl[2] br[2] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_3 bl[3] br[3] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_4 bl[4] br[4] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_5 bl[5] br[5] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_6 bl[6] br[6] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_7 bl[7] br[7] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_8 bl[8] br[8] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_9 bl[9] br[9] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_10 bl[10] br[10] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_11 bl[11] br[11] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_12 bl[12] br[12] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_13 bl[13] br[13] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_14 bl[14] br[14] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_15 bl[15] br[15] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_16 bl[16] br[16] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_17 bl[17] br[17] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_18 bl[18] br[18] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_19 bl[19] br[19] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_20 bl[20] br[20] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_21 bl[21] br[21] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_22 bl[22] br[22] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_23 bl[23] br[23] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_24 bl[24] br[24] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_25 bl[25] br[25] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_26 bl[26] br[26] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_27 bl[27] br[27] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_28 bl[28] br[28] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_29 bl[29] br[29] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_30 bl[30] br[30] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_31 bl[31] br[31] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_32 bl[32] br[32] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_33 bl[33] br[33] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_34 bl[34] br[34] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_35 bl[35] br[35] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_36 bl[36] br[36] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_37 bl[37] br[37] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_38 bl[38] br[38] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_39 bl[39] br[39] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_40 bl[40] br[40] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_41 bl[41] br[41] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_42 bl[42] br[42] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_43 bl[43] br[43] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_44 bl[44] br[44] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_45 bl[45] br[45] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_46 bl[46] br[46] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_47 bl[47] br[47] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_48 bl[48] br[48] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_49 bl[49] br[49] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_50 bl[50] br[50] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_51 bl[51] br[51] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_52 bl[52] br[52] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_53 bl[53] br[53] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_54 bl[54] br[54] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_55 bl[55] br[55] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_56 bl[56] br[56] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_57 bl[57] br[57] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_58 bl[58] br[58] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_59 bl[59] br[59] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_60 bl[60] br[60] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_61 bl[61] br[61] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_62 bl[62] br[62] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_63 bl[63] br[63] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_64 bl[64] br[64] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_65 bl[65] br[65] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_66 bl[66] br[66] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_67 bl[67] br[67] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_68 bl[68] br[68] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_69 bl[69] br[69] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_70 bl[70] br[70] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_71 bl[71] br[71] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_72 bl[72] br[72] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_73 bl[73] br[73] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_74 bl[74] br[74] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_75 bl[75] br[75] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_76 bl[76] br[76] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_77 bl[77] br[77] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_78 bl[78] br[78] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_79 bl[79] br[79] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_80 bl[80] br[80] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_81 bl[81] br[81] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_82 bl[82] br[82] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_83 bl[83] br[83] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_84 bl[84] br[84] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_85 bl[85] br[85] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_86 bl[86] br[86] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_87 bl[87] br[87] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_88 bl[88] br[88] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_89 bl[89] br[89] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_90 bl[90] br[90] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_91 bl[91] br[91] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_92 bl[92] br[92] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_93 bl[93] br[93] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_94 bl[94] br[94] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_95 bl[95] br[95] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_96 bl[96] br[96] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_97 bl[97] br[97] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_98 bl[98] br[98] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_99 bl[99] br[99] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_100 bl[100] br[100] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_101 bl[101] br[101] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_102 bl[102] br[102] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_103 bl[103] br[103] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_104 bl[104] br[104] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_105 bl[105] br[105] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_106 bl[106] br[106] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_107 bl[107] br[107] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_108 bl[108] br[108] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_109 bl[109] br[109] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_110 bl[110] br[110] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_111 bl[111] br[111] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_112 bl[112] br[112] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_113 bl[113] br[113] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_114 bl[114] br[114] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_115 bl[115] br[115] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_116 bl[116] br[116] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_117 bl[117] br[117] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_118 bl[118] br[118] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_119 bl[119] br[119] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_120 bl[120] br[120] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_121 bl[121] br[121] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_122 bl[122] br[122] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_123 bl[123] br[123] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_124 bl[124] br[124] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_125 bl[125] br[125] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_126 bl[126] br[126] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_127 bl[127] br[127] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_128 bl[128] br[128] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_129 bl[129] br[129] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_130 bl[130] br[130] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_131 bl[131] br[131] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_132 bl[132] br[132] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_133 bl[133] br[133] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_134 bl[134] br[134] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_135 bl[135] br[135] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_136 bl[136] br[136] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_137 bl[137] br[137] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_138 bl[138] br[138] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_139 bl[139] br[139] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_140 bl[140] br[140] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_141 bl[141] br[141] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_142 bl[142] br[142] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_143 bl[143] br[143] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_144 bl[144] br[144] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_145 bl[145] br[145] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_146 bl[146] br[146] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_147 bl[147] br[147] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_148 bl[148] br[148] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_149 bl[149] br[149] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_150 bl[150] br[150] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_151 bl[151] br[151] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_152 bl[152] br[152] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_153 bl[153] br[153] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_154 bl[154] br[154] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_155 bl[155] br[155] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_156 bl[156] br[156] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_157 bl[157] br[157] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_158 bl[158] br[158] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_159 bl[159] br[159] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_160 bl[160] br[160] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_161 bl[161] br[161] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_162 bl[162] br[162] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_163 bl[163] br[163] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_164 bl[164] br[164] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_165 bl[165] br[165] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_166 bl[166] br[166] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_167 bl[167] br[167] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_168 bl[168] br[168] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_169 bl[169] br[169] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_170 bl[170] br[170] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_171 bl[171] br[171] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_172 bl[172] br[172] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_173 bl[173] br[173] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_174 bl[174] br[174] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_175 bl[175] br[175] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_176 bl[176] br[176] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_177 bl[177] br[177] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_178 bl[178] br[178] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_179 bl[179] br[179] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_180 bl[180] br[180] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_181 bl[181] br[181] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_182 bl[182] br[182] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_183 bl[183] br[183] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_184 bl[184] br[184] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_185 bl[185] br[185] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_186 bl[186] br[186] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_187 bl[187] br[187] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_188 bl[188] br[188] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_189 bl[189] br[189] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_190 bl[190] br[190] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_191 bl[191] br[191] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_192 bl[192] br[192] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_193 bl[193] br[193] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_194 bl[194] br[194] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_195 bl[195] br[195] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_196 bl[196] br[196] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_197 bl[197] br[197] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_198 bl[198] br[198] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_199 bl[199] br[199] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_200 bl[200] br[200] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_201 bl[201] br[201] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_202 bl[202] br[202] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_203 bl[203] br[203] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_204 bl[204] br[204] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_205 bl[205] br[205] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_206 bl[206] br[206] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_207 bl[207] br[207] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_208 bl[208] br[208] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_209 bl[209] br[209] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_210 bl[210] br[210] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_211 bl[211] br[211] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_212 bl[212] br[212] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_213 bl[213] br[213] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_214 bl[214] br[214] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_215 bl[215] br[215] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_216 bl[216] br[216] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_217 bl[217] br[217] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_218 bl[218] br[218] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_219 bl[219] br[219] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_220 bl[220] br[220] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_221 bl[221] br[221] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_222 bl[222] br[222] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_223 bl[223] br[223] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_224 bl[224] br[224] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_225 bl[225] br[225] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_226 bl[226] br[226] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_227 bl[227] br[227] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_228 bl[228] br[228] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_229 bl[229] br[229] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_230 bl[230] br[230] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_231 bl[231] br[231] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_232 bl[232] br[232] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_233 bl[233] br[233] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_234 bl[234] br[234] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_235 bl[235] br[235] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_236 bl[236] br[236] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_237 bl[237] br[237] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_238 bl[238] br[238] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_239 bl[239] br[239] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_240 bl[240] br[240] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_241 bl[241] br[241] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_242 bl[242] br[242] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_243 bl[243] br[243] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_244 bl[244] br[244] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_245 bl[245] br[245] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_246 bl[246] br[246] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_247 bl[247] br[247] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_248 bl[248] br[248] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_249 bl[249] br[249] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_250 bl[250] br[250] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_251 bl[251] br[251] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_252 bl[252] br[252] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_253 bl[253] br[253] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_254 bl[254] br[254] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_255 bl[255] br[255] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_10_0 bl[0] br[0] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_1 bl[1] br[1] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_2 bl[2] br[2] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_3 bl[3] br[3] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_4 bl[4] br[4] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_5 bl[5] br[5] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_6 bl[6] br[6] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_7 bl[7] br[7] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_8 bl[8] br[8] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_9 bl[9] br[9] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_10 bl[10] br[10] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_11 bl[11] br[11] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_12 bl[12] br[12] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_13 bl[13] br[13] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_14 bl[14] br[14] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_15 bl[15] br[15] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_16 bl[16] br[16] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_17 bl[17] br[17] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_18 bl[18] br[18] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_19 bl[19] br[19] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_20 bl[20] br[20] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_21 bl[21] br[21] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_22 bl[22] br[22] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_23 bl[23] br[23] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_24 bl[24] br[24] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_25 bl[25] br[25] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_26 bl[26] br[26] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_27 bl[27] br[27] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_28 bl[28] br[28] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_29 bl[29] br[29] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_30 bl[30] br[30] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_31 bl[31] br[31] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_32 bl[32] br[32] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_33 bl[33] br[33] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_34 bl[34] br[34] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_35 bl[35] br[35] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_36 bl[36] br[36] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_37 bl[37] br[37] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_38 bl[38] br[38] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_39 bl[39] br[39] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_40 bl[40] br[40] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_41 bl[41] br[41] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_42 bl[42] br[42] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_43 bl[43] br[43] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_44 bl[44] br[44] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_45 bl[45] br[45] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_46 bl[46] br[46] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_47 bl[47] br[47] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_48 bl[48] br[48] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_49 bl[49] br[49] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_50 bl[50] br[50] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_51 bl[51] br[51] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_52 bl[52] br[52] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_53 bl[53] br[53] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_54 bl[54] br[54] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_55 bl[55] br[55] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_56 bl[56] br[56] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_57 bl[57] br[57] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_58 bl[58] br[58] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_59 bl[59] br[59] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_60 bl[60] br[60] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_61 bl[61] br[61] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_62 bl[62] br[62] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_63 bl[63] br[63] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_64 bl[64] br[64] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_65 bl[65] br[65] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_66 bl[66] br[66] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_67 bl[67] br[67] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_68 bl[68] br[68] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_69 bl[69] br[69] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_70 bl[70] br[70] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_71 bl[71] br[71] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_72 bl[72] br[72] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_73 bl[73] br[73] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_74 bl[74] br[74] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_75 bl[75] br[75] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_76 bl[76] br[76] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_77 bl[77] br[77] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_78 bl[78] br[78] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_79 bl[79] br[79] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_80 bl[80] br[80] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_81 bl[81] br[81] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_82 bl[82] br[82] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_83 bl[83] br[83] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_84 bl[84] br[84] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_85 bl[85] br[85] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_86 bl[86] br[86] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_87 bl[87] br[87] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_88 bl[88] br[88] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_89 bl[89] br[89] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_90 bl[90] br[90] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_91 bl[91] br[91] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_92 bl[92] br[92] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_93 bl[93] br[93] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_94 bl[94] br[94] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_95 bl[95] br[95] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_96 bl[96] br[96] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_97 bl[97] br[97] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_98 bl[98] br[98] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_99 bl[99] br[99] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_100 bl[100] br[100] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_101 bl[101] br[101] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_102 bl[102] br[102] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_103 bl[103] br[103] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_104 bl[104] br[104] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_105 bl[105] br[105] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_106 bl[106] br[106] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_107 bl[107] br[107] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_108 bl[108] br[108] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_109 bl[109] br[109] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_110 bl[110] br[110] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_111 bl[111] br[111] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_112 bl[112] br[112] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_113 bl[113] br[113] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_114 bl[114] br[114] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_115 bl[115] br[115] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_116 bl[116] br[116] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_117 bl[117] br[117] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_118 bl[118] br[118] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_119 bl[119] br[119] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_120 bl[120] br[120] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_121 bl[121] br[121] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_122 bl[122] br[122] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_123 bl[123] br[123] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_124 bl[124] br[124] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_125 bl[125] br[125] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_126 bl[126] br[126] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_127 bl[127] br[127] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_128 bl[128] br[128] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_129 bl[129] br[129] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_130 bl[130] br[130] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_131 bl[131] br[131] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_132 bl[132] br[132] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_133 bl[133] br[133] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_134 bl[134] br[134] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_135 bl[135] br[135] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_136 bl[136] br[136] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_137 bl[137] br[137] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_138 bl[138] br[138] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_139 bl[139] br[139] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_140 bl[140] br[140] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_141 bl[141] br[141] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_142 bl[142] br[142] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_143 bl[143] br[143] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_144 bl[144] br[144] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_145 bl[145] br[145] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_146 bl[146] br[146] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_147 bl[147] br[147] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_148 bl[148] br[148] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_149 bl[149] br[149] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_150 bl[150] br[150] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_151 bl[151] br[151] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_152 bl[152] br[152] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_153 bl[153] br[153] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_154 bl[154] br[154] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_155 bl[155] br[155] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_156 bl[156] br[156] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_157 bl[157] br[157] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_158 bl[158] br[158] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_159 bl[159] br[159] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_160 bl[160] br[160] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_161 bl[161] br[161] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_162 bl[162] br[162] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_163 bl[163] br[163] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_164 bl[164] br[164] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_165 bl[165] br[165] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_166 bl[166] br[166] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_167 bl[167] br[167] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_168 bl[168] br[168] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_169 bl[169] br[169] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_170 bl[170] br[170] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_171 bl[171] br[171] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_172 bl[172] br[172] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_173 bl[173] br[173] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_174 bl[174] br[174] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_175 bl[175] br[175] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_176 bl[176] br[176] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_177 bl[177] br[177] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_178 bl[178] br[178] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_179 bl[179] br[179] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_180 bl[180] br[180] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_181 bl[181] br[181] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_182 bl[182] br[182] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_183 bl[183] br[183] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_184 bl[184] br[184] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_185 bl[185] br[185] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_186 bl[186] br[186] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_187 bl[187] br[187] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_188 bl[188] br[188] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_189 bl[189] br[189] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_190 bl[190] br[190] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_191 bl[191] br[191] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_192 bl[192] br[192] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_193 bl[193] br[193] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_194 bl[194] br[194] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_195 bl[195] br[195] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_196 bl[196] br[196] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_197 bl[197] br[197] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_198 bl[198] br[198] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_199 bl[199] br[199] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_200 bl[200] br[200] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_201 bl[201] br[201] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_202 bl[202] br[202] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_203 bl[203] br[203] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_204 bl[204] br[204] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_205 bl[205] br[205] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_206 bl[206] br[206] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_207 bl[207] br[207] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_208 bl[208] br[208] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_209 bl[209] br[209] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_210 bl[210] br[210] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_211 bl[211] br[211] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_212 bl[212] br[212] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_213 bl[213] br[213] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_214 bl[214] br[214] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_215 bl[215] br[215] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_216 bl[216] br[216] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_217 bl[217] br[217] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_218 bl[218] br[218] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_219 bl[219] br[219] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_220 bl[220] br[220] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_221 bl[221] br[221] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_222 bl[222] br[222] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_223 bl[223] br[223] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_224 bl[224] br[224] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_225 bl[225] br[225] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_226 bl[226] br[226] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_227 bl[227] br[227] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_228 bl[228] br[228] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_229 bl[229] br[229] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_230 bl[230] br[230] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_231 bl[231] br[231] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_232 bl[232] br[232] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_233 bl[233] br[233] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_234 bl[234] br[234] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_235 bl[235] br[235] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_236 bl[236] br[236] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_237 bl[237] br[237] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_238 bl[238] br[238] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_239 bl[239] br[239] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_240 bl[240] br[240] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_241 bl[241] br[241] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_242 bl[242] br[242] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_243 bl[243] br[243] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_244 bl[244] br[244] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_245 bl[245] br[245] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_246 bl[246] br[246] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_247 bl[247] br[247] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_248 bl[248] br[248] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_249 bl[249] br[249] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_250 bl[250] br[250] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_251 bl[251] br[251] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_252 bl[252] br[252] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_253 bl[253] br[253] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_254 bl[254] br[254] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_255 bl[255] br[255] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_11_0 bl[0] br[0] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_1 bl[1] br[1] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_2 bl[2] br[2] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_3 bl[3] br[3] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_4 bl[4] br[4] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_5 bl[5] br[5] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_6 bl[6] br[6] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_7 bl[7] br[7] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_8 bl[8] br[8] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_9 bl[9] br[9] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_10 bl[10] br[10] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_11 bl[11] br[11] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_12 bl[12] br[12] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_13 bl[13] br[13] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_14 bl[14] br[14] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_15 bl[15] br[15] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_16 bl[16] br[16] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_17 bl[17] br[17] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_18 bl[18] br[18] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_19 bl[19] br[19] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_20 bl[20] br[20] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_21 bl[21] br[21] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_22 bl[22] br[22] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_23 bl[23] br[23] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_24 bl[24] br[24] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_25 bl[25] br[25] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_26 bl[26] br[26] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_27 bl[27] br[27] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_28 bl[28] br[28] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_29 bl[29] br[29] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_30 bl[30] br[30] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_31 bl[31] br[31] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_32 bl[32] br[32] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_33 bl[33] br[33] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_34 bl[34] br[34] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_35 bl[35] br[35] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_36 bl[36] br[36] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_37 bl[37] br[37] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_38 bl[38] br[38] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_39 bl[39] br[39] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_40 bl[40] br[40] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_41 bl[41] br[41] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_42 bl[42] br[42] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_43 bl[43] br[43] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_44 bl[44] br[44] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_45 bl[45] br[45] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_46 bl[46] br[46] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_47 bl[47] br[47] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_48 bl[48] br[48] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_49 bl[49] br[49] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_50 bl[50] br[50] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_51 bl[51] br[51] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_52 bl[52] br[52] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_53 bl[53] br[53] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_54 bl[54] br[54] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_55 bl[55] br[55] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_56 bl[56] br[56] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_57 bl[57] br[57] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_58 bl[58] br[58] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_59 bl[59] br[59] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_60 bl[60] br[60] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_61 bl[61] br[61] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_62 bl[62] br[62] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_63 bl[63] br[63] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_64 bl[64] br[64] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_65 bl[65] br[65] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_66 bl[66] br[66] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_67 bl[67] br[67] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_68 bl[68] br[68] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_69 bl[69] br[69] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_70 bl[70] br[70] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_71 bl[71] br[71] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_72 bl[72] br[72] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_73 bl[73] br[73] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_74 bl[74] br[74] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_75 bl[75] br[75] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_76 bl[76] br[76] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_77 bl[77] br[77] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_78 bl[78] br[78] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_79 bl[79] br[79] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_80 bl[80] br[80] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_81 bl[81] br[81] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_82 bl[82] br[82] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_83 bl[83] br[83] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_84 bl[84] br[84] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_85 bl[85] br[85] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_86 bl[86] br[86] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_87 bl[87] br[87] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_88 bl[88] br[88] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_89 bl[89] br[89] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_90 bl[90] br[90] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_91 bl[91] br[91] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_92 bl[92] br[92] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_93 bl[93] br[93] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_94 bl[94] br[94] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_95 bl[95] br[95] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_96 bl[96] br[96] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_97 bl[97] br[97] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_98 bl[98] br[98] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_99 bl[99] br[99] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_100 bl[100] br[100] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_101 bl[101] br[101] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_102 bl[102] br[102] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_103 bl[103] br[103] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_104 bl[104] br[104] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_105 bl[105] br[105] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_106 bl[106] br[106] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_107 bl[107] br[107] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_108 bl[108] br[108] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_109 bl[109] br[109] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_110 bl[110] br[110] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_111 bl[111] br[111] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_112 bl[112] br[112] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_113 bl[113] br[113] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_114 bl[114] br[114] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_115 bl[115] br[115] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_116 bl[116] br[116] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_117 bl[117] br[117] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_118 bl[118] br[118] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_119 bl[119] br[119] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_120 bl[120] br[120] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_121 bl[121] br[121] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_122 bl[122] br[122] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_123 bl[123] br[123] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_124 bl[124] br[124] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_125 bl[125] br[125] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_126 bl[126] br[126] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_127 bl[127] br[127] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_128 bl[128] br[128] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_129 bl[129] br[129] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_130 bl[130] br[130] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_131 bl[131] br[131] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_132 bl[132] br[132] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_133 bl[133] br[133] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_134 bl[134] br[134] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_135 bl[135] br[135] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_136 bl[136] br[136] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_137 bl[137] br[137] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_138 bl[138] br[138] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_139 bl[139] br[139] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_140 bl[140] br[140] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_141 bl[141] br[141] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_142 bl[142] br[142] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_143 bl[143] br[143] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_144 bl[144] br[144] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_145 bl[145] br[145] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_146 bl[146] br[146] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_147 bl[147] br[147] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_148 bl[148] br[148] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_149 bl[149] br[149] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_150 bl[150] br[150] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_151 bl[151] br[151] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_152 bl[152] br[152] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_153 bl[153] br[153] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_154 bl[154] br[154] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_155 bl[155] br[155] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_156 bl[156] br[156] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_157 bl[157] br[157] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_158 bl[158] br[158] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_159 bl[159] br[159] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_160 bl[160] br[160] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_161 bl[161] br[161] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_162 bl[162] br[162] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_163 bl[163] br[163] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_164 bl[164] br[164] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_165 bl[165] br[165] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_166 bl[166] br[166] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_167 bl[167] br[167] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_168 bl[168] br[168] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_169 bl[169] br[169] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_170 bl[170] br[170] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_171 bl[171] br[171] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_172 bl[172] br[172] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_173 bl[173] br[173] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_174 bl[174] br[174] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_175 bl[175] br[175] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_176 bl[176] br[176] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_177 bl[177] br[177] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_178 bl[178] br[178] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_179 bl[179] br[179] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_180 bl[180] br[180] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_181 bl[181] br[181] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_182 bl[182] br[182] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_183 bl[183] br[183] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_184 bl[184] br[184] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_185 bl[185] br[185] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_186 bl[186] br[186] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_187 bl[187] br[187] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_188 bl[188] br[188] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_189 bl[189] br[189] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_190 bl[190] br[190] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_191 bl[191] br[191] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_192 bl[192] br[192] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_193 bl[193] br[193] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_194 bl[194] br[194] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_195 bl[195] br[195] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_196 bl[196] br[196] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_197 bl[197] br[197] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_198 bl[198] br[198] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_199 bl[199] br[199] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_200 bl[200] br[200] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_201 bl[201] br[201] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_202 bl[202] br[202] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_203 bl[203] br[203] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_204 bl[204] br[204] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_205 bl[205] br[205] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_206 bl[206] br[206] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_207 bl[207] br[207] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_208 bl[208] br[208] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_209 bl[209] br[209] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_210 bl[210] br[210] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_211 bl[211] br[211] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_212 bl[212] br[212] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_213 bl[213] br[213] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_214 bl[214] br[214] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_215 bl[215] br[215] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_216 bl[216] br[216] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_217 bl[217] br[217] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_218 bl[218] br[218] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_219 bl[219] br[219] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_220 bl[220] br[220] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_221 bl[221] br[221] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_222 bl[222] br[222] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_223 bl[223] br[223] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_224 bl[224] br[224] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_225 bl[225] br[225] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_226 bl[226] br[226] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_227 bl[227] br[227] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_228 bl[228] br[228] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_229 bl[229] br[229] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_230 bl[230] br[230] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_231 bl[231] br[231] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_232 bl[232] br[232] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_233 bl[233] br[233] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_234 bl[234] br[234] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_235 bl[235] br[235] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_236 bl[236] br[236] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_237 bl[237] br[237] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_238 bl[238] br[238] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_239 bl[239] br[239] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_240 bl[240] br[240] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_241 bl[241] br[241] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_242 bl[242] br[242] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_243 bl[243] br[243] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_244 bl[244] br[244] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_245 bl[245] br[245] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_246 bl[246] br[246] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_247 bl[247] br[247] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_248 bl[248] br[248] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_249 bl[249] br[249] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_250 bl[250] br[250] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_251 bl[251] br[251] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_252 bl[252] br[252] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_253 bl[253] br[253] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_254 bl[254] br[254] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_255 bl[255] br[255] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_12_0 bl[0] br[0] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_1 bl[1] br[1] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_2 bl[2] br[2] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_3 bl[3] br[3] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_4 bl[4] br[4] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_5 bl[5] br[5] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_6 bl[6] br[6] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_7 bl[7] br[7] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_8 bl[8] br[8] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_9 bl[9] br[9] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_10 bl[10] br[10] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_11 bl[11] br[11] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_12 bl[12] br[12] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_13 bl[13] br[13] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_14 bl[14] br[14] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_15 bl[15] br[15] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_16 bl[16] br[16] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_17 bl[17] br[17] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_18 bl[18] br[18] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_19 bl[19] br[19] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_20 bl[20] br[20] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_21 bl[21] br[21] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_22 bl[22] br[22] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_23 bl[23] br[23] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_24 bl[24] br[24] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_25 bl[25] br[25] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_26 bl[26] br[26] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_27 bl[27] br[27] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_28 bl[28] br[28] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_29 bl[29] br[29] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_30 bl[30] br[30] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_31 bl[31] br[31] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_32 bl[32] br[32] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_33 bl[33] br[33] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_34 bl[34] br[34] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_35 bl[35] br[35] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_36 bl[36] br[36] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_37 bl[37] br[37] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_38 bl[38] br[38] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_39 bl[39] br[39] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_40 bl[40] br[40] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_41 bl[41] br[41] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_42 bl[42] br[42] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_43 bl[43] br[43] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_44 bl[44] br[44] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_45 bl[45] br[45] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_46 bl[46] br[46] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_47 bl[47] br[47] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_48 bl[48] br[48] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_49 bl[49] br[49] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_50 bl[50] br[50] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_51 bl[51] br[51] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_52 bl[52] br[52] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_53 bl[53] br[53] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_54 bl[54] br[54] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_55 bl[55] br[55] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_56 bl[56] br[56] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_57 bl[57] br[57] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_58 bl[58] br[58] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_59 bl[59] br[59] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_60 bl[60] br[60] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_61 bl[61] br[61] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_62 bl[62] br[62] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_63 bl[63] br[63] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_64 bl[64] br[64] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_65 bl[65] br[65] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_66 bl[66] br[66] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_67 bl[67] br[67] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_68 bl[68] br[68] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_69 bl[69] br[69] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_70 bl[70] br[70] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_71 bl[71] br[71] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_72 bl[72] br[72] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_73 bl[73] br[73] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_74 bl[74] br[74] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_75 bl[75] br[75] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_76 bl[76] br[76] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_77 bl[77] br[77] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_78 bl[78] br[78] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_79 bl[79] br[79] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_80 bl[80] br[80] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_81 bl[81] br[81] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_82 bl[82] br[82] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_83 bl[83] br[83] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_84 bl[84] br[84] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_85 bl[85] br[85] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_86 bl[86] br[86] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_87 bl[87] br[87] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_88 bl[88] br[88] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_89 bl[89] br[89] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_90 bl[90] br[90] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_91 bl[91] br[91] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_92 bl[92] br[92] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_93 bl[93] br[93] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_94 bl[94] br[94] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_95 bl[95] br[95] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_96 bl[96] br[96] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_97 bl[97] br[97] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_98 bl[98] br[98] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_99 bl[99] br[99] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_100 bl[100] br[100] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_101 bl[101] br[101] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_102 bl[102] br[102] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_103 bl[103] br[103] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_104 bl[104] br[104] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_105 bl[105] br[105] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_106 bl[106] br[106] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_107 bl[107] br[107] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_108 bl[108] br[108] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_109 bl[109] br[109] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_110 bl[110] br[110] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_111 bl[111] br[111] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_112 bl[112] br[112] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_113 bl[113] br[113] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_114 bl[114] br[114] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_115 bl[115] br[115] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_116 bl[116] br[116] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_117 bl[117] br[117] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_118 bl[118] br[118] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_119 bl[119] br[119] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_120 bl[120] br[120] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_121 bl[121] br[121] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_122 bl[122] br[122] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_123 bl[123] br[123] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_124 bl[124] br[124] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_125 bl[125] br[125] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_126 bl[126] br[126] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_127 bl[127] br[127] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_128 bl[128] br[128] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_129 bl[129] br[129] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_130 bl[130] br[130] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_131 bl[131] br[131] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_132 bl[132] br[132] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_133 bl[133] br[133] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_134 bl[134] br[134] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_135 bl[135] br[135] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_136 bl[136] br[136] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_137 bl[137] br[137] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_138 bl[138] br[138] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_139 bl[139] br[139] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_140 bl[140] br[140] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_141 bl[141] br[141] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_142 bl[142] br[142] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_143 bl[143] br[143] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_144 bl[144] br[144] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_145 bl[145] br[145] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_146 bl[146] br[146] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_147 bl[147] br[147] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_148 bl[148] br[148] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_149 bl[149] br[149] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_150 bl[150] br[150] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_151 bl[151] br[151] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_152 bl[152] br[152] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_153 bl[153] br[153] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_154 bl[154] br[154] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_155 bl[155] br[155] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_156 bl[156] br[156] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_157 bl[157] br[157] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_158 bl[158] br[158] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_159 bl[159] br[159] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_160 bl[160] br[160] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_161 bl[161] br[161] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_162 bl[162] br[162] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_163 bl[163] br[163] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_164 bl[164] br[164] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_165 bl[165] br[165] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_166 bl[166] br[166] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_167 bl[167] br[167] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_168 bl[168] br[168] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_169 bl[169] br[169] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_170 bl[170] br[170] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_171 bl[171] br[171] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_172 bl[172] br[172] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_173 bl[173] br[173] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_174 bl[174] br[174] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_175 bl[175] br[175] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_176 bl[176] br[176] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_177 bl[177] br[177] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_178 bl[178] br[178] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_179 bl[179] br[179] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_180 bl[180] br[180] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_181 bl[181] br[181] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_182 bl[182] br[182] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_183 bl[183] br[183] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_184 bl[184] br[184] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_185 bl[185] br[185] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_186 bl[186] br[186] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_187 bl[187] br[187] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_188 bl[188] br[188] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_189 bl[189] br[189] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_190 bl[190] br[190] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_191 bl[191] br[191] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_192 bl[192] br[192] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_193 bl[193] br[193] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_194 bl[194] br[194] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_195 bl[195] br[195] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_196 bl[196] br[196] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_197 bl[197] br[197] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_198 bl[198] br[198] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_199 bl[199] br[199] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_200 bl[200] br[200] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_201 bl[201] br[201] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_202 bl[202] br[202] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_203 bl[203] br[203] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_204 bl[204] br[204] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_205 bl[205] br[205] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_206 bl[206] br[206] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_207 bl[207] br[207] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_208 bl[208] br[208] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_209 bl[209] br[209] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_210 bl[210] br[210] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_211 bl[211] br[211] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_212 bl[212] br[212] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_213 bl[213] br[213] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_214 bl[214] br[214] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_215 bl[215] br[215] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_216 bl[216] br[216] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_217 bl[217] br[217] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_218 bl[218] br[218] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_219 bl[219] br[219] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_220 bl[220] br[220] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_221 bl[221] br[221] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_222 bl[222] br[222] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_223 bl[223] br[223] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_224 bl[224] br[224] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_225 bl[225] br[225] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_226 bl[226] br[226] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_227 bl[227] br[227] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_228 bl[228] br[228] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_229 bl[229] br[229] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_230 bl[230] br[230] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_231 bl[231] br[231] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_232 bl[232] br[232] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_233 bl[233] br[233] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_234 bl[234] br[234] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_235 bl[235] br[235] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_236 bl[236] br[236] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_237 bl[237] br[237] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_238 bl[238] br[238] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_239 bl[239] br[239] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_240 bl[240] br[240] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_241 bl[241] br[241] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_242 bl[242] br[242] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_243 bl[243] br[243] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_244 bl[244] br[244] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_245 bl[245] br[245] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_246 bl[246] br[246] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_247 bl[247] br[247] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_248 bl[248] br[248] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_249 bl[249] br[249] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_250 bl[250] br[250] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_251 bl[251] br[251] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_252 bl[252] br[252] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_253 bl[253] br[253] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_254 bl[254] br[254] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_255 bl[255] br[255] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_13_0 bl[0] br[0] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_1 bl[1] br[1] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_2 bl[2] br[2] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_3 bl[3] br[3] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_4 bl[4] br[4] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_5 bl[5] br[5] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_6 bl[6] br[6] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_7 bl[7] br[7] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_8 bl[8] br[8] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_9 bl[9] br[9] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_10 bl[10] br[10] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_11 bl[11] br[11] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_12 bl[12] br[12] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_13 bl[13] br[13] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_14 bl[14] br[14] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_15 bl[15] br[15] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_16 bl[16] br[16] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_17 bl[17] br[17] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_18 bl[18] br[18] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_19 bl[19] br[19] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_20 bl[20] br[20] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_21 bl[21] br[21] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_22 bl[22] br[22] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_23 bl[23] br[23] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_24 bl[24] br[24] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_25 bl[25] br[25] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_26 bl[26] br[26] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_27 bl[27] br[27] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_28 bl[28] br[28] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_29 bl[29] br[29] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_30 bl[30] br[30] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_31 bl[31] br[31] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_32 bl[32] br[32] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_33 bl[33] br[33] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_34 bl[34] br[34] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_35 bl[35] br[35] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_36 bl[36] br[36] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_37 bl[37] br[37] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_38 bl[38] br[38] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_39 bl[39] br[39] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_40 bl[40] br[40] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_41 bl[41] br[41] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_42 bl[42] br[42] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_43 bl[43] br[43] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_44 bl[44] br[44] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_45 bl[45] br[45] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_46 bl[46] br[46] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_47 bl[47] br[47] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_48 bl[48] br[48] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_49 bl[49] br[49] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_50 bl[50] br[50] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_51 bl[51] br[51] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_52 bl[52] br[52] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_53 bl[53] br[53] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_54 bl[54] br[54] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_55 bl[55] br[55] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_56 bl[56] br[56] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_57 bl[57] br[57] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_58 bl[58] br[58] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_59 bl[59] br[59] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_60 bl[60] br[60] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_61 bl[61] br[61] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_62 bl[62] br[62] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_63 bl[63] br[63] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_64 bl[64] br[64] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_65 bl[65] br[65] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_66 bl[66] br[66] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_67 bl[67] br[67] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_68 bl[68] br[68] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_69 bl[69] br[69] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_70 bl[70] br[70] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_71 bl[71] br[71] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_72 bl[72] br[72] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_73 bl[73] br[73] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_74 bl[74] br[74] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_75 bl[75] br[75] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_76 bl[76] br[76] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_77 bl[77] br[77] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_78 bl[78] br[78] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_79 bl[79] br[79] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_80 bl[80] br[80] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_81 bl[81] br[81] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_82 bl[82] br[82] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_83 bl[83] br[83] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_84 bl[84] br[84] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_85 bl[85] br[85] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_86 bl[86] br[86] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_87 bl[87] br[87] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_88 bl[88] br[88] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_89 bl[89] br[89] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_90 bl[90] br[90] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_91 bl[91] br[91] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_92 bl[92] br[92] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_93 bl[93] br[93] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_94 bl[94] br[94] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_95 bl[95] br[95] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_96 bl[96] br[96] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_97 bl[97] br[97] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_98 bl[98] br[98] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_99 bl[99] br[99] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_100 bl[100] br[100] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_101 bl[101] br[101] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_102 bl[102] br[102] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_103 bl[103] br[103] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_104 bl[104] br[104] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_105 bl[105] br[105] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_106 bl[106] br[106] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_107 bl[107] br[107] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_108 bl[108] br[108] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_109 bl[109] br[109] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_110 bl[110] br[110] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_111 bl[111] br[111] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_112 bl[112] br[112] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_113 bl[113] br[113] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_114 bl[114] br[114] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_115 bl[115] br[115] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_116 bl[116] br[116] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_117 bl[117] br[117] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_118 bl[118] br[118] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_119 bl[119] br[119] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_120 bl[120] br[120] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_121 bl[121] br[121] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_122 bl[122] br[122] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_123 bl[123] br[123] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_124 bl[124] br[124] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_125 bl[125] br[125] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_126 bl[126] br[126] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_127 bl[127] br[127] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_128 bl[128] br[128] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_129 bl[129] br[129] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_130 bl[130] br[130] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_131 bl[131] br[131] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_132 bl[132] br[132] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_133 bl[133] br[133] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_134 bl[134] br[134] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_135 bl[135] br[135] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_136 bl[136] br[136] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_137 bl[137] br[137] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_138 bl[138] br[138] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_139 bl[139] br[139] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_140 bl[140] br[140] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_141 bl[141] br[141] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_142 bl[142] br[142] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_143 bl[143] br[143] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_144 bl[144] br[144] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_145 bl[145] br[145] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_146 bl[146] br[146] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_147 bl[147] br[147] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_148 bl[148] br[148] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_149 bl[149] br[149] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_150 bl[150] br[150] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_151 bl[151] br[151] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_152 bl[152] br[152] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_153 bl[153] br[153] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_154 bl[154] br[154] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_155 bl[155] br[155] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_156 bl[156] br[156] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_157 bl[157] br[157] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_158 bl[158] br[158] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_159 bl[159] br[159] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_160 bl[160] br[160] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_161 bl[161] br[161] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_162 bl[162] br[162] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_163 bl[163] br[163] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_164 bl[164] br[164] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_165 bl[165] br[165] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_166 bl[166] br[166] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_167 bl[167] br[167] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_168 bl[168] br[168] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_169 bl[169] br[169] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_170 bl[170] br[170] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_171 bl[171] br[171] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_172 bl[172] br[172] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_173 bl[173] br[173] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_174 bl[174] br[174] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_175 bl[175] br[175] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_176 bl[176] br[176] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_177 bl[177] br[177] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_178 bl[178] br[178] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_179 bl[179] br[179] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_180 bl[180] br[180] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_181 bl[181] br[181] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_182 bl[182] br[182] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_183 bl[183] br[183] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_184 bl[184] br[184] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_185 bl[185] br[185] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_186 bl[186] br[186] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_187 bl[187] br[187] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_188 bl[188] br[188] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_189 bl[189] br[189] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_190 bl[190] br[190] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_191 bl[191] br[191] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_192 bl[192] br[192] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_193 bl[193] br[193] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_194 bl[194] br[194] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_195 bl[195] br[195] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_196 bl[196] br[196] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_197 bl[197] br[197] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_198 bl[198] br[198] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_199 bl[199] br[199] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_200 bl[200] br[200] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_201 bl[201] br[201] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_202 bl[202] br[202] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_203 bl[203] br[203] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_204 bl[204] br[204] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_205 bl[205] br[205] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_206 bl[206] br[206] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_207 bl[207] br[207] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_208 bl[208] br[208] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_209 bl[209] br[209] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_210 bl[210] br[210] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_211 bl[211] br[211] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_212 bl[212] br[212] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_213 bl[213] br[213] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_214 bl[214] br[214] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_215 bl[215] br[215] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_216 bl[216] br[216] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_217 bl[217] br[217] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_218 bl[218] br[218] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_219 bl[219] br[219] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_220 bl[220] br[220] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_221 bl[221] br[221] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_222 bl[222] br[222] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_223 bl[223] br[223] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_224 bl[224] br[224] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_225 bl[225] br[225] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_226 bl[226] br[226] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_227 bl[227] br[227] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_228 bl[228] br[228] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_229 bl[229] br[229] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_230 bl[230] br[230] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_231 bl[231] br[231] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_232 bl[232] br[232] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_233 bl[233] br[233] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_234 bl[234] br[234] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_235 bl[235] br[235] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_236 bl[236] br[236] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_237 bl[237] br[237] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_238 bl[238] br[238] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_239 bl[239] br[239] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_240 bl[240] br[240] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_241 bl[241] br[241] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_242 bl[242] br[242] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_243 bl[243] br[243] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_244 bl[244] br[244] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_245 bl[245] br[245] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_246 bl[246] br[246] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_247 bl[247] br[247] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_248 bl[248] br[248] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_249 bl[249] br[249] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_250 bl[250] br[250] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_251 bl[251] br[251] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_252 bl[252] br[252] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_253 bl[253] br[253] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_254 bl[254] br[254] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_255 bl[255] br[255] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_14_0 bl[0] br[0] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_1 bl[1] br[1] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_2 bl[2] br[2] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_3 bl[3] br[3] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_4 bl[4] br[4] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_5 bl[5] br[5] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_6 bl[6] br[6] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_7 bl[7] br[7] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_8 bl[8] br[8] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_9 bl[9] br[9] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_10 bl[10] br[10] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_11 bl[11] br[11] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_12 bl[12] br[12] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_13 bl[13] br[13] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_14 bl[14] br[14] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_15 bl[15] br[15] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_16 bl[16] br[16] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_17 bl[17] br[17] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_18 bl[18] br[18] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_19 bl[19] br[19] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_20 bl[20] br[20] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_21 bl[21] br[21] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_22 bl[22] br[22] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_23 bl[23] br[23] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_24 bl[24] br[24] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_25 bl[25] br[25] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_26 bl[26] br[26] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_27 bl[27] br[27] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_28 bl[28] br[28] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_29 bl[29] br[29] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_30 bl[30] br[30] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_31 bl[31] br[31] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_32 bl[32] br[32] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_33 bl[33] br[33] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_34 bl[34] br[34] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_35 bl[35] br[35] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_36 bl[36] br[36] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_37 bl[37] br[37] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_38 bl[38] br[38] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_39 bl[39] br[39] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_40 bl[40] br[40] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_41 bl[41] br[41] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_42 bl[42] br[42] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_43 bl[43] br[43] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_44 bl[44] br[44] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_45 bl[45] br[45] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_46 bl[46] br[46] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_47 bl[47] br[47] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_48 bl[48] br[48] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_49 bl[49] br[49] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_50 bl[50] br[50] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_51 bl[51] br[51] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_52 bl[52] br[52] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_53 bl[53] br[53] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_54 bl[54] br[54] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_55 bl[55] br[55] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_56 bl[56] br[56] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_57 bl[57] br[57] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_58 bl[58] br[58] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_59 bl[59] br[59] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_60 bl[60] br[60] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_61 bl[61] br[61] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_62 bl[62] br[62] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_63 bl[63] br[63] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_64 bl[64] br[64] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_65 bl[65] br[65] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_66 bl[66] br[66] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_67 bl[67] br[67] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_68 bl[68] br[68] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_69 bl[69] br[69] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_70 bl[70] br[70] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_71 bl[71] br[71] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_72 bl[72] br[72] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_73 bl[73] br[73] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_74 bl[74] br[74] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_75 bl[75] br[75] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_76 bl[76] br[76] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_77 bl[77] br[77] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_78 bl[78] br[78] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_79 bl[79] br[79] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_80 bl[80] br[80] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_81 bl[81] br[81] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_82 bl[82] br[82] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_83 bl[83] br[83] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_84 bl[84] br[84] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_85 bl[85] br[85] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_86 bl[86] br[86] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_87 bl[87] br[87] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_88 bl[88] br[88] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_89 bl[89] br[89] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_90 bl[90] br[90] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_91 bl[91] br[91] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_92 bl[92] br[92] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_93 bl[93] br[93] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_94 bl[94] br[94] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_95 bl[95] br[95] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_96 bl[96] br[96] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_97 bl[97] br[97] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_98 bl[98] br[98] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_99 bl[99] br[99] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_100 bl[100] br[100] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_101 bl[101] br[101] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_102 bl[102] br[102] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_103 bl[103] br[103] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_104 bl[104] br[104] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_105 bl[105] br[105] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_106 bl[106] br[106] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_107 bl[107] br[107] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_108 bl[108] br[108] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_109 bl[109] br[109] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_110 bl[110] br[110] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_111 bl[111] br[111] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_112 bl[112] br[112] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_113 bl[113] br[113] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_114 bl[114] br[114] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_115 bl[115] br[115] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_116 bl[116] br[116] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_117 bl[117] br[117] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_118 bl[118] br[118] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_119 bl[119] br[119] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_120 bl[120] br[120] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_121 bl[121] br[121] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_122 bl[122] br[122] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_123 bl[123] br[123] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_124 bl[124] br[124] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_125 bl[125] br[125] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_126 bl[126] br[126] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_127 bl[127] br[127] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_128 bl[128] br[128] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_129 bl[129] br[129] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_130 bl[130] br[130] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_131 bl[131] br[131] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_132 bl[132] br[132] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_133 bl[133] br[133] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_134 bl[134] br[134] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_135 bl[135] br[135] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_136 bl[136] br[136] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_137 bl[137] br[137] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_138 bl[138] br[138] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_139 bl[139] br[139] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_140 bl[140] br[140] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_141 bl[141] br[141] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_142 bl[142] br[142] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_143 bl[143] br[143] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_144 bl[144] br[144] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_145 bl[145] br[145] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_146 bl[146] br[146] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_147 bl[147] br[147] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_148 bl[148] br[148] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_149 bl[149] br[149] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_150 bl[150] br[150] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_151 bl[151] br[151] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_152 bl[152] br[152] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_153 bl[153] br[153] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_154 bl[154] br[154] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_155 bl[155] br[155] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_156 bl[156] br[156] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_157 bl[157] br[157] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_158 bl[158] br[158] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_159 bl[159] br[159] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_160 bl[160] br[160] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_161 bl[161] br[161] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_162 bl[162] br[162] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_163 bl[163] br[163] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_164 bl[164] br[164] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_165 bl[165] br[165] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_166 bl[166] br[166] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_167 bl[167] br[167] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_168 bl[168] br[168] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_169 bl[169] br[169] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_170 bl[170] br[170] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_171 bl[171] br[171] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_172 bl[172] br[172] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_173 bl[173] br[173] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_174 bl[174] br[174] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_175 bl[175] br[175] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_176 bl[176] br[176] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_177 bl[177] br[177] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_178 bl[178] br[178] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_179 bl[179] br[179] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_180 bl[180] br[180] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_181 bl[181] br[181] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_182 bl[182] br[182] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_183 bl[183] br[183] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_184 bl[184] br[184] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_185 bl[185] br[185] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_186 bl[186] br[186] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_187 bl[187] br[187] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_188 bl[188] br[188] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_189 bl[189] br[189] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_190 bl[190] br[190] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_191 bl[191] br[191] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_192 bl[192] br[192] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_193 bl[193] br[193] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_194 bl[194] br[194] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_195 bl[195] br[195] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_196 bl[196] br[196] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_197 bl[197] br[197] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_198 bl[198] br[198] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_199 bl[199] br[199] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_200 bl[200] br[200] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_201 bl[201] br[201] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_202 bl[202] br[202] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_203 bl[203] br[203] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_204 bl[204] br[204] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_205 bl[205] br[205] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_206 bl[206] br[206] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_207 bl[207] br[207] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_208 bl[208] br[208] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_209 bl[209] br[209] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_210 bl[210] br[210] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_211 bl[211] br[211] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_212 bl[212] br[212] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_213 bl[213] br[213] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_214 bl[214] br[214] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_215 bl[215] br[215] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_216 bl[216] br[216] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_217 bl[217] br[217] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_218 bl[218] br[218] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_219 bl[219] br[219] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_220 bl[220] br[220] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_221 bl[221] br[221] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_222 bl[222] br[222] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_223 bl[223] br[223] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_224 bl[224] br[224] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_225 bl[225] br[225] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_226 bl[226] br[226] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_227 bl[227] br[227] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_228 bl[228] br[228] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_229 bl[229] br[229] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_230 bl[230] br[230] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_231 bl[231] br[231] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_232 bl[232] br[232] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_233 bl[233] br[233] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_234 bl[234] br[234] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_235 bl[235] br[235] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_236 bl[236] br[236] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_237 bl[237] br[237] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_238 bl[238] br[238] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_239 bl[239] br[239] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_240 bl[240] br[240] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_241 bl[241] br[241] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_242 bl[242] br[242] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_243 bl[243] br[243] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_244 bl[244] br[244] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_245 bl[245] br[245] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_246 bl[246] br[246] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_247 bl[247] br[247] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_248 bl[248] br[248] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_249 bl[249] br[249] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_250 bl[250] br[250] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_251 bl[251] br[251] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_252 bl[252] br[252] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_253 bl[253] br[253] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_254 bl[254] br[254] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_255 bl[255] br[255] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_15_0 bl[0] br[0] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_1 bl[1] br[1] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_2 bl[2] br[2] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_3 bl[3] br[3] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_4 bl[4] br[4] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_5 bl[5] br[5] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_6 bl[6] br[6] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_7 bl[7] br[7] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_8 bl[8] br[8] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_9 bl[9] br[9] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_10 bl[10] br[10] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_11 bl[11] br[11] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_12 bl[12] br[12] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_13 bl[13] br[13] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_14 bl[14] br[14] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_15 bl[15] br[15] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_16 bl[16] br[16] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_17 bl[17] br[17] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_18 bl[18] br[18] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_19 bl[19] br[19] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_20 bl[20] br[20] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_21 bl[21] br[21] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_22 bl[22] br[22] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_23 bl[23] br[23] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_24 bl[24] br[24] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_25 bl[25] br[25] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_26 bl[26] br[26] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_27 bl[27] br[27] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_28 bl[28] br[28] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_29 bl[29] br[29] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_30 bl[30] br[30] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_31 bl[31] br[31] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_32 bl[32] br[32] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_33 bl[33] br[33] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_34 bl[34] br[34] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_35 bl[35] br[35] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_36 bl[36] br[36] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_37 bl[37] br[37] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_38 bl[38] br[38] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_39 bl[39] br[39] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_40 bl[40] br[40] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_41 bl[41] br[41] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_42 bl[42] br[42] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_43 bl[43] br[43] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_44 bl[44] br[44] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_45 bl[45] br[45] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_46 bl[46] br[46] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_47 bl[47] br[47] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_48 bl[48] br[48] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_49 bl[49] br[49] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_50 bl[50] br[50] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_51 bl[51] br[51] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_52 bl[52] br[52] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_53 bl[53] br[53] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_54 bl[54] br[54] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_55 bl[55] br[55] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_56 bl[56] br[56] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_57 bl[57] br[57] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_58 bl[58] br[58] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_59 bl[59] br[59] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_60 bl[60] br[60] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_61 bl[61] br[61] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_62 bl[62] br[62] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_63 bl[63] br[63] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_64 bl[64] br[64] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_65 bl[65] br[65] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_66 bl[66] br[66] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_67 bl[67] br[67] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_68 bl[68] br[68] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_69 bl[69] br[69] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_70 bl[70] br[70] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_71 bl[71] br[71] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_72 bl[72] br[72] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_73 bl[73] br[73] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_74 bl[74] br[74] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_75 bl[75] br[75] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_76 bl[76] br[76] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_77 bl[77] br[77] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_78 bl[78] br[78] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_79 bl[79] br[79] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_80 bl[80] br[80] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_81 bl[81] br[81] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_82 bl[82] br[82] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_83 bl[83] br[83] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_84 bl[84] br[84] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_85 bl[85] br[85] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_86 bl[86] br[86] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_87 bl[87] br[87] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_88 bl[88] br[88] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_89 bl[89] br[89] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_90 bl[90] br[90] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_91 bl[91] br[91] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_92 bl[92] br[92] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_93 bl[93] br[93] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_94 bl[94] br[94] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_95 bl[95] br[95] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_96 bl[96] br[96] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_97 bl[97] br[97] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_98 bl[98] br[98] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_99 bl[99] br[99] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_100 bl[100] br[100] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_101 bl[101] br[101] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_102 bl[102] br[102] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_103 bl[103] br[103] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_104 bl[104] br[104] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_105 bl[105] br[105] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_106 bl[106] br[106] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_107 bl[107] br[107] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_108 bl[108] br[108] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_109 bl[109] br[109] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_110 bl[110] br[110] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_111 bl[111] br[111] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_112 bl[112] br[112] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_113 bl[113] br[113] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_114 bl[114] br[114] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_115 bl[115] br[115] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_116 bl[116] br[116] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_117 bl[117] br[117] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_118 bl[118] br[118] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_119 bl[119] br[119] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_120 bl[120] br[120] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_121 bl[121] br[121] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_122 bl[122] br[122] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_123 bl[123] br[123] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_124 bl[124] br[124] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_125 bl[125] br[125] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_126 bl[126] br[126] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_127 bl[127] br[127] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_128 bl[128] br[128] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_129 bl[129] br[129] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_130 bl[130] br[130] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_131 bl[131] br[131] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_132 bl[132] br[132] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_133 bl[133] br[133] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_134 bl[134] br[134] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_135 bl[135] br[135] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_136 bl[136] br[136] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_137 bl[137] br[137] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_138 bl[138] br[138] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_139 bl[139] br[139] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_140 bl[140] br[140] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_141 bl[141] br[141] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_142 bl[142] br[142] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_143 bl[143] br[143] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_144 bl[144] br[144] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_145 bl[145] br[145] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_146 bl[146] br[146] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_147 bl[147] br[147] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_148 bl[148] br[148] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_149 bl[149] br[149] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_150 bl[150] br[150] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_151 bl[151] br[151] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_152 bl[152] br[152] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_153 bl[153] br[153] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_154 bl[154] br[154] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_155 bl[155] br[155] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_156 bl[156] br[156] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_157 bl[157] br[157] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_158 bl[158] br[158] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_159 bl[159] br[159] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_160 bl[160] br[160] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_161 bl[161] br[161] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_162 bl[162] br[162] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_163 bl[163] br[163] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_164 bl[164] br[164] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_165 bl[165] br[165] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_166 bl[166] br[166] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_167 bl[167] br[167] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_168 bl[168] br[168] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_169 bl[169] br[169] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_170 bl[170] br[170] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_171 bl[171] br[171] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_172 bl[172] br[172] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_173 bl[173] br[173] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_174 bl[174] br[174] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_175 bl[175] br[175] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_176 bl[176] br[176] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_177 bl[177] br[177] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_178 bl[178] br[178] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_179 bl[179] br[179] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_180 bl[180] br[180] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_181 bl[181] br[181] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_182 bl[182] br[182] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_183 bl[183] br[183] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_184 bl[184] br[184] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_185 bl[185] br[185] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_186 bl[186] br[186] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_187 bl[187] br[187] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_188 bl[188] br[188] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_189 bl[189] br[189] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_190 bl[190] br[190] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_191 bl[191] br[191] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_192 bl[192] br[192] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_193 bl[193] br[193] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_194 bl[194] br[194] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_195 bl[195] br[195] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_196 bl[196] br[196] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_197 bl[197] br[197] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_198 bl[198] br[198] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_199 bl[199] br[199] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_200 bl[200] br[200] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_201 bl[201] br[201] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_202 bl[202] br[202] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_203 bl[203] br[203] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_204 bl[204] br[204] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_205 bl[205] br[205] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_206 bl[206] br[206] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_207 bl[207] br[207] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_208 bl[208] br[208] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_209 bl[209] br[209] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_210 bl[210] br[210] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_211 bl[211] br[211] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_212 bl[212] br[212] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_213 bl[213] br[213] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_214 bl[214] br[214] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_215 bl[215] br[215] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_216 bl[216] br[216] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_217 bl[217] br[217] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_218 bl[218] br[218] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_219 bl[219] br[219] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_220 bl[220] br[220] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_221 bl[221] br[221] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_222 bl[222] br[222] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_223 bl[223] br[223] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_224 bl[224] br[224] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_225 bl[225] br[225] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_226 bl[226] br[226] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_227 bl[227] br[227] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_228 bl[228] br[228] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_229 bl[229] br[229] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_230 bl[230] br[230] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_231 bl[231] br[231] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_232 bl[232] br[232] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_233 bl[233] br[233] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_234 bl[234] br[234] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_235 bl[235] br[235] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_236 bl[236] br[236] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_237 bl[237] br[237] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_238 bl[238] br[238] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_239 bl[239] br[239] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_240 bl[240] br[240] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_241 bl[241] br[241] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_242 bl[242] br[242] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_243 bl[243] br[243] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_244 bl[244] br[244] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_245 bl[245] br[245] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_246 bl[246] br[246] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_247 bl[247] br[247] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_248 bl[248] br[248] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_249 bl[249] br[249] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_250 bl[250] br[250] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_251 bl[251] br[251] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_252 bl[252] br[252] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_253 bl[253] br[253] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_254 bl[254] br[254] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_255 bl[255] br[255] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_16_0 bl[0] br[0] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_1 bl[1] br[1] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_2 bl[2] br[2] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_3 bl[3] br[3] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_4 bl[4] br[4] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_5 bl[5] br[5] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_6 bl[6] br[6] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_7 bl[7] br[7] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_8 bl[8] br[8] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_9 bl[9] br[9] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_10 bl[10] br[10] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_11 bl[11] br[11] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_12 bl[12] br[12] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_13 bl[13] br[13] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_14 bl[14] br[14] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_15 bl[15] br[15] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_16 bl[16] br[16] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_17 bl[17] br[17] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_18 bl[18] br[18] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_19 bl[19] br[19] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_20 bl[20] br[20] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_21 bl[21] br[21] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_22 bl[22] br[22] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_23 bl[23] br[23] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_24 bl[24] br[24] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_25 bl[25] br[25] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_26 bl[26] br[26] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_27 bl[27] br[27] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_28 bl[28] br[28] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_29 bl[29] br[29] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_30 bl[30] br[30] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_31 bl[31] br[31] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_32 bl[32] br[32] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_33 bl[33] br[33] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_34 bl[34] br[34] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_35 bl[35] br[35] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_36 bl[36] br[36] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_37 bl[37] br[37] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_38 bl[38] br[38] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_39 bl[39] br[39] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_40 bl[40] br[40] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_41 bl[41] br[41] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_42 bl[42] br[42] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_43 bl[43] br[43] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_44 bl[44] br[44] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_45 bl[45] br[45] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_46 bl[46] br[46] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_47 bl[47] br[47] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_48 bl[48] br[48] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_49 bl[49] br[49] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_50 bl[50] br[50] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_51 bl[51] br[51] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_52 bl[52] br[52] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_53 bl[53] br[53] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_54 bl[54] br[54] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_55 bl[55] br[55] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_56 bl[56] br[56] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_57 bl[57] br[57] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_58 bl[58] br[58] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_59 bl[59] br[59] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_60 bl[60] br[60] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_61 bl[61] br[61] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_62 bl[62] br[62] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_63 bl[63] br[63] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_64 bl[64] br[64] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_65 bl[65] br[65] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_66 bl[66] br[66] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_67 bl[67] br[67] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_68 bl[68] br[68] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_69 bl[69] br[69] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_70 bl[70] br[70] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_71 bl[71] br[71] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_72 bl[72] br[72] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_73 bl[73] br[73] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_74 bl[74] br[74] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_75 bl[75] br[75] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_76 bl[76] br[76] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_77 bl[77] br[77] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_78 bl[78] br[78] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_79 bl[79] br[79] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_80 bl[80] br[80] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_81 bl[81] br[81] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_82 bl[82] br[82] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_83 bl[83] br[83] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_84 bl[84] br[84] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_85 bl[85] br[85] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_86 bl[86] br[86] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_87 bl[87] br[87] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_88 bl[88] br[88] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_89 bl[89] br[89] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_90 bl[90] br[90] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_91 bl[91] br[91] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_92 bl[92] br[92] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_93 bl[93] br[93] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_94 bl[94] br[94] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_95 bl[95] br[95] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_96 bl[96] br[96] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_97 bl[97] br[97] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_98 bl[98] br[98] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_99 bl[99] br[99] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_100 bl[100] br[100] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_101 bl[101] br[101] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_102 bl[102] br[102] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_103 bl[103] br[103] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_104 bl[104] br[104] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_105 bl[105] br[105] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_106 bl[106] br[106] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_107 bl[107] br[107] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_108 bl[108] br[108] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_109 bl[109] br[109] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_110 bl[110] br[110] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_111 bl[111] br[111] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_112 bl[112] br[112] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_113 bl[113] br[113] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_114 bl[114] br[114] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_115 bl[115] br[115] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_116 bl[116] br[116] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_117 bl[117] br[117] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_118 bl[118] br[118] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_119 bl[119] br[119] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_120 bl[120] br[120] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_121 bl[121] br[121] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_122 bl[122] br[122] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_123 bl[123] br[123] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_124 bl[124] br[124] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_125 bl[125] br[125] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_126 bl[126] br[126] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_127 bl[127] br[127] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_128 bl[128] br[128] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_129 bl[129] br[129] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_130 bl[130] br[130] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_131 bl[131] br[131] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_132 bl[132] br[132] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_133 bl[133] br[133] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_134 bl[134] br[134] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_135 bl[135] br[135] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_136 bl[136] br[136] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_137 bl[137] br[137] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_138 bl[138] br[138] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_139 bl[139] br[139] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_140 bl[140] br[140] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_141 bl[141] br[141] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_142 bl[142] br[142] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_143 bl[143] br[143] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_144 bl[144] br[144] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_145 bl[145] br[145] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_146 bl[146] br[146] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_147 bl[147] br[147] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_148 bl[148] br[148] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_149 bl[149] br[149] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_150 bl[150] br[150] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_151 bl[151] br[151] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_152 bl[152] br[152] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_153 bl[153] br[153] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_154 bl[154] br[154] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_155 bl[155] br[155] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_156 bl[156] br[156] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_157 bl[157] br[157] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_158 bl[158] br[158] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_159 bl[159] br[159] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_160 bl[160] br[160] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_161 bl[161] br[161] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_162 bl[162] br[162] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_163 bl[163] br[163] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_164 bl[164] br[164] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_165 bl[165] br[165] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_166 bl[166] br[166] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_167 bl[167] br[167] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_168 bl[168] br[168] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_169 bl[169] br[169] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_170 bl[170] br[170] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_171 bl[171] br[171] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_172 bl[172] br[172] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_173 bl[173] br[173] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_174 bl[174] br[174] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_175 bl[175] br[175] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_176 bl[176] br[176] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_177 bl[177] br[177] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_178 bl[178] br[178] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_179 bl[179] br[179] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_180 bl[180] br[180] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_181 bl[181] br[181] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_182 bl[182] br[182] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_183 bl[183] br[183] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_184 bl[184] br[184] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_185 bl[185] br[185] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_186 bl[186] br[186] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_187 bl[187] br[187] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_188 bl[188] br[188] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_189 bl[189] br[189] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_190 bl[190] br[190] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_191 bl[191] br[191] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_192 bl[192] br[192] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_193 bl[193] br[193] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_194 bl[194] br[194] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_195 bl[195] br[195] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_196 bl[196] br[196] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_197 bl[197] br[197] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_198 bl[198] br[198] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_199 bl[199] br[199] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_200 bl[200] br[200] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_201 bl[201] br[201] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_202 bl[202] br[202] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_203 bl[203] br[203] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_204 bl[204] br[204] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_205 bl[205] br[205] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_206 bl[206] br[206] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_207 bl[207] br[207] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_208 bl[208] br[208] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_209 bl[209] br[209] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_210 bl[210] br[210] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_211 bl[211] br[211] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_212 bl[212] br[212] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_213 bl[213] br[213] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_214 bl[214] br[214] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_215 bl[215] br[215] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_216 bl[216] br[216] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_217 bl[217] br[217] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_218 bl[218] br[218] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_219 bl[219] br[219] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_220 bl[220] br[220] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_221 bl[221] br[221] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_222 bl[222] br[222] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_223 bl[223] br[223] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_224 bl[224] br[224] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_225 bl[225] br[225] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_226 bl[226] br[226] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_227 bl[227] br[227] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_228 bl[228] br[228] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_229 bl[229] br[229] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_230 bl[230] br[230] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_231 bl[231] br[231] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_232 bl[232] br[232] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_233 bl[233] br[233] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_234 bl[234] br[234] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_235 bl[235] br[235] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_236 bl[236] br[236] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_237 bl[237] br[237] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_238 bl[238] br[238] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_239 bl[239] br[239] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_240 bl[240] br[240] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_241 bl[241] br[241] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_242 bl[242] br[242] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_243 bl[243] br[243] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_244 bl[244] br[244] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_245 bl[245] br[245] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_246 bl[246] br[246] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_247 bl[247] br[247] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_248 bl[248] br[248] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_249 bl[249] br[249] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_250 bl[250] br[250] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_251 bl[251] br[251] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_252 bl[252] br[252] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_253 bl[253] br[253] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_254 bl[254] br[254] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_255 bl[255] br[255] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_17_0 bl[0] br[0] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_1 bl[1] br[1] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_2 bl[2] br[2] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_3 bl[3] br[3] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_4 bl[4] br[4] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_5 bl[5] br[5] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_6 bl[6] br[6] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_7 bl[7] br[7] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_8 bl[8] br[8] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_9 bl[9] br[9] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_10 bl[10] br[10] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_11 bl[11] br[11] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_12 bl[12] br[12] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_13 bl[13] br[13] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_14 bl[14] br[14] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_15 bl[15] br[15] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_16 bl[16] br[16] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_17 bl[17] br[17] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_18 bl[18] br[18] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_19 bl[19] br[19] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_20 bl[20] br[20] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_21 bl[21] br[21] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_22 bl[22] br[22] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_23 bl[23] br[23] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_24 bl[24] br[24] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_25 bl[25] br[25] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_26 bl[26] br[26] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_27 bl[27] br[27] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_28 bl[28] br[28] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_29 bl[29] br[29] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_30 bl[30] br[30] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_31 bl[31] br[31] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_32 bl[32] br[32] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_33 bl[33] br[33] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_34 bl[34] br[34] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_35 bl[35] br[35] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_36 bl[36] br[36] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_37 bl[37] br[37] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_38 bl[38] br[38] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_39 bl[39] br[39] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_40 bl[40] br[40] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_41 bl[41] br[41] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_42 bl[42] br[42] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_43 bl[43] br[43] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_44 bl[44] br[44] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_45 bl[45] br[45] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_46 bl[46] br[46] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_47 bl[47] br[47] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_48 bl[48] br[48] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_49 bl[49] br[49] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_50 bl[50] br[50] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_51 bl[51] br[51] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_52 bl[52] br[52] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_53 bl[53] br[53] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_54 bl[54] br[54] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_55 bl[55] br[55] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_56 bl[56] br[56] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_57 bl[57] br[57] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_58 bl[58] br[58] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_59 bl[59] br[59] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_60 bl[60] br[60] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_61 bl[61] br[61] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_62 bl[62] br[62] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_63 bl[63] br[63] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_64 bl[64] br[64] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_65 bl[65] br[65] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_66 bl[66] br[66] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_67 bl[67] br[67] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_68 bl[68] br[68] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_69 bl[69] br[69] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_70 bl[70] br[70] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_71 bl[71] br[71] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_72 bl[72] br[72] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_73 bl[73] br[73] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_74 bl[74] br[74] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_75 bl[75] br[75] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_76 bl[76] br[76] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_77 bl[77] br[77] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_78 bl[78] br[78] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_79 bl[79] br[79] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_80 bl[80] br[80] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_81 bl[81] br[81] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_82 bl[82] br[82] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_83 bl[83] br[83] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_84 bl[84] br[84] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_85 bl[85] br[85] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_86 bl[86] br[86] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_87 bl[87] br[87] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_88 bl[88] br[88] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_89 bl[89] br[89] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_90 bl[90] br[90] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_91 bl[91] br[91] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_92 bl[92] br[92] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_93 bl[93] br[93] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_94 bl[94] br[94] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_95 bl[95] br[95] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_96 bl[96] br[96] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_97 bl[97] br[97] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_98 bl[98] br[98] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_99 bl[99] br[99] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_100 bl[100] br[100] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_101 bl[101] br[101] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_102 bl[102] br[102] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_103 bl[103] br[103] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_104 bl[104] br[104] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_105 bl[105] br[105] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_106 bl[106] br[106] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_107 bl[107] br[107] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_108 bl[108] br[108] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_109 bl[109] br[109] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_110 bl[110] br[110] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_111 bl[111] br[111] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_112 bl[112] br[112] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_113 bl[113] br[113] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_114 bl[114] br[114] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_115 bl[115] br[115] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_116 bl[116] br[116] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_117 bl[117] br[117] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_118 bl[118] br[118] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_119 bl[119] br[119] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_120 bl[120] br[120] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_121 bl[121] br[121] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_122 bl[122] br[122] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_123 bl[123] br[123] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_124 bl[124] br[124] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_125 bl[125] br[125] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_126 bl[126] br[126] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_127 bl[127] br[127] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_128 bl[128] br[128] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_129 bl[129] br[129] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_130 bl[130] br[130] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_131 bl[131] br[131] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_132 bl[132] br[132] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_133 bl[133] br[133] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_134 bl[134] br[134] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_135 bl[135] br[135] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_136 bl[136] br[136] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_137 bl[137] br[137] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_138 bl[138] br[138] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_139 bl[139] br[139] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_140 bl[140] br[140] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_141 bl[141] br[141] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_142 bl[142] br[142] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_143 bl[143] br[143] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_144 bl[144] br[144] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_145 bl[145] br[145] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_146 bl[146] br[146] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_147 bl[147] br[147] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_148 bl[148] br[148] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_149 bl[149] br[149] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_150 bl[150] br[150] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_151 bl[151] br[151] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_152 bl[152] br[152] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_153 bl[153] br[153] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_154 bl[154] br[154] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_155 bl[155] br[155] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_156 bl[156] br[156] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_157 bl[157] br[157] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_158 bl[158] br[158] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_159 bl[159] br[159] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_160 bl[160] br[160] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_161 bl[161] br[161] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_162 bl[162] br[162] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_163 bl[163] br[163] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_164 bl[164] br[164] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_165 bl[165] br[165] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_166 bl[166] br[166] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_167 bl[167] br[167] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_168 bl[168] br[168] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_169 bl[169] br[169] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_170 bl[170] br[170] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_171 bl[171] br[171] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_172 bl[172] br[172] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_173 bl[173] br[173] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_174 bl[174] br[174] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_175 bl[175] br[175] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_176 bl[176] br[176] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_177 bl[177] br[177] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_178 bl[178] br[178] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_179 bl[179] br[179] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_180 bl[180] br[180] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_181 bl[181] br[181] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_182 bl[182] br[182] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_183 bl[183] br[183] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_184 bl[184] br[184] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_185 bl[185] br[185] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_186 bl[186] br[186] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_187 bl[187] br[187] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_188 bl[188] br[188] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_189 bl[189] br[189] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_190 bl[190] br[190] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_191 bl[191] br[191] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_192 bl[192] br[192] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_193 bl[193] br[193] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_194 bl[194] br[194] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_195 bl[195] br[195] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_196 bl[196] br[196] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_197 bl[197] br[197] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_198 bl[198] br[198] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_199 bl[199] br[199] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_200 bl[200] br[200] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_201 bl[201] br[201] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_202 bl[202] br[202] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_203 bl[203] br[203] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_204 bl[204] br[204] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_205 bl[205] br[205] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_206 bl[206] br[206] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_207 bl[207] br[207] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_208 bl[208] br[208] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_209 bl[209] br[209] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_210 bl[210] br[210] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_211 bl[211] br[211] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_212 bl[212] br[212] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_213 bl[213] br[213] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_214 bl[214] br[214] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_215 bl[215] br[215] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_216 bl[216] br[216] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_217 bl[217] br[217] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_218 bl[218] br[218] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_219 bl[219] br[219] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_220 bl[220] br[220] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_221 bl[221] br[221] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_222 bl[222] br[222] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_223 bl[223] br[223] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_224 bl[224] br[224] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_225 bl[225] br[225] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_226 bl[226] br[226] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_227 bl[227] br[227] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_228 bl[228] br[228] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_229 bl[229] br[229] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_230 bl[230] br[230] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_231 bl[231] br[231] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_232 bl[232] br[232] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_233 bl[233] br[233] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_234 bl[234] br[234] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_235 bl[235] br[235] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_236 bl[236] br[236] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_237 bl[237] br[237] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_238 bl[238] br[238] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_239 bl[239] br[239] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_240 bl[240] br[240] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_241 bl[241] br[241] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_242 bl[242] br[242] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_243 bl[243] br[243] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_244 bl[244] br[244] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_245 bl[245] br[245] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_246 bl[246] br[246] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_247 bl[247] br[247] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_248 bl[248] br[248] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_249 bl[249] br[249] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_250 bl[250] br[250] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_251 bl[251] br[251] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_252 bl[252] br[252] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_253 bl[253] br[253] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_254 bl[254] br[254] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_255 bl[255] br[255] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_18_0 bl[0] br[0] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_1 bl[1] br[1] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_2 bl[2] br[2] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_3 bl[3] br[3] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_4 bl[4] br[4] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_5 bl[5] br[5] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_6 bl[6] br[6] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_7 bl[7] br[7] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_8 bl[8] br[8] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_9 bl[9] br[9] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_10 bl[10] br[10] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_11 bl[11] br[11] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_12 bl[12] br[12] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_13 bl[13] br[13] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_14 bl[14] br[14] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_15 bl[15] br[15] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_16 bl[16] br[16] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_17 bl[17] br[17] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_18 bl[18] br[18] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_19 bl[19] br[19] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_20 bl[20] br[20] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_21 bl[21] br[21] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_22 bl[22] br[22] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_23 bl[23] br[23] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_24 bl[24] br[24] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_25 bl[25] br[25] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_26 bl[26] br[26] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_27 bl[27] br[27] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_28 bl[28] br[28] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_29 bl[29] br[29] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_30 bl[30] br[30] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_31 bl[31] br[31] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_32 bl[32] br[32] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_33 bl[33] br[33] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_34 bl[34] br[34] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_35 bl[35] br[35] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_36 bl[36] br[36] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_37 bl[37] br[37] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_38 bl[38] br[38] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_39 bl[39] br[39] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_40 bl[40] br[40] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_41 bl[41] br[41] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_42 bl[42] br[42] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_43 bl[43] br[43] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_44 bl[44] br[44] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_45 bl[45] br[45] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_46 bl[46] br[46] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_47 bl[47] br[47] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_48 bl[48] br[48] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_49 bl[49] br[49] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_50 bl[50] br[50] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_51 bl[51] br[51] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_52 bl[52] br[52] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_53 bl[53] br[53] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_54 bl[54] br[54] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_55 bl[55] br[55] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_56 bl[56] br[56] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_57 bl[57] br[57] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_58 bl[58] br[58] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_59 bl[59] br[59] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_60 bl[60] br[60] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_61 bl[61] br[61] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_62 bl[62] br[62] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_63 bl[63] br[63] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_64 bl[64] br[64] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_65 bl[65] br[65] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_66 bl[66] br[66] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_67 bl[67] br[67] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_68 bl[68] br[68] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_69 bl[69] br[69] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_70 bl[70] br[70] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_71 bl[71] br[71] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_72 bl[72] br[72] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_73 bl[73] br[73] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_74 bl[74] br[74] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_75 bl[75] br[75] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_76 bl[76] br[76] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_77 bl[77] br[77] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_78 bl[78] br[78] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_79 bl[79] br[79] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_80 bl[80] br[80] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_81 bl[81] br[81] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_82 bl[82] br[82] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_83 bl[83] br[83] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_84 bl[84] br[84] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_85 bl[85] br[85] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_86 bl[86] br[86] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_87 bl[87] br[87] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_88 bl[88] br[88] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_89 bl[89] br[89] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_90 bl[90] br[90] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_91 bl[91] br[91] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_92 bl[92] br[92] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_93 bl[93] br[93] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_94 bl[94] br[94] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_95 bl[95] br[95] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_96 bl[96] br[96] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_97 bl[97] br[97] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_98 bl[98] br[98] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_99 bl[99] br[99] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_100 bl[100] br[100] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_101 bl[101] br[101] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_102 bl[102] br[102] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_103 bl[103] br[103] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_104 bl[104] br[104] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_105 bl[105] br[105] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_106 bl[106] br[106] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_107 bl[107] br[107] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_108 bl[108] br[108] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_109 bl[109] br[109] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_110 bl[110] br[110] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_111 bl[111] br[111] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_112 bl[112] br[112] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_113 bl[113] br[113] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_114 bl[114] br[114] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_115 bl[115] br[115] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_116 bl[116] br[116] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_117 bl[117] br[117] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_118 bl[118] br[118] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_119 bl[119] br[119] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_120 bl[120] br[120] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_121 bl[121] br[121] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_122 bl[122] br[122] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_123 bl[123] br[123] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_124 bl[124] br[124] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_125 bl[125] br[125] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_126 bl[126] br[126] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_127 bl[127] br[127] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_128 bl[128] br[128] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_129 bl[129] br[129] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_130 bl[130] br[130] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_131 bl[131] br[131] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_132 bl[132] br[132] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_133 bl[133] br[133] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_134 bl[134] br[134] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_135 bl[135] br[135] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_136 bl[136] br[136] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_137 bl[137] br[137] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_138 bl[138] br[138] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_139 bl[139] br[139] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_140 bl[140] br[140] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_141 bl[141] br[141] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_142 bl[142] br[142] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_143 bl[143] br[143] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_144 bl[144] br[144] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_145 bl[145] br[145] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_146 bl[146] br[146] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_147 bl[147] br[147] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_148 bl[148] br[148] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_149 bl[149] br[149] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_150 bl[150] br[150] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_151 bl[151] br[151] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_152 bl[152] br[152] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_153 bl[153] br[153] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_154 bl[154] br[154] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_155 bl[155] br[155] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_156 bl[156] br[156] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_157 bl[157] br[157] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_158 bl[158] br[158] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_159 bl[159] br[159] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_160 bl[160] br[160] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_161 bl[161] br[161] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_162 bl[162] br[162] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_163 bl[163] br[163] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_164 bl[164] br[164] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_165 bl[165] br[165] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_166 bl[166] br[166] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_167 bl[167] br[167] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_168 bl[168] br[168] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_169 bl[169] br[169] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_170 bl[170] br[170] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_171 bl[171] br[171] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_172 bl[172] br[172] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_173 bl[173] br[173] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_174 bl[174] br[174] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_175 bl[175] br[175] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_176 bl[176] br[176] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_177 bl[177] br[177] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_178 bl[178] br[178] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_179 bl[179] br[179] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_180 bl[180] br[180] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_181 bl[181] br[181] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_182 bl[182] br[182] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_183 bl[183] br[183] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_184 bl[184] br[184] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_185 bl[185] br[185] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_186 bl[186] br[186] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_187 bl[187] br[187] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_188 bl[188] br[188] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_189 bl[189] br[189] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_190 bl[190] br[190] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_191 bl[191] br[191] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_192 bl[192] br[192] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_193 bl[193] br[193] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_194 bl[194] br[194] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_195 bl[195] br[195] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_196 bl[196] br[196] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_197 bl[197] br[197] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_198 bl[198] br[198] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_199 bl[199] br[199] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_200 bl[200] br[200] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_201 bl[201] br[201] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_202 bl[202] br[202] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_203 bl[203] br[203] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_204 bl[204] br[204] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_205 bl[205] br[205] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_206 bl[206] br[206] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_207 bl[207] br[207] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_208 bl[208] br[208] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_209 bl[209] br[209] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_210 bl[210] br[210] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_211 bl[211] br[211] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_212 bl[212] br[212] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_213 bl[213] br[213] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_214 bl[214] br[214] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_215 bl[215] br[215] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_216 bl[216] br[216] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_217 bl[217] br[217] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_218 bl[218] br[218] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_219 bl[219] br[219] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_220 bl[220] br[220] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_221 bl[221] br[221] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_222 bl[222] br[222] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_223 bl[223] br[223] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_224 bl[224] br[224] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_225 bl[225] br[225] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_226 bl[226] br[226] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_227 bl[227] br[227] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_228 bl[228] br[228] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_229 bl[229] br[229] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_230 bl[230] br[230] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_231 bl[231] br[231] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_232 bl[232] br[232] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_233 bl[233] br[233] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_234 bl[234] br[234] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_235 bl[235] br[235] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_236 bl[236] br[236] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_237 bl[237] br[237] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_238 bl[238] br[238] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_239 bl[239] br[239] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_240 bl[240] br[240] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_241 bl[241] br[241] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_242 bl[242] br[242] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_243 bl[243] br[243] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_244 bl[244] br[244] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_245 bl[245] br[245] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_246 bl[246] br[246] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_247 bl[247] br[247] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_248 bl[248] br[248] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_249 bl[249] br[249] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_250 bl[250] br[250] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_251 bl[251] br[251] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_252 bl[252] br[252] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_253 bl[253] br[253] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_254 bl[254] br[254] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_255 bl[255] br[255] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_19_0 bl[0] br[0] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_1 bl[1] br[1] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_2 bl[2] br[2] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_3 bl[3] br[3] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_4 bl[4] br[4] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_5 bl[5] br[5] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_6 bl[6] br[6] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_7 bl[7] br[7] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_8 bl[8] br[8] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_9 bl[9] br[9] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_10 bl[10] br[10] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_11 bl[11] br[11] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_12 bl[12] br[12] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_13 bl[13] br[13] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_14 bl[14] br[14] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_15 bl[15] br[15] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_16 bl[16] br[16] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_17 bl[17] br[17] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_18 bl[18] br[18] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_19 bl[19] br[19] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_20 bl[20] br[20] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_21 bl[21] br[21] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_22 bl[22] br[22] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_23 bl[23] br[23] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_24 bl[24] br[24] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_25 bl[25] br[25] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_26 bl[26] br[26] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_27 bl[27] br[27] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_28 bl[28] br[28] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_29 bl[29] br[29] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_30 bl[30] br[30] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_31 bl[31] br[31] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_32 bl[32] br[32] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_33 bl[33] br[33] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_34 bl[34] br[34] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_35 bl[35] br[35] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_36 bl[36] br[36] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_37 bl[37] br[37] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_38 bl[38] br[38] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_39 bl[39] br[39] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_40 bl[40] br[40] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_41 bl[41] br[41] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_42 bl[42] br[42] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_43 bl[43] br[43] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_44 bl[44] br[44] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_45 bl[45] br[45] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_46 bl[46] br[46] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_47 bl[47] br[47] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_48 bl[48] br[48] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_49 bl[49] br[49] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_50 bl[50] br[50] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_51 bl[51] br[51] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_52 bl[52] br[52] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_53 bl[53] br[53] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_54 bl[54] br[54] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_55 bl[55] br[55] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_56 bl[56] br[56] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_57 bl[57] br[57] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_58 bl[58] br[58] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_59 bl[59] br[59] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_60 bl[60] br[60] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_61 bl[61] br[61] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_62 bl[62] br[62] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_63 bl[63] br[63] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_64 bl[64] br[64] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_65 bl[65] br[65] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_66 bl[66] br[66] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_67 bl[67] br[67] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_68 bl[68] br[68] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_69 bl[69] br[69] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_70 bl[70] br[70] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_71 bl[71] br[71] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_72 bl[72] br[72] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_73 bl[73] br[73] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_74 bl[74] br[74] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_75 bl[75] br[75] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_76 bl[76] br[76] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_77 bl[77] br[77] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_78 bl[78] br[78] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_79 bl[79] br[79] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_80 bl[80] br[80] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_81 bl[81] br[81] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_82 bl[82] br[82] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_83 bl[83] br[83] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_84 bl[84] br[84] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_85 bl[85] br[85] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_86 bl[86] br[86] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_87 bl[87] br[87] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_88 bl[88] br[88] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_89 bl[89] br[89] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_90 bl[90] br[90] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_91 bl[91] br[91] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_92 bl[92] br[92] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_93 bl[93] br[93] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_94 bl[94] br[94] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_95 bl[95] br[95] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_96 bl[96] br[96] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_97 bl[97] br[97] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_98 bl[98] br[98] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_99 bl[99] br[99] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_100 bl[100] br[100] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_101 bl[101] br[101] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_102 bl[102] br[102] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_103 bl[103] br[103] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_104 bl[104] br[104] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_105 bl[105] br[105] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_106 bl[106] br[106] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_107 bl[107] br[107] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_108 bl[108] br[108] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_109 bl[109] br[109] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_110 bl[110] br[110] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_111 bl[111] br[111] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_112 bl[112] br[112] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_113 bl[113] br[113] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_114 bl[114] br[114] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_115 bl[115] br[115] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_116 bl[116] br[116] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_117 bl[117] br[117] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_118 bl[118] br[118] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_119 bl[119] br[119] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_120 bl[120] br[120] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_121 bl[121] br[121] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_122 bl[122] br[122] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_123 bl[123] br[123] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_124 bl[124] br[124] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_125 bl[125] br[125] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_126 bl[126] br[126] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_127 bl[127] br[127] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_128 bl[128] br[128] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_129 bl[129] br[129] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_130 bl[130] br[130] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_131 bl[131] br[131] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_132 bl[132] br[132] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_133 bl[133] br[133] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_134 bl[134] br[134] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_135 bl[135] br[135] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_136 bl[136] br[136] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_137 bl[137] br[137] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_138 bl[138] br[138] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_139 bl[139] br[139] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_140 bl[140] br[140] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_141 bl[141] br[141] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_142 bl[142] br[142] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_143 bl[143] br[143] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_144 bl[144] br[144] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_145 bl[145] br[145] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_146 bl[146] br[146] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_147 bl[147] br[147] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_148 bl[148] br[148] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_149 bl[149] br[149] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_150 bl[150] br[150] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_151 bl[151] br[151] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_152 bl[152] br[152] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_153 bl[153] br[153] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_154 bl[154] br[154] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_155 bl[155] br[155] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_156 bl[156] br[156] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_157 bl[157] br[157] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_158 bl[158] br[158] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_159 bl[159] br[159] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_160 bl[160] br[160] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_161 bl[161] br[161] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_162 bl[162] br[162] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_163 bl[163] br[163] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_164 bl[164] br[164] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_165 bl[165] br[165] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_166 bl[166] br[166] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_167 bl[167] br[167] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_168 bl[168] br[168] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_169 bl[169] br[169] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_170 bl[170] br[170] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_171 bl[171] br[171] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_172 bl[172] br[172] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_173 bl[173] br[173] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_174 bl[174] br[174] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_175 bl[175] br[175] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_176 bl[176] br[176] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_177 bl[177] br[177] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_178 bl[178] br[178] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_179 bl[179] br[179] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_180 bl[180] br[180] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_181 bl[181] br[181] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_182 bl[182] br[182] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_183 bl[183] br[183] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_184 bl[184] br[184] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_185 bl[185] br[185] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_186 bl[186] br[186] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_187 bl[187] br[187] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_188 bl[188] br[188] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_189 bl[189] br[189] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_190 bl[190] br[190] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_191 bl[191] br[191] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_192 bl[192] br[192] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_193 bl[193] br[193] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_194 bl[194] br[194] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_195 bl[195] br[195] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_196 bl[196] br[196] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_197 bl[197] br[197] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_198 bl[198] br[198] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_199 bl[199] br[199] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_200 bl[200] br[200] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_201 bl[201] br[201] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_202 bl[202] br[202] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_203 bl[203] br[203] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_204 bl[204] br[204] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_205 bl[205] br[205] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_206 bl[206] br[206] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_207 bl[207] br[207] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_208 bl[208] br[208] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_209 bl[209] br[209] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_210 bl[210] br[210] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_211 bl[211] br[211] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_212 bl[212] br[212] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_213 bl[213] br[213] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_214 bl[214] br[214] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_215 bl[215] br[215] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_216 bl[216] br[216] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_217 bl[217] br[217] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_218 bl[218] br[218] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_219 bl[219] br[219] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_220 bl[220] br[220] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_221 bl[221] br[221] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_222 bl[222] br[222] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_223 bl[223] br[223] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_224 bl[224] br[224] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_225 bl[225] br[225] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_226 bl[226] br[226] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_227 bl[227] br[227] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_228 bl[228] br[228] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_229 bl[229] br[229] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_230 bl[230] br[230] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_231 bl[231] br[231] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_232 bl[232] br[232] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_233 bl[233] br[233] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_234 bl[234] br[234] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_235 bl[235] br[235] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_236 bl[236] br[236] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_237 bl[237] br[237] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_238 bl[238] br[238] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_239 bl[239] br[239] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_240 bl[240] br[240] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_241 bl[241] br[241] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_242 bl[242] br[242] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_243 bl[243] br[243] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_244 bl[244] br[244] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_245 bl[245] br[245] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_246 bl[246] br[246] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_247 bl[247] br[247] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_248 bl[248] br[248] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_249 bl[249] br[249] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_250 bl[250] br[250] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_251 bl[251] br[251] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_252 bl[252] br[252] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_253 bl[253] br[253] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_254 bl[254] br[254] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_255 bl[255] br[255] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_20_0 bl[0] br[0] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_1 bl[1] br[1] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_2 bl[2] br[2] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_3 bl[3] br[3] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_4 bl[4] br[4] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_5 bl[5] br[5] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_6 bl[6] br[6] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_7 bl[7] br[7] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_8 bl[8] br[8] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_9 bl[9] br[9] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_10 bl[10] br[10] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_11 bl[11] br[11] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_12 bl[12] br[12] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_13 bl[13] br[13] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_14 bl[14] br[14] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_15 bl[15] br[15] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_16 bl[16] br[16] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_17 bl[17] br[17] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_18 bl[18] br[18] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_19 bl[19] br[19] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_20 bl[20] br[20] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_21 bl[21] br[21] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_22 bl[22] br[22] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_23 bl[23] br[23] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_24 bl[24] br[24] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_25 bl[25] br[25] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_26 bl[26] br[26] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_27 bl[27] br[27] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_28 bl[28] br[28] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_29 bl[29] br[29] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_30 bl[30] br[30] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_31 bl[31] br[31] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_32 bl[32] br[32] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_33 bl[33] br[33] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_34 bl[34] br[34] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_35 bl[35] br[35] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_36 bl[36] br[36] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_37 bl[37] br[37] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_38 bl[38] br[38] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_39 bl[39] br[39] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_40 bl[40] br[40] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_41 bl[41] br[41] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_42 bl[42] br[42] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_43 bl[43] br[43] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_44 bl[44] br[44] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_45 bl[45] br[45] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_46 bl[46] br[46] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_47 bl[47] br[47] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_48 bl[48] br[48] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_49 bl[49] br[49] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_50 bl[50] br[50] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_51 bl[51] br[51] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_52 bl[52] br[52] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_53 bl[53] br[53] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_54 bl[54] br[54] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_55 bl[55] br[55] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_56 bl[56] br[56] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_57 bl[57] br[57] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_58 bl[58] br[58] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_59 bl[59] br[59] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_60 bl[60] br[60] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_61 bl[61] br[61] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_62 bl[62] br[62] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_63 bl[63] br[63] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_64 bl[64] br[64] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_65 bl[65] br[65] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_66 bl[66] br[66] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_67 bl[67] br[67] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_68 bl[68] br[68] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_69 bl[69] br[69] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_70 bl[70] br[70] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_71 bl[71] br[71] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_72 bl[72] br[72] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_73 bl[73] br[73] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_74 bl[74] br[74] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_75 bl[75] br[75] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_76 bl[76] br[76] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_77 bl[77] br[77] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_78 bl[78] br[78] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_79 bl[79] br[79] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_80 bl[80] br[80] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_81 bl[81] br[81] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_82 bl[82] br[82] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_83 bl[83] br[83] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_84 bl[84] br[84] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_85 bl[85] br[85] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_86 bl[86] br[86] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_87 bl[87] br[87] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_88 bl[88] br[88] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_89 bl[89] br[89] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_90 bl[90] br[90] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_91 bl[91] br[91] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_92 bl[92] br[92] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_93 bl[93] br[93] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_94 bl[94] br[94] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_95 bl[95] br[95] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_96 bl[96] br[96] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_97 bl[97] br[97] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_98 bl[98] br[98] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_99 bl[99] br[99] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_100 bl[100] br[100] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_101 bl[101] br[101] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_102 bl[102] br[102] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_103 bl[103] br[103] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_104 bl[104] br[104] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_105 bl[105] br[105] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_106 bl[106] br[106] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_107 bl[107] br[107] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_108 bl[108] br[108] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_109 bl[109] br[109] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_110 bl[110] br[110] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_111 bl[111] br[111] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_112 bl[112] br[112] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_113 bl[113] br[113] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_114 bl[114] br[114] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_115 bl[115] br[115] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_116 bl[116] br[116] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_117 bl[117] br[117] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_118 bl[118] br[118] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_119 bl[119] br[119] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_120 bl[120] br[120] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_121 bl[121] br[121] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_122 bl[122] br[122] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_123 bl[123] br[123] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_124 bl[124] br[124] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_125 bl[125] br[125] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_126 bl[126] br[126] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_127 bl[127] br[127] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_128 bl[128] br[128] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_129 bl[129] br[129] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_130 bl[130] br[130] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_131 bl[131] br[131] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_132 bl[132] br[132] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_133 bl[133] br[133] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_134 bl[134] br[134] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_135 bl[135] br[135] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_136 bl[136] br[136] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_137 bl[137] br[137] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_138 bl[138] br[138] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_139 bl[139] br[139] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_140 bl[140] br[140] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_141 bl[141] br[141] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_142 bl[142] br[142] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_143 bl[143] br[143] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_144 bl[144] br[144] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_145 bl[145] br[145] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_146 bl[146] br[146] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_147 bl[147] br[147] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_148 bl[148] br[148] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_149 bl[149] br[149] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_150 bl[150] br[150] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_151 bl[151] br[151] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_152 bl[152] br[152] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_153 bl[153] br[153] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_154 bl[154] br[154] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_155 bl[155] br[155] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_156 bl[156] br[156] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_157 bl[157] br[157] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_158 bl[158] br[158] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_159 bl[159] br[159] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_160 bl[160] br[160] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_161 bl[161] br[161] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_162 bl[162] br[162] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_163 bl[163] br[163] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_164 bl[164] br[164] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_165 bl[165] br[165] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_166 bl[166] br[166] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_167 bl[167] br[167] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_168 bl[168] br[168] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_169 bl[169] br[169] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_170 bl[170] br[170] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_171 bl[171] br[171] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_172 bl[172] br[172] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_173 bl[173] br[173] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_174 bl[174] br[174] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_175 bl[175] br[175] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_176 bl[176] br[176] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_177 bl[177] br[177] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_178 bl[178] br[178] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_179 bl[179] br[179] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_180 bl[180] br[180] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_181 bl[181] br[181] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_182 bl[182] br[182] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_183 bl[183] br[183] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_184 bl[184] br[184] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_185 bl[185] br[185] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_186 bl[186] br[186] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_187 bl[187] br[187] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_188 bl[188] br[188] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_189 bl[189] br[189] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_190 bl[190] br[190] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_191 bl[191] br[191] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_192 bl[192] br[192] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_193 bl[193] br[193] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_194 bl[194] br[194] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_195 bl[195] br[195] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_196 bl[196] br[196] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_197 bl[197] br[197] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_198 bl[198] br[198] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_199 bl[199] br[199] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_200 bl[200] br[200] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_201 bl[201] br[201] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_202 bl[202] br[202] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_203 bl[203] br[203] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_204 bl[204] br[204] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_205 bl[205] br[205] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_206 bl[206] br[206] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_207 bl[207] br[207] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_208 bl[208] br[208] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_209 bl[209] br[209] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_210 bl[210] br[210] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_211 bl[211] br[211] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_212 bl[212] br[212] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_213 bl[213] br[213] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_214 bl[214] br[214] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_215 bl[215] br[215] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_216 bl[216] br[216] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_217 bl[217] br[217] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_218 bl[218] br[218] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_219 bl[219] br[219] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_220 bl[220] br[220] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_221 bl[221] br[221] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_222 bl[222] br[222] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_223 bl[223] br[223] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_224 bl[224] br[224] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_225 bl[225] br[225] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_226 bl[226] br[226] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_227 bl[227] br[227] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_228 bl[228] br[228] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_229 bl[229] br[229] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_230 bl[230] br[230] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_231 bl[231] br[231] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_232 bl[232] br[232] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_233 bl[233] br[233] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_234 bl[234] br[234] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_235 bl[235] br[235] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_236 bl[236] br[236] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_237 bl[237] br[237] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_238 bl[238] br[238] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_239 bl[239] br[239] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_240 bl[240] br[240] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_241 bl[241] br[241] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_242 bl[242] br[242] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_243 bl[243] br[243] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_244 bl[244] br[244] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_245 bl[245] br[245] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_246 bl[246] br[246] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_247 bl[247] br[247] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_248 bl[248] br[248] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_249 bl[249] br[249] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_250 bl[250] br[250] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_251 bl[251] br[251] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_252 bl[252] br[252] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_253 bl[253] br[253] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_254 bl[254] br[254] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_255 bl[255] br[255] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_21_0 bl[0] br[0] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_1 bl[1] br[1] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_2 bl[2] br[2] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_3 bl[3] br[3] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_4 bl[4] br[4] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_5 bl[5] br[5] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_6 bl[6] br[6] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_7 bl[7] br[7] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_8 bl[8] br[8] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_9 bl[9] br[9] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_10 bl[10] br[10] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_11 bl[11] br[11] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_12 bl[12] br[12] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_13 bl[13] br[13] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_14 bl[14] br[14] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_15 bl[15] br[15] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_16 bl[16] br[16] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_17 bl[17] br[17] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_18 bl[18] br[18] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_19 bl[19] br[19] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_20 bl[20] br[20] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_21 bl[21] br[21] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_22 bl[22] br[22] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_23 bl[23] br[23] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_24 bl[24] br[24] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_25 bl[25] br[25] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_26 bl[26] br[26] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_27 bl[27] br[27] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_28 bl[28] br[28] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_29 bl[29] br[29] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_30 bl[30] br[30] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_31 bl[31] br[31] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_32 bl[32] br[32] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_33 bl[33] br[33] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_34 bl[34] br[34] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_35 bl[35] br[35] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_36 bl[36] br[36] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_37 bl[37] br[37] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_38 bl[38] br[38] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_39 bl[39] br[39] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_40 bl[40] br[40] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_41 bl[41] br[41] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_42 bl[42] br[42] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_43 bl[43] br[43] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_44 bl[44] br[44] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_45 bl[45] br[45] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_46 bl[46] br[46] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_47 bl[47] br[47] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_48 bl[48] br[48] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_49 bl[49] br[49] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_50 bl[50] br[50] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_51 bl[51] br[51] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_52 bl[52] br[52] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_53 bl[53] br[53] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_54 bl[54] br[54] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_55 bl[55] br[55] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_56 bl[56] br[56] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_57 bl[57] br[57] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_58 bl[58] br[58] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_59 bl[59] br[59] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_60 bl[60] br[60] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_61 bl[61] br[61] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_62 bl[62] br[62] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_63 bl[63] br[63] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_64 bl[64] br[64] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_65 bl[65] br[65] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_66 bl[66] br[66] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_67 bl[67] br[67] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_68 bl[68] br[68] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_69 bl[69] br[69] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_70 bl[70] br[70] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_71 bl[71] br[71] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_72 bl[72] br[72] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_73 bl[73] br[73] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_74 bl[74] br[74] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_75 bl[75] br[75] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_76 bl[76] br[76] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_77 bl[77] br[77] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_78 bl[78] br[78] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_79 bl[79] br[79] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_80 bl[80] br[80] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_81 bl[81] br[81] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_82 bl[82] br[82] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_83 bl[83] br[83] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_84 bl[84] br[84] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_85 bl[85] br[85] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_86 bl[86] br[86] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_87 bl[87] br[87] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_88 bl[88] br[88] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_89 bl[89] br[89] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_90 bl[90] br[90] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_91 bl[91] br[91] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_92 bl[92] br[92] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_93 bl[93] br[93] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_94 bl[94] br[94] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_95 bl[95] br[95] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_96 bl[96] br[96] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_97 bl[97] br[97] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_98 bl[98] br[98] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_99 bl[99] br[99] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_100 bl[100] br[100] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_101 bl[101] br[101] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_102 bl[102] br[102] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_103 bl[103] br[103] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_104 bl[104] br[104] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_105 bl[105] br[105] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_106 bl[106] br[106] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_107 bl[107] br[107] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_108 bl[108] br[108] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_109 bl[109] br[109] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_110 bl[110] br[110] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_111 bl[111] br[111] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_112 bl[112] br[112] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_113 bl[113] br[113] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_114 bl[114] br[114] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_115 bl[115] br[115] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_116 bl[116] br[116] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_117 bl[117] br[117] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_118 bl[118] br[118] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_119 bl[119] br[119] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_120 bl[120] br[120] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_121 bl[121] br[121] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_122 bl[122] br[122] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_123 bl[123] br[123] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_124 bl[124] br[124] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_125 bl[125] br[125] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_126 bl[126] br[126] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_127 bl[127] br[127] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_128 bl[128] br[128] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_129 bl[129] br[129] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_130 bl[130] br[130] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_131 bl[131] br[131] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_132 bl[132] br[132] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_133 bl[133] br[133] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_134 bl[134] br[134] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_135 bl[135] br[135] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_136 bl[136] br[136] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_137 bl[137] br[137] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_138 bl[138] br[138] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_139 bl[139] br[139] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_140 bl[140] br[140] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_141 bl[141] br[141] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_142 bl[142] br[142] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_143 bl[143] br[143] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_144 bl[144] br[144] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_145 bl[145] br[145] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_146 bl[146] br[146] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_147 bl[147] br[147] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_148 bl[148] br[148] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_149 bl[149] br[149] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_150 bl[150] br[150] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_151 bl[151] br[151] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_152 bl[152] br[152] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_153 bl[153] br[153] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_154 bl[154] br[154] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_155 bl[155] br[155] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_156 bl[156] br[156] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_157 bl[157] br[157] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_158 bl[158] br[158] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_159 bl[159] br[159] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_160 bl[160] br[160] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_161 bl[161] br[161] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_162 bl[162] br[162] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_163 bl[163] br[163] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_164 bl[164] br[164] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_165 bl[165] br[165] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_166 bl[166] br[166] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_167 bl[167] br[167] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_168 bl[168] br[168] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_169 bl[169] br[169] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_170 bl[170] br[170] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_171 bl[171] br[171] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_172 bl[172] br[172] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_173 bl[173] br[173] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_174 bl[174] br[174] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_175 bl[175] br[175] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_176 bl[176] br[176] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_177 bl[177] br[177] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_178 bl[178] br[178] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_179 bl[179] br[179] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_180 bl[180] br[180] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_181 bl[181] br[181] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_182 bl[182] br[182] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_183 bl[183] br[183] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_184 bl[184] br[184] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_185 bl[185] br[185] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_186 bl[186] br[186] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_187 bl[187] br[187] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_188 bl[188] br[188] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_189 bl[189] br[189] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_190 bl[190] br[190] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_191 bl[191] br[191] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_192 bl[192] br[192] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_193 bl[193] br[193] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_194 bl[194] br[194] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_195 bl[195] br[195] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_196 bl[196] br[196] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_197 bl[197] br[197] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_198 bl[198] br[198] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_199 bl[199] br[199] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_200 bl[200] br[200] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_201 bl[201] br[201] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_202 bl[202] br[202] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_203 bl[203] br[203] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_204 bl[204] br[204] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_205 bl[205] br[205] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_206 bl[206] br[206] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_207 bl[207] br[207] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_208 bl[208] br[208] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_209 bl[209] br[209] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_210 bl[210] br[210] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_211 bl[211] br[211] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_212 bl[212] br[212] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_213 bl[213] br[213] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_214 bl[214] br[214] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_215 bl[215] br[215] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_216 bl[216] br[216] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_217 bl[217] br[217] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_218 bl[218] br[218] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_219 bl[219] br[219] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_220 bl[220] br[220] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_221 bl[221] br[221] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_222 bl[222] br[222] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_223 bl[223] br[223] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_224 bl[224] br[224] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_225 bl[225] br[225] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_226 bl[226] br[226] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_227 bl[227] br[227] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_228 bl[228] br[228] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_229 bl[229] br[229] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_230 bl[230] br[230] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_231 bl[231] br[231] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_232 bl[232] br[232] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_233 bl[233] br[233] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_234 bl[234] br[234] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_235 bl[235] br[235] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_236 bl[236] br[236] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_237 bl[237] br[237] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_238 bl[238] br[238] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_239 bl[239] br[239] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_240 bl[240] br[240] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_241 bl[241] br[241] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_242 bl[242] br[242] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_243 bl[243] br[243] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_244 bl[244] br[244] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_245 bl[245] br[245] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_246 bl[246] br[246] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_247 bl[247] br[247] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_248 bl[248] br[248] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_249 bl[249] br[249] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_250 bl[250] br[250] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_251 bl[251] br[251] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_252 bl[252] br[252] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_253 bl[253] br[253] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_254 bl[254] br[254] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_255 bl[255] br[255] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_22_0 bl[0] br[0] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_1 bl[1] br[1] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_2 bl[2] br[2] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_3 bl[3] br[3] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_4 bl[4] br[4] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_5 bl[5] br[5] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_6 bl[6] br[6] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_7 bl[7] br[7] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_8 bl[8] br[8] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_9 bl[9] br[9] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_10 bl[10] br[10] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_11 bl[11] br[11] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_12 bl[12] br[12] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_13 bl[13] br[13] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_14 bl[14] br[14] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_15 bl[15] br[15] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_16 bl[16] br[16] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_17 bl[17] br[17] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_18 bl[18] br[18] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_19 bl[19] br[19] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_20 bl[20] br[20] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_21 bl[21] br[21] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_22 bl[22] br[22] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_23 bl[23] br[23] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_24 bl[24] br[24] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_25 bl[25] br[25] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_26 bl[26] br[26] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_27 bl[27] br[27] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_28 bl[28] br[28] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_29 bl[29] br[29] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_30 bl[30] br[30] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_31 bl[31] br[31] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_32 bl[32] br[32] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_33 bl[33] br[33] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_34 bl[34] br[34] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_35 bl[35] br[35] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_36 bl[36] br[36] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_37 bl[37] br[37] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_38 bl[38] br[38] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_39 bl[39] br[39] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_40 bl[40] br[40] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_41 bl[41] br[41] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_42 bl[42] br[42] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_43 bl[43] br[43] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_44 bl[44] br[44] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_45 bl[45] br[45] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_46 bl[46] br[46] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_47 bl[47] br[47] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_48 bl[48] br[48] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_49 bl[49] br[49] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_50 bl[50] br[50] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_51 bl[51] br[51] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_52 bl[52] br[52] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_53 bl[53] br[53] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_54 bl[54] br[54] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_55 bl[55] br[55] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_56 bl[56] br[56] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_57 bl[57] br[57] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_58 bl[58] br[58] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_59 bl[59] br[59] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_60 bl[60] br[60] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_61 bl[61] br[61] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_62 bl[62] br[62] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_63 bl[63] br[63] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_64 bl[64] br[64] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_65 bl[65] br[65] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_66 bl[66] br[66] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_67 bl[67] br[67] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_68 bl[68] br[68] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_69 bl[69] br[69] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_70 bl[70] br[70] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_71 bl[71] br[71] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_72 bl[72] br[72] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_73 bl[73] br[73] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_74 bl[74] br[74] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_75 bl[75] br[75] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_76 bl[76] br[76] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_77 bl[77] br[77] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_78 bl[78] br[78] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_79 bl[79] br[79] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_80 bl[80] br[80] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_81 bl[81] br[81] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_82 bl[82] br[82] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_83 bl[83] br[83] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_84 bl[84] br[84] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_85 bl[85] br[85] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_86 bl[86] br[86] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_87 bl[87] br[87] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_88 bl[88] br[88] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_89 bl[89] br[89] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_90 bl[90] br[90] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_91 bl[91] br[91] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_92 bl[92] br[92] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_93 bl[93] br[93] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_94 bl[94] br[94] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_95 bl[95] br[95] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_96 bl[96] br[96] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_97 bl[97] br[97] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_98 bl[98] br[98] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_99 bl[99] br[99] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_100 bl[100] br[100] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_101 bl[101] br[101] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_102 bl[102] br[102] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_103 bl[103] br[103] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_104 bl[104] br[104] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_105 bl[105] br[105] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_106 bl[106] br[106] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_107 bl[107] br[107] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_108 bl[108] br[108] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_109 bl[109] br[109] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_110 bl[110] br[110] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_111 bl[111] br[111] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_112 bl[112] br[112] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_113 bl[113] br[113] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_114 bl[114] br[114] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_115 bl[115] br[115] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_116 bl[116] br[116] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_117 bl[117] br[117] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_118 bl[118] br[118] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_119 bl[119] br[119] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_120 bl[120] br[120] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_121 bl[121] br[121] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_122 bl[122] br[122] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_123 bl[123] br[123] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_124 bl[124] br[124] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_125 bl[125] br[125] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_126 bl[126] br[126] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_127 bl[127] br[127] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_128 bl[128] br[128] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_129 bl[129] br[129] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_130 bl[130] br[130] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_131 bl[131] br[131] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_132 bl[132] br[132] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_133 bl[133] br[133] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_134 bl[134] br[134] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_135 bl[135] br[135] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_136 bl[136] br[136] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_137 bl[137] br[137] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_138 bl[138] br[138] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_139 bl[139] br[139] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_140 bl[140] br[140] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_141 bl[141] br[141] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_142 bl[142] br[142] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_143 bl[143] br[143] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_144 bl[144] br[144] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_145 bl[145] br[145] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_146 bl[146] br[146] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_147 bl[147] br[147] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_148 bl[148] br[148] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_149 bl[149] br[149] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_150 bl[150] br[150] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_151 bl[151] br[151] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_152 bl[152] br[152] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_153 bl[153] br[153] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_154 bl[154] br[154] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_155 bl[155] br[155] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_156 bl[156] br[156] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_157 bl[157] br[157] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_158 bl[158] br[158] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_159 bl[159] br[159] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_160 bl[160] br[160] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_161 bl[161] br[161] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_162 bl[162] br[162] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_163 bl[163] br[163] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_164 bl[164] br[164] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_165 bl[165] br[165] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_166 bl[166] br[166] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_167 bl[167] br[167] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_168 bl[168] br[168] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_169 bl[169] br[169] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_170 bl[170] br[170] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_171 bl[171] br[171] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_172 bl[172] br[172] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_173 bl[173] br[173] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_174 bl[174] br[174] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_175 bl[175] br[175] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_176 bl[176] br[176] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_177 bl[177] br[177] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_178 bl[178] br[178] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_179 bl[179] br[179] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_180 bl[180] br[180] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_181 bl[181] br[181] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_182 bl[182] br[182] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_183 bl[183] br[183] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_184 bl[184] br[184] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_185 bl[185] br[185] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_186 bl[186] br[186] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_187 bl[187] br[187] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_188 bl[188] br[188] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_189 bl[189] br[189] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_190 bl[190] br[190] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_191 bl[191] br[191] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_192 bl[192] br[192] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_193 bl[193] br[193] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_194 bl[194] br[194] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_195 bl[195] br[195] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_196 bl[196] br[196] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_197 bl[197] br[197] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_198 bl[198] br[198] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_199 bl[199] br[199] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_200 bl[200] br[200] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_201 bl[201] br[201] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_202 bl[202] br[202] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_203 bl[203] br[203] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_204 bl[204] br[204] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_205 bl[205] br[205] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_206 bl[206] br[206] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_207 bl[207] br[207] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_208 bl[208] br[208] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_209 bl[209] br[209] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_210 bl[210] br[210] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_211 bl[211] br[211] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_212 bl[212] br[212] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_213 bl[213] br[213] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_214 bl[214] br[214] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_215 bl[215] br[215] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_216 bl[216] br[216] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_217 bl[217] br[217] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_218 bl[218] br[218] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_219 bl[219] br[219] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_220 bl[220] br[220] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_221 bl[221] br[221] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_222 bl[222] br[222] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_223 bl[223] br[223] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_224 bl[224] br[224] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_225 bl[225] br[225] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_226 bl[226] br[226] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_227 bl[227] br[227] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_228 bl[228] br[228] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_229 bl[229] br[229] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_230 bl[230] br[230] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_231 bl[231] br[231] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_232 bl[232] br[232] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_233 bl[233] br[233] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_234 bl[234] br[234] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_235 bl[235] br[235] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_236 bl[236] br[236] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_237 bl[237] br[237] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_238 bl[238] br[238] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_239 bl[239] br[239] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_240 bl[240] br[240] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_241 bl[241] br[241] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_242 bl[242] br[242] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_243 bl[243] br[243] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_244 bl[244] br[244] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_245 bl[245] br[245] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_246 bl[246] br[246] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_247 bl[247] br[247] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_248 bl[248] br[248] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_249 bl[249] br[249] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_250 bl[250] br[250] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_251 bl[251] br[251] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_252 bl[252] br[252] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_253 bl[253] br[253] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_254 bl[254] br[254] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_255 bl[255] br[255] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_23_0 bl[0] br[0] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_1 bl[1] br[1] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_2 bl[2] br[2] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_3 bl[3] br[3] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_4 bl[4] br[4] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_5 bl[5] br[5] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_6 bl[6] br[6] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_7 bl[7] br[7] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_8 bl[8] br[8] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_9 bl[9] br[9] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_10 bl[10] br[10] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_11 bl[11] br[11] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_12 bl[12] br[12] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_13 bl[13] br[13] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_14 bl[14] br[14] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_15 bl[15] br[15] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_16 bl[16] br[16] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_17 bl[17] br[17] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_18 bl[18] br[18] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_19 bl[19] br[19] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_20 bl[20] br[20] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_21 bl[21] br[21] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_22 bl[22] br[22] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_23 bl[23] br[23] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_24 bl[24] br[24] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_25 bl[25] br[25] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_26 bl[26] br[26] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_27 bl[27] br[27] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_28 bl[28] br[28] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_29 bl[29] br[29] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_30 bl[30] br[30] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_31 bl[31] br[31] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_32 bl[32] br[32] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_33 bl[33] br[33] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_34 bl[34] br[34] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_35 bl[35] br[35] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_36 bl[36] br[36] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_37 bl[37] br[37] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_38 bl[38] br[38] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_39 bl[39] br[39] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_40 bl[40] br[40] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_41 bl[41] br[41] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_42 bl[42] br[42] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_43 bl[43] br[43] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_44 bl[44] br[44] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_45 bl[45] br[45] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_46 bl[46] br[46] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_47 bl[47] br[47] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_48 bl[48] br[48] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_49 bl[49] br[49] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_50 bl[50] br[50] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_51 bl[51] br[51] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_52 bl[52] br[52] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_53 bl[53] br[53] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_54 bl[54] br[54] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_55 bl[55] br[55] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_56 bl[56] br[56] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_57 bl[57] br[57] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_58 bl[58] br[58] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_59 bl[59] br[59] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_60 bl[60] br[60] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_61 bl[61] br[61] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_62 bl[62] br[62] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_63 bl[63] br[63] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_64 bl[64] br[64] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_65 bl[65] br[65] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_66 bl[66] br[66] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_67 bl[67] br[67] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_68 bl[68] br[68] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_69 bl[69] br[69] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_70 bl[70] br[70] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_71 bl[71] br[71] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_72 bl[72] br[72] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_73 bl[73] br[73] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_74 bl[74] br[74] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_75 bl[75] br[75] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_76 bl[76] br[76] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_77 bl[77] br[77] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_78 bl[78] br[78] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_79 bl[79] br[79] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_80 bl[80] br[80] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_81 bl[81] br[81] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_82 bl[82] br[82] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_83 bl[83] br[83] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_84 bl[84] br[84] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_85 bl[85] br[85] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_86 bl[86] br[86] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_87 bl[87] br[87] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_88 bl[88] br[88] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_89 bl[89] br[89] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_90 bl[90] br[90] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_91 bl[91] br[91] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_92 bl[92] br[92] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_93 bl[93] br[93] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_94 bl[94] br[94] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_95 bl[95] br[95] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_96 bl[96] br[96] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_97 bl[97] br[97] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_98 bl[98] br[98] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_99 bl[99] br[99] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_100 bl[100] br[100] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_101 bl[101] br[101] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_102 bl[102] br[102] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_103 bl[103] br[103] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_104 bl[104] br[104] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_105 bl[105] br[105] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_106 bl[106] br[106] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_107 bl[107] br[107] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_108 bl[108] br[108] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_109 bl[109] br[109] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_110 bl[110] br[110] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_111 bl[111] br[111] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_112 bl[112] br[112] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_113 bl[113] br[113] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_114 bl[114] br[114] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_115 bl[115] br[115] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_116 bl[116] br[116] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_117 bl[117] br[117] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_118 bl[118] br[118] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_119 bl[119] br[119] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_120 bl[120] br[120] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_121 bl[121] br[121] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_122 bl[122] br[122] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_123 bl[123] br[123] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_124 bl[124] br[124] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_125 bl[125] br[125] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_126 bl[126] br[126] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_127 bl[127] br[127] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_128 bl[128] br[128] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_129 bl[129] br[129] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_130 bl[130] br[130] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_131 bl[131] br[131] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_132 bl[132] br[132] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_133 bl[133] br[133] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_134 bl[134] br[134] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_135 bl[135] br[135] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_136 bl[136] br[136] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_137 bl[137] br[137] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_138 bl[138] br[138] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_139 bl[139] br[139] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_140 bl[140] br[140] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_141 bl[141] br[141] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_142 bl[142] br[142] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_143 bl[143] br[143] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_144 bl[144] br[144] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_145 bl[145] br[145] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_146 bl[146] br[146] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_147 bl[147] br[147] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_148 bl[148] br[148] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_149 bl[149] br[149] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_150 bl[150] br[150] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_151 bl[151] br[151] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_152 bl[152] br[152] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_153 bl[153] br[153] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_154 bl[154] br[154] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_155 bl[155] br[155] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_156 bl[156] br[156] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_157 bl[157] br[157] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_158 bl[158] br[158] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_159 bl[159] br[159] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_160 bl[160] br[160] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_161 bl[161] br[161] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_162 bl[162] br[162] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_163 bl[163] br[163] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_164 bl[164] br[164] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_165 bl[165] br[165] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_166 bl[166] br[166] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_167 bl[167] br[167] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_168 bl[168] br[168] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_169 bl[169] br[169] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_170 bl[170] br[170] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_171 bl[171] br[171] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_172 bl[172] br[172] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_173 bl[173] br[173] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_174 bl[174] br[174] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_175 bl[175] br[175] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_176 bl[176] br[176] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_177 bl[177] br[177] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_178 bl[178] br[178] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_179 bl[179] br[179] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_180 bl[180] br[180] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_181 bl[181] br[181] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_182 bl[182] br[182] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_183 bl[183] br[183] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_184 bl[184] br[184] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_185 bl[185] br[185] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_186 bl[186] br[186] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_187 bl[187] br[187] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_188 bl[188] br[188] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_189 bl[189] br[189] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_190 bl[190] br[190] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_191 bl[191] br[191] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_192 bl[192] br[192] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_193 bl[193] br[193] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_194 bl[194] br[194] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_195 bl[195] br[195] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_196 bl[196] br[196] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_197 bl[197] br[197] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_198 bl[198] br[198] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_199 bl[199] br[199] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_200 bl[200] br[200] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_201 bl[201] br[201] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_202 bl[202] br[202] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_203 bl[203] br[203] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_204 bl[204] br[204] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_205 bl[205] br[205] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_206 bl[206] br[206] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_207 bl[207] br[207] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_208 bl[208] br[208] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_209 bl[209] br[209] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_210 bl[210] br[210] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_211 bl[211] br[211] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_212 bl[212] br[212] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_213 bl[213] br[213] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_214 bl[214] br[214] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_215 bl[215] br[215] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_216 bl[216] br[216] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_217 bl[217] br[217] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_218 bl[218] br[218] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_219 bl[219] br[219] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_220 bl[220] br[220] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_221 bl[221] br[221] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_222 bl[222] br[222] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_223 bl[223] br[223] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_224 bl[224] br[224] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_225 bl[225] br[225] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_226 bl[226] br[226] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_227 bl[227] br[227] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_228 bl[228] br[228] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_229 bl[229] br[229] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_230 bl[230] br[230] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_231 bl[231] br[231] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_232 bl[232] br[232] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_233 bl[233] br[233] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_234 bl[234] br[234] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_235 bl[235] br[235] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_236 bl[236] br[236] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_237 bl[237] br[237] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_238 bl[238] br[238] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_239 bl[239] br[239] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_240 bl[240] br[240] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_241 bl[241] br[241] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_242 bl[242] br[242] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_243 bl[243] br[243] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_244 bl[244] br[244] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_245 bl[245] br[245] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_246 bl[246] br[246] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_247 bl[247] br[247] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_248 bl[248] br[248] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_249 bl[249] br[249] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_250 bl[250] br[250] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_251 bl[251] br[251] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_252 bl[252] br[252] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_253 bl[253] br[253] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_254 bl[254] br[254] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_255 bl[255] br[255] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_24_0 bl[0] br[0] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_1 bl[1] br[1] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_2 bl[2] br[2] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_3 bl[3] br[3] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_4 bl[4] br[4] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_5 bl[5] br[5] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_6 bl[6] br[6] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_7 bl[7] br[7] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_8 bl[8] br[8] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_9 bl[9] br[9] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_10 bl[10] br[10] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_11 bl[11] br[11] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_12 bl[12] br[12] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_13 bl[13] br[13] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_14 bl[14] br[14] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_15 bl[15] br[15] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_16 bl[16] br[16] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_17 bl[17] br[17] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_18 bl[18] br[18] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_19 bl[19] br[19] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_20 bl[20] br[20] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_21 bl[21] br[21] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_22 bl[22] br[22] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_23 bl[23] br[23] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_24 bl[24] br[24] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_25 bl[25] br[25] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_26 bl[26] br[26] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_27 bl[27] br[27] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_28 bl[28] br[28] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_29 bl[29] br[29] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_30 bl[30] br[30] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_31 bl[31] br[31] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_32 bl[32] br[32] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_33 bl[33] br[33] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_34 bl[34] br[34] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_35 bl[35] br[35] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_36 bl[36] br[36] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_37 bl[37] br[37] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_38 bl[38] br[38] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_39 bl[39] br[39] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_40 bl[40] br[40] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_41 bl[41] br[41] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_42 bl[42] br[42] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_43 bl[43] br[43] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_44 bl[44] br[44] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_45 bl[45] br[45] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_46 bl[46] br[46] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_47 bl[47] br[47] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_48 bl[48] br[48] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_49 bl[49] br[49] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_50 bl[50] br[50] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_51 bl[51] br[51] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_52 bl[52] br[52] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_53 bl[53] br[53] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_54 bl[54] br[54] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_55 bl[55] br[55] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_56 bl[56] br[56] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_57 bl[57] br[57] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_58 bl[58] br[58] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_59 bl[59] br[59] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_60 bl[60] br[60] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_61 bl[61] br[61] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_62 bl[62] br[62] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_63 bl[63] br[63] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_64 bl[64] br[64] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_65 bl[65] br[65] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_66 bl[66] br[66] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_67 bl[67] br[67] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_68 bl[68] br[68] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_69 bl[69] br[69] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_70 bl[70] br[70] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_71 bl[71] br[71] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_72 bl[72] br[72] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_73 bl[73] br[73] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_74 bl[74] br[74] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_75 bl[75] br[75] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_76 bl[76] br[76] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_77 bl[77] br[77] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_78 bl[78] br[78] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_79 bl[79] br[79] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_80 bl[80] br[80] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_81 bl[81] br[81] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_82 bl[82] br[82] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_83 bl[83] br[83] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_84 bl[84] br[84] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_85 bl[85] br[85] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_86 bl[86] br[86] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_87 bl[87] br[87] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_88 bl[88] br[88] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_89 bl[89] br[89] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_90 bl[90] br[90] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_91 bl[91] br[91] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_92 bl[92] br[92] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_93 bl[93] br[93] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_94 bl[94] br[94] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_95 bl[95] br[95] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_96 bl[96] br[96] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_97 bl[97] br[97] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_98 bl[98] br[98] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_99 bl[99] br[99] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_100 bl[100] br[100] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_101 bl[101] br[101] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_102 bl[102] br[102] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_103 bl[103] br[103] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_104 bl[104] br[104] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_105 bl[105] br[105] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_106 bl[106] br[106] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_107 bl[107] br[107] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_108 bl[108] br[108] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_109 bl[109] br[109] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_110 bl[110] br[110] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_111 bl[111] br[111] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_112 bl[112] br[112] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_113 bl[113] br[113] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_114 bl[114] br[114] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_115 bl[115] br[115] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_116 bl[116] br[116] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_117 bl[117] br[117] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_118 bl[118] br[118] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_119 bl[119] br[119] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_120 bl[120] br[120] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_121 bl[121] br[121] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_122 bl[122] br[122] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_123 bl[123] br[123] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_124 bl[124] br[124] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_125 bl[125] br[125] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_126 bl[126] br[126] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_127 bl[127] br[127] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_128 bl[128] br[128] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_129 bl[129] br[129] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_130 bl[130] br[130] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_131 bl[131] br[131] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_132 bl[132] br[132] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_133 bl[133] br[133] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_134 bl[134] br[134] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_135 bl[135] br[135] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_136 bl[136] br[136] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_137 bl[137] br[137] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_138 bl[138] br[138] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_139 bl[139] br[139] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_140 bl[140] br[140] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_141 bl[141] br[141] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_142 bl[142] br[142] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_143 bl[143] br[143] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_144 bl[144] br[144] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_145 bl[145] br[145] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_146 bl[146] br[146] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_147 bl[147] br[147] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_148 bl[148] br[148] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_149 bl[149] br[149] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_150 bl[150] br[150] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_151 bl[151] br[151] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_152 bl[152] br[152] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_153 bl[153] br[153] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_154 bl[154] br[154] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_155 bl[155] br[155] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_156 bl[156] br[156] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_157 bl[157] br[157] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_158 bl[158] br[158] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_159 bl[159] br[159] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_160 bl[160] br[160] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_161 bl[161] br[161] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_162 bl[162] br[162] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_163 bl[163] br[163] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_164 bl[164] br[164] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_165 bl[165] br[165] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_166 bl[166] br[166] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_167 bl[167] br[167] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_168 bl[168] br[168] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_169 bl[169] br[169] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_170 bl[170] br[170] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_171 bl[171] br[171] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_172 bl[172] br[172] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_173 bl[173] br[173] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_174 bl[174] br[174] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_175 bl[175] br[175] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_176 bl[176] br[176] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_177 bl[177] br[177] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_178 bl[178] br[178] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_179 bl[179] br[179] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_180 bl[180] br[180] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_181 bl[181] br[181] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_182 bl[182] br[182] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_183 bl[183] br[183] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_184 bl[184] br[184] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_185 bl[185] br[185] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_186 bl[186] br[186] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_187 bl[187] br[187] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_188 bl[188] br[188] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_189 bl[189] br[189] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_190 bl[190] br[190] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_191 bl[191] br[191] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_192 bl[192] br[192] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_193 bl[193] br[193] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_194 bl[194] br[194] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_195 bl[195] br[195] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_196 bl[196] br[196] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_197 bl[197] br[197] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_198 bl[198] br[198] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_199 bl[199] br[199] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_200 bl[200] br[200] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_201 bl[201] br[201] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_202 bl[202] br[202] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_203 bl[203] br[203] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_204 bl[204] br[204] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_205 bl[205] br[205] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_206 bl[206] br[206] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_207 bl[207] br[207] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_208 bl[208] br[208] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_209 bl[209] br[209] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_210 bl[210] br[210] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_211 bl[211] br[211] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_212 bl[212] br[212] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_213 bl[213] br[213] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_214 bl[214] br[214] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_215 bl[215] br[215] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_216 bl[216] br[216] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_217 bl[217] br[217] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_218 bl[218] br[218] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_219 bl[219] br[219] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_220 bl[220] br[220] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_221 bl[221] br[221] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_222 bl[222] br[222] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_223 bl[223] br[223] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_224 bl[224] br[224] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_225 bl[225] br[225] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_226 bl[226] br[226] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_227 bl[227] br[227] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_228 bl[228] br[228] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_229 bl[229] br[229] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_230 bl[230] br[230] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_231 bl[231] br[231] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_232 bl[232] br[232] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_233 bl[233] br[233] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_234 bl[234] br[234] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_235 bl[235] br[235] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_236 bl[236] br[236] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_237 bl[237] br[237] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_238 bl[238] br[238] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_239 bl[239] br[239] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_240 bl[240] br[240] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_241 bl[241] br[241] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_242 bl[242] br[242] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_243 bl[243] br[243] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_244 bl[244] br[244] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_245 bl[245] br[245] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_246 bl[246] br[246] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_247 bl[247] br[247] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_248 bl[248] br[248] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_249 bl[249] br[249] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_250 bl[250] br[250] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_251 bl[251] br[251] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_252 bl[252] br[252] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_253 bl[253] br[253] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_254 bl[254] br[254] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_255 bl[255] br[255] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_25_0 bl[0] br[0] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_1 bl[1] br[1] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_2 bl[2] br[2] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_3 bl[3] br[3] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_4 bl[4] br[4] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_5 bl[5] br[5] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_6 bl[6] br[6] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_7 bl[7] br[7] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_8 bl[8] br[8] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_9 bl[9] br[9] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_10 bl[10] br[10] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_11 bl[11] br[11] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_12 bl[12] br[12] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_13 bl[13] br[13] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_14 bl[14] br[14] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_15 bl[15] br[15] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_16 bl[16] br[16] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_17 bl[17] br[17] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_18 bl[18] br[18] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_19 bl[19] br[19] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_20 bl[20] br[20] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_21 bl[21] br[21] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_22 bl[22] br[22] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_23 bl[23] br[23] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_24 bl[24] br[24] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_25 bl[25] br[25] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_26 bl[26] br[26] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_27 bl[27] br[27] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_28 bl[28] br[28] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_29 bl[29] br[29] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_30 bl[30] br[30] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_31 bl[31] br[31] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_32 bl[32] br[32] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_33 bl[33] br[33] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_34 bl[34] br[34] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_35 bl[35] br[35] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_36 bl[36] br[36] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_37 bl[37] br[37] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_38 bl[38] br[38] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_39 bl[39] br[39] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_40 bl[40] br[40] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_41 bl[41] br[41] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_42 bl[42] br[42] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_43 bl[43] br[43] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_44 bl[44] br[44] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_45 bl[45] br[45] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_46 bl[46] br[46] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_47 bl[47] br[47] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_48 bl[48] br[48] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_49 bl[49] br[49] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_50 bl[50] br[50] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_51 bl[51] br[51] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_52 bl[52] br[52] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_53 bl[53] br[53] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_54 bl[54] br[54] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_55 bl[55] br[55] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_56 bl[56] br[56] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_57 bl[57] br[57] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_58 bl[58] br[58] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_59 bl[59] br[59] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_60 bl[60] br[60] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_61 bl[61] br[61] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_62 bl[62] br[62] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_63 bl[63] br[63] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_64 bl[64] br[64] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_65 bl[65] br[65] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_66 bl[66] br[66] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_67 bl[67] br[67] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_68 bl[68] br[68] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_69 bl[69] br[69] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_70 bl[70] br[70] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_71 bl[71] br[71] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_72 bl[72] br[72] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_73 bl[73] br[73] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_74 bl[74] br[74] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_75 bl[75] br[75] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_76 bl[76] br[76] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_77 bl[77] br[77] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_78 bl[78] br[78] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_79 bl[79] br[79] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_80 bl[80] br[80] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_81 bl[81] br[81] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_82 bl[82] br[82] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_83 bl[83] br[83] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_84 bl[84] br[84] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_85 bl[85] br[85] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_86 bl[86] br[86] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_87 bl[87] br[87] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_88 bl[88] br[88] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_89 bl[89] br[89] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_90 bl[90] br[90] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_91 bl[91] br[91] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_92 bl[92] br[92] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_93 bl[93] br[93] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_94 bl[94] br[94] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_95 bl[95] br[95] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_96 bl[96] br[96] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_97 bl[97] br[97] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_98 bl[98] br[98] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_99 bl[99] br[99] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_100 bl[100] br[100] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_101 bl[101] br[101] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_102 bl[102] br[102] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_103 bl[103] br[103] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_104 bl[104] br[104] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_105 bl[105] br[105] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_106 bl[106] br[106] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_107 bl[107] br[107] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_108 bl[108] br[108] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_109 bl[109] br[109] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_110 bl[110] br[110] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_111 bl[111] br[111] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_112 bl[112] br[112] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_113 bl[113] br[113] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_114 bl[114] br[114] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_115 bl[115] br[115] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_116 bl[116] br[116] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_117 bl[117] br[117] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_118 bl[118] br[118] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_119 bl[119] br[119] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_120 bl[120] br[120] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_121 bl[121] br[121] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_122 bl[122] br[122] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_123 bl[123] br[123] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_124 bl[124] br[124] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_125 bl[125] br[125] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_126 bl[126] br[126] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_127 bl[127] br[127] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_128 bl[128] br[128] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_129 bl[129] br[129] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_130 bl[130] br[130] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_131 bl[131] br[131] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_132 bl[132] br[132] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_133 bl[133] br[133] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_134 bl[134] br[134] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_135 bl[135] br[135] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_136 bl[136] br[136] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_137 bl[137] br[137] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_138 bl[138] br[138] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_139 bl[139] br[139] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_140 bl[140] br[140] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_141 bl[141] br[141] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_142 bl[142] br[142] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_143 bl[143] br[143] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_144 bl[144] br[144] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_145 bl[145] br[145] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_146 bl[146] br[146] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_147 bl[147] br[147] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_148 bl[148] br[148] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_149 bl[149] br[149] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_150 bl[150] br[150] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_151 bl[151] br[151] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_152 bl[152] br[152] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_153 bl[153] br[153] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_154 bl[154] br[154] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_155 bl[155] br[155] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_156 bl[156] br[156] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_157 bl[157] br[157] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_158 bl[158] br[158] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_159 bl[159] br[159] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_160 bl[160] br[160] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_161 bl[161] br[161] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_162 bl[162] br[162] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_163 bl[163] br[163] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_164 bl[164] br[164] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_165 bl[165] br[165] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_166 bl[166] br[166] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_167 bl[167] br[167] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_168 bl[168] br[168] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_169 bl[169] br[169] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_170 bl[170] br[170] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_171 bl[171] br[171] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_172 bl[172] br[172] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_173 bl[173] br[173] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_174 bl[174] br[174] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_175 bl[175] br[175] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_176 bl[176] br[176] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_177 bl[177] br[177] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_178 bl[178] br[178] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_179 bl[179] br[179] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_180 bl[180] br[180] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_181 bl[181] br[181] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_182 bl[182] br[182] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_183 bl[183] br[183] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_184 bl[184] br[184] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_185 bl[185] br[185] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_186 bl[186] br[186] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_187 bl[187] br[187] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_188 bl[188] br[188] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_189 bl[189] br[189] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_190 bl[190] br[190] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_191 bl[191] br[191] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_192 bl[192] br[192] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_193 bl[193] br[193] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_194 bl[194] br[194] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_195 bl[195] br[195] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_196 bl[196] br[196] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_197 bl[197] br[197] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_198 bl[198] br[198] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_199 bl[199] br[199] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_200 bl[200] br[200] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_201 bl[201] br[201] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_202 bl[202] br[202] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_203 bl[203] br[203] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_204 bl[204] br[204] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_205 bl[205] br[205] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_206 bl[206] br[206] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_207 bl[207] br[207] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_208 bl[208] br[208] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_209 bl[209] br[209] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_210 bl[210] br[210] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_211 bl[211] br[211] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_212 bl[212] br[212] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_213 bl[213] br[213] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_214 bl[214] br[214] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_215 bl[215] br[215] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_216 bl[216] br[216] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_217 bl[217] br[217] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_218 bl[218] br[218] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_219 bl[219] br[219] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_220 bl[220] br[220] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_221 bl[221] br[221] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_222 bl[222] br[222] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_223 bl[223] br[223] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_224 bl[224] br[224] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_225 bl[225] br[225] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_226 bl[226] br[226] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_227 bl[227] br[227] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_228 bl[228] br[228] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_229 bl[229] br[229] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_230 bl[230] br[230] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_231 bl[231] br[231] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_232 bl[232] br[232] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_233 bl[233] br[233] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_234 bl[234] br[234] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_235 bl[235] br[235] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_236 bl[236] br[236] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_237 bl[237] br[237] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_238 bl[238] br[238] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_239 bl[239] br[239] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_240 bl[240] br[240] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_241 bl[241] br[241] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_242 bl[242] br[242] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_243 bl[243] br[243] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_244 bl[244] br[244] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_245 bl[245] br[245] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_246 bl[246] br[246] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_247 bl[247] br[247] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_248 bl[248] br[248] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_249 bl[249] br[249] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_250 bl[250] br[250] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_251 bl[251] br[251] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_252 bl[252] br[252] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_253 bl[253] br[253] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_254 bl[254] br[254] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_255 bl[255] br[255] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_26_0 bl[0] br[0] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_1 bl[1] br[1] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_2 bl[2] br[2] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_3 bl[3] br[3] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_4 bl[4] br[4] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_5 bl[5] br[5] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_6 bl[6] br[6] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_7 bl[7] br[7] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_8 bl[8] br[8] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_9 bl[9] br[9] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_10 bl[10] br[10] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_11 bl[11] br[11] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_12 bl[12] br[12] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_13 bl[13] br[13] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_14 bl[14] br[14] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_15 bl[15] br[15] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_16 bl[16] br[16] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_17 bl[17] br[17] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_18 bl[18] br[18] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_19 bl[19] br[19] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_20 bl[20] br[20] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_21 bl[21] br[21] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_22 bl[22] br[22] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_23 bl[23] br[23] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_24 bl[24] br[24] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_25 bl[25] br[25] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_26 bl[26] br[26] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_27 bl[27] br[27] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_28 bl[28] br[28] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_29 bl[29] br[29] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_30 bl[30] br[30] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_31 bl[31] br[31] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_32 bl[32] br[32] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_33 bl[33] br[33] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_34 bl[34] br[34] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_35 bl[35] br[35] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_36 bl[36] br[36] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_37 bl[37] br[37] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_38 bl[38] br[38] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_39 bl[39] br[39] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_40 bl[40] br[40] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_41 bl[41] br[41] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_42 bl[42] br[42] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_43 bl[43] br[43] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_44 bl[44] br[44] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_45 bl[45] br[45] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_46 bl[46] br[46] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_47 bl[47] br[47] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_48 bl[48] br[48] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_49 bl[49] br[49] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_50 bl[50] br[50] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_51 bl[51] br[51] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_52 bl[52] br[52] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_53 bl[53] br[53] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_54 bl[54] br[54] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_55 bl[55] br[55] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_56 bl[56] br[56] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_57 bl[57] br[57] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_58 bl[58] br[58] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_59 bl[59] br[59] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_60 bl[60] br[60] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_61 bl[61] br[61] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_62 bl[62] br[62] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_63 bl[63] br[63] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_64 bl[64] br[64] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_65 bl[65] br[65] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_66 bl[66] br[66] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_67 bl[67] br[67] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_68 bl[68] br[68] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_69 bl[69] br[69] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_70 bl[70] br[70] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_71 bl[71] br[71] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_72 bl[72] br[72] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_73 bl[73] br[73] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_74 bl[74] br[74] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_75 bl[75] br[75] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_76 bl[76] br[76] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_77 bl[77] br[77] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_78 bl[78] br[78] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_79 bl[79] br[79] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_80 bl[80] br[80] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_81 bl[81] br[81] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_82 bl[82] br[82] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_83 bl[83] br[83] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_84 bl[84] br[84] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_85 bl[85] br[85] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_86 bl[86] br[86] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_87 bl[87] br[87] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_88 bl[88] br[88] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_89 bl[89] br[89] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_90 bl[90] br[90] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_91 bl[91] br[91] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_92 bl[92] br[92] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_93 bl[93] br[93] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_94 bl[94] br[94] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_95 bl[95] br[95] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_96 bl[96] br[96] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_97 bl[97] br[97] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_98 bl[98] br[98] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_99 bl[99] br[99] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_100 bl[100] br[100] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_101 bl[101] br[101] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_102 bl[102] br[102] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_103 bl[103] br[103] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_104 bl[104] br[104] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_105 bl[105] br[105] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_106 bl[106] br[106] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_107 bl[107] br[107] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_108 bl[108] br[108] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_109 bl[109] br[109] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_110 bl[110] br[110] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_111 bl[111] br[111] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_112 bl[112] br[112] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_113 bl[113] br[113] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_114 bl[114] br[114] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_115 bl[115] br[115] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_116 bl[116] br[116] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_117 bl[117] br[117] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_118 bl[118] br[118] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_119 bl[119] br[119] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_120 bl[120] br[120] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_121 bl[121] br[121] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_122 bl[122] br[122] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_123 bl[123] br[123] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_124 bl[124] br[124] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_125 bl[125] br[125] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_126 bl[126] br[126] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_127 bl[127] br[127] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_128 bl[128] br[128] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_129 bl[129] br[129] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_130 bl[130] br[130] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_131 bl[131] br[131] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_132 bl[132] br[132] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_133 bl[133] br[133] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_134 bl[134] br[134] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_135 bl[135] br[135] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_136 bl[136] br[136] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_137 bl[137] br[137] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_138 bl[138] br[138] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_139 bl[139] br[139] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_140 bl[140] br[140] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_141 bl[141] br[141] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_142 bl[142] br[142] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_143 bl[143] br[143] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_144 bl[144] br[144] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_145 bl[145] br[145] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_146 bl[146] br[146] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_147 bl[147] br[147] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_148 bl[148] br[148] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_149 bl[149] br[149] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_150 bl[150] br[150] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_151 bl[151] br[151] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_152 bl[152] br[152] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_153 bl[153] br[153] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_154 bl[154] br[154] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_155 bl[155] br[155] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_156 bl[156] br[156] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_157 bl[157] br[157] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_158 bl[158] br[158] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_159 bl[159] br[159] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_160 bl[160] br[160] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_161 bl[161] br[161] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_162 bl[162] br[162] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_163 bl[163] br[163] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_164 bl[164] br[164] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_165 bl[165] br[165] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_166 bl[166] br[166] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_167 bl[167] br[167] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_168 bl[168] br[168] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_169 bl[169] br[169] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_170 bl[170] br[170] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_171 bl[171] br[171] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_172 bl[172] br[172] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_173 bl[173] br[173] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_174 bl[174] br[174] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_175 bl[175] br[175] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_176 bl[176] br[176] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_177 bl[177] br[177] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_178 bl[178] br[178] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_179 bl[179] br[179] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_180 bl[180] br[180] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_181 bl[181] br[181] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_182 bl[182] br[182] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_183 bl[183] br[183] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_184 bl[184] br[184] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_185 bl[185] br[185] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_186 bl[186] br[186] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_187 bl[187] br[187] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_188 bl[188] br[188] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_189 bl[189] br[189] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_190 bl[190] br[190] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_191 bl[191] br[191] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_192 bl[192] br[192] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_193 bl[193] br[193] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_194 bl[194] br[194] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_195 bl[195] br[195] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_196 bl[196] br[196] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_197 bl[197] br[197] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_198 bl[198] br[198] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_199 bl[199] br[199] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_200 bl[200] br[200] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_201 bl[201] br[201] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_202 bl[202] br[202] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_203 bl[203] br[203] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_204 bl[204] br[204] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_205 bl[205] br[205] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_206 bl[206] br[206] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_207 bl[207] br[207] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_208 bl[208] br[208] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_209 bl[209] br[209] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_210 bl[210] br[210] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_211 bl[211] br[211] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_212 bl[212] br[212] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_213 bl[213] br[213] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_214 bl[214] br[214] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_215 bl[215] br[215] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_216 bl[216] br[216] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_217 bl[217] br[217] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_218 bl[218] br[218] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_219 bl[219] br[219] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_220 bl[220] br[220] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_221 bl[221] br[221] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_222 bl[222] br[222] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_223 bl[223] br[223] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_224 bl[224] br[224] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_225 bl[225] br[225] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_226 bl[226] br[226] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_227 bl[227] br[227] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_228 bl[228] br[228] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_229 bl[229] br[229] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_230 bl[230] br[230] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_231 bl[231] br[231] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_232 bl[232] br[232] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_233 bl[233] br[233] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_234 bl[234] br[234] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_235 bl[235] br[235] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_236 bl[236] br[236] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_237 bl[237] br[237] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_238 bl[238] br[238] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_239 bl[239] br[239] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_240 bl[240] br[240] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_241 bl[241] br[241] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_242 bl[242] br[242] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_243 bl[243] br[243] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_244 bl[244] br[244] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_245 bl[245] br[245] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_246 bl[246] br[246] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_247 bl[247] br[247] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_248 bl[248] br[248] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_249 bl[249] br[249] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_250 bl[250] br[250] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_251 bl[251] br[251] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_252 bl[252] br[252] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_253 bl[253] br[253] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_254 bl[254] br[254] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_255 bl[255] br[255] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_27_0 bl[0] br[0] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_1 bl[1] br[1] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_2 bl[2] br[2] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_3 bl[3] br[3] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_4 bl[4] br[4] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_5 bl[5] br[5] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_6 bl[6] br[6] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_7 bl[7] br[7] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_8 bl[8] br[8] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_9 bl[9] br[9] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_10 bl[10] br[10] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_11 bl[11] br[11] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_12 bl[12] br[12] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_13 bl[13] br[13] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_14 bl[14] br[14] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_15 bl[15] br[15] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_16 bl[16] br[16] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_17 bl[17] br[17] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_18 bl[18] br[18] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_19 bl[19] br[19] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_20 bl[20] br[20] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_21 bl[21] br[21] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_22 bl[22] br[22] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_23 bl[23] br[23] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_24 bl[24] br[24] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_25 bl[25] br[25] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_26 bl[26] br[26] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_27 bl[27] br[27] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_28 bl[28] br[28] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_29 bl[29] br[29] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_30 bl[30] br[30] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_31 bl[31] br[31] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_32 bl[32] br[32] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_33 bl[33] br[33] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_34 bl[34] br[34] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_35 bl[35] br[35] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_36 bl[36] br[36] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_37 bl[37] br[37] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_38 bl[38] br[38] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_39 bl[39] br[39] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_40 bl[40] br[40] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_41 bl[41] br[41] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_42 bl[42] br[42] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_43 bl[43] br[43] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_44 bl[44] br[44] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_45 bl[45] br[45] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_46 bl[46] br[46] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_47 bl[47] br[47] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_48 bl[48] br[48] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_49 bl[49] br[49] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_50 bl[50] br[50] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_51 bl[51] br[51] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_52 bl[52] br[52] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_53 bl[53] br[53] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_54 bl[54] br[54] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_55 bl[55] br[55] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_56 bl[56] br[56] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_57 bl[57] br[57] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_58 bl[58] br[58] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_59 bl[59] br[59] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_60 bl[60] br[60] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_61 bl[61] br[61] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_62 bl[62] br[62] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_63 bl[63] br[63] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_64 bl[64] br[64] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_65 bl[65] br[65] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_66 bl[66] br[66] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_67 bl[67] br[67] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_68 bl[68] br[68] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_69 bl[69] br[69] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_70 bl[70] br[70] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_71 bl[71] br[71] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_72 bl[72] br[72] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_73 bl[73] br[73] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_74 bl[74] br[74] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_75 bl[75] br[75] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_76 bl[76] br[76] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_77 bl[77] br[77] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_78 bl[78] br[78] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_79 bl[79] br[79] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_80 bl[80] br[80] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_81 bl[81] br[81] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_82 bl[82] br[82] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_83 bl[83] br[83] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_84 bl[84] br[84] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_85 bl[85] br[85] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_86 bl[86] br[86] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_87 bl[87] br[87] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_88 bl[88] br[88] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_89 bl[89] br[89] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_90 bl[90] br[90] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_91 bl[91] br[91] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_92 bl[92] br[92] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_93 bl[93] br[93] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_94 bl[94] br[94] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_95 bl[95] br[95] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_96 bl[96] br[96] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_97 bl[97] br[97] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_98 bl[98] br[98] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_99 bl[99] br[99] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_100 bl[100] br[100] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_101 bl[101] br[101] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_102 bl[102] br[102] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_103 bl[103] br[103] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_104 bl[104] br[104] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_105 bl[105] br[105] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_106 bl[106] br[106] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_107 bl[107] br[107] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_108 bl[108] br[108] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_109 bl[109] br[109] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_110 bl[110] br[110] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_111 bl[111] br[111] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_112 bl[112] br[112] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_113 bl[113] br[113] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_114 bl[114] br[114] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_115 bl[115] br[115] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_116 bl[116] br[116] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_117 bl[117] br[117] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_118 bl[118] br[118] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_119 bl[119] br[119] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_120 bl[120] br[120] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_121 bl[121] br[121] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_122 bl[122] br[122] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_123 bl[123] br[123] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_124 bl[124] br[124] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_125 bl[125] br[125] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_126 bl[126] br[126] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_127 bl[127] br[127] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_128 bl[128] br[128] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_129 bl[129] br[129] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_130 bl[130] br[130] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_131 bl[131] br[131] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_132 bl[132] br[132] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_133 bl[133] br[133] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_134 bl[134] br[134] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_135 bl[135] br[135] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_136 bl[136] br[136] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_137 bl[137] br[137] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_138 bl[138] br[138] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_139 bl[139] br[139] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_140 bl[140] br[140] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_141 bl[141] br[141] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_142 bl[142] br[142] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_143 bl[143] br[143] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_144 bl[144] br[144] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_145 bl[145] br[145] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_146 bl[146] br[146] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_147 bl[147] br[147] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_148 bl[148] br[148] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_149 bl[149] br[149] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_150 bl[150] br[150] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_151 bl[151] br[151] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_152 bl[152] br[152] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_153 bl[153] br[153] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_154 bl[154] br[154] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_155 bl[155] br[155] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_156 bl[156] br[156] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_157 bl[157] br[157] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_158 bl[158] br[158] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_159 bl[159] br[159] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_160 bl[160] br[160] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_161 bl[161] br[161] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_162 bl[162] br[162] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_163 bl[163] br[163] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_164 bl[164] br[164] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_165 bl[165] br[165] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_166 bl[166] br[166] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_167 bl[167] br[167] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_168 bl[168] br[168] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_169 bl[169] br[169] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_170 bl[170] br[170] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_171 bl[171] br[171] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_172 bl[172] br[172] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_173 bl[173] br[173] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_174 bl[174] br[174] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_175 bl[175] br[175] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_176 bl[176] br[176] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_177 bl[177] br[177] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_178 bl[178] br[178] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_179 bl[179] br[179] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_180 bl[180] br[180] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_181 bl[181] br[181] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_182 bl[182] br[182] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_183 bl[183] br[183] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_184 bl[184] br[184] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_185 bl[185] br[185] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_186 bl[186] br[186] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_187 bl[187] br[187] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_188 bl[188] br[188] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_189 bl[189] br[189] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_190 bl[190] br[190] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_191 bl[191] br[191] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_192 bl[192] br[192] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_193 bl[193] br[193] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_194 bl[194] br[194] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_195 bl[195] br[195] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_196 bl[196] br[196] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_197 bl[197] br[197] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_198 bl[198] br[198] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_199 bl[199] br[199] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_200 bl[200] br[200] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_201 bl[201] br[201] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_202 bl[202] br[202] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_203 bl[203] br[203] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_204 bl[204] br[204] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_205 bl[205] br[205] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_206 bl[206] br[206] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_207 bl[207] br[207] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_208 bl[208] br[208] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_209 bl[209] br[209] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_210 bl[210] br[210] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_211 bl[211] br[211] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_212 bl[212] br[212] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_213 bl[213] br[213] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_214 bl[214] br[214] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_215 bl[215] br[215] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_216 bl[216] br[216] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_217 bl[217] br[217] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_218 bl[218] br[218] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_219 bl[219] br[219] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_220 bl[220] br[220] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_221 bl[221] br[221] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_222 bl[222] br[222] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_223 bl[223] br[223] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_224 bl[224] br[224] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_225 bl[225] br[225] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_226 bl[226] br[226] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_227 bl[227] br[227] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_228 bl[228] br[228] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_229 bl[229] br[229] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_230 bl[230] br[230] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_231 bl[231] br[231] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_232 bl[232] br[232] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_233 bl[233] br[233] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_234 bl[234] br[234] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_235 bl[235] br[235] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_236 bl[236] br[236] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_237 bl[237] br[237] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_238 bl[238] br[238] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_239 bl[239] br[239] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_240 bl[240] br[240] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_241 bl[241] br[241] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_242 bl[242] br[242] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_243 bl[243] br[243] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_244 bl[244] br[244] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_245 bl[245] br[245] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_246 bl[246] br[246] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_247 bl[247] br[247] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_248 bl[248] br[248] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_249 bl[249] br[249] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_250 bl[250] br[250] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_251 bl[251] br[251] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_252 bl[252] br[252] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_253 bl[253] br[253] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_254 bl[254] br[254] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_255 bl[255] br[255] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_28_0 bl[0] br[0] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_1 bl[1] br[1] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_2 bl[2] br[2] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_3 bl[3] br[3] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_4 bl[4] br[4] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_5 bl[5] br[5] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_6 bl[6] br[6] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_7 bl[7] br[7] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_8 bl[8] br[8] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_9 bl[9] br[9] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_10 bl[10] br[10] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_11 bl[11] br[11] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_12 bl[12] br[12] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_13 bl[13] br[13] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_14 bl[14] br[14] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_15 bl[15] br[15] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_16 bl[16] br[16] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_17 bl[17] br[17] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_18 bl[18] br[18] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_19 bl[19] br[19] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_20 bl[20] br[20] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_21 bl[21] br[21] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_22 bl[22] br[22] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_23 bl[23] br[23] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_24 bl[24] br[24] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_25 bl[25] br[25] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_26 bl[26] br[26] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_27 bl[27] br[27] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_28 bl[28] br[28] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_29 bl[29] br[29] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_30 bl[30] br[30] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_31 bl[31] br[31] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_32 bl[32] br[32] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_33 bl[33] br[33] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_34 bl[34] br[34] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_35 bl[35] br[35] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_36 bl[36] br[36] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_37 bl[37] br[37] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_38 bl[38] br[38] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_39 bl[39] br[39] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_40 bl[40] br[40] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_41 bl[41] br[41] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_42 bl[42] br[42] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_43 bl[43] br[43] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_44 bl[44] br[44] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_45 bl[45] br[45] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_46 bl[46] br[46] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_47 bl[47] br[47] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_48 bl[48] br[48] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_49 bl[49] br[49] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_50 bl[50] br[50] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_51 bl[51] br[51] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_52 bl[52] br[52] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_53 bl[53] br[53] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_54 bl[54] br[54] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_55 bl[55] br[55] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_56 bl[56] br[56] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_57 bl[57] br[57] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_58 bl[58] br[58] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_59 bl[59] br[59] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_60 bl[60] br[60] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_61 bl[61] br[61] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_62 bl[62] br[62] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_63 bl[63] br[63] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_64 bl[64] br[64] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_65 bl[65] br[65] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_66 bl[66] br[66] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_67 bl[67] br[67] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_68 bl[68] br[68] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_69 bl[69] br[69] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_70 bl[70] br[70] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_71 bl[71] br[71] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_72 bl[72] br[72] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_73 bl[73] br[73] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_74 bl[74] br[74] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_75 bl[75] br[75] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_76 bl[76] br[76] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_77 bl[77] br[77] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_78 bl[78] br[78] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_79 bl[79] br[79] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_80 bl[80] br[80] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_81 bl[81] br[81] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_82 bl[82] br[82] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_83 bl[83] br[83] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_84 bl[84] br[84] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_85 bl[85] br[85] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_86 bl[86] br[86] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_87 bl[87] br[87] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_88 bl[88] br[88] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_89 bl[89] br[89] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_90 bl[90] br[90] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_91 bl[91] br[91] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_92 bl[92] br[92] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_93 bl[93] br[93] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_94 bl[94] br[94] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_95 bl[95] br[95] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_96 bl[96] br[96] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_97 bl[97] br[97] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_98 bl[98] br[98] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_99 bl[99] br[99] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_100 bl[100] br[100] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_101 bl[101] br[101] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_102 bl[102] br[102] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_103 bl[103] br[103] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_104 bl[104] br[104] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_105 bl[105] br[105] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_106 bl[106] br[106] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_107 bl[107] br[107] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_108 bl[108] br[108] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_109 bl[109] br[109] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_110 bl[110] br[110] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_111 bl[111] br[111] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_112 bl[112] br[112] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_113 bl[113] br[113] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_114 bl[114] br[114] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_115 bl[115] br[115] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_116 bl[116] br[116] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_117 bl[117] br[117] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_118 bl[118] br[118] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_119 bl[119] br[119] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_120 bl[120] br[120] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_121 bl[121] br[121] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_122 bl[122] br[122] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_123 bl[123] br[123] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_124 bl[124] br[124] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_125 bl[125] br[125] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_126 bl[126] br[126] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_127 bl[127] br[127] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_128 bl[128] br[128] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_129 bl[129] br[129] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_130 bl[130] br[130] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_131 bl[131] br[131] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_132 bl[132] br[132] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_133 bl[133] br[133] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_134 bl[134] br[134] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_135 bl[135] br[135] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_136 bl[136] br[136] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_137 bl[137] br[137] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_138 bl[138] br[138] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_139 bl[139] br[139] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_140 bl[140] br[140] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_141 bl[141] br[141] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_142 bl[142] br[142] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_143 bl[143] br[143] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_144 bl[144] br[144] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_145 bl[145] br[145] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_146 bl[146] br[146] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_147 bl[147] br[147] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_148 bl[148] br[148] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_149 bl[149] br[149] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_150 bl[150] br[150] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_151 bl[151] br[151] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_152 bl[152] br[152] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_153 bl[153] br[153] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_154 bl[154] br[154] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_155 bl[155] br[155] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_156 bl[156] br[156] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_157 bl[157] br[157] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_158 bl[158] br[158] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_159 bl[159] br[159] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_160 bl[160] br[160] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_161 bl[161] br[161] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_162 bl[162] br[162] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_163 bl[163] br[163] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_164 bl[164] br[164] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_165 bl[165] br[165] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_166 bl[166] br[166] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_167 bl[167] br[167] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_168 bl[168] br[168] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_169 bl[169] br[169] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_170 bl[170] br[170] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_171 bl[171] br[171] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_172 bl[172] br[172] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_173 bl[173] br[173] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_174 bl[174] br[174] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_175 bl[175] br[175] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_176 bl[176] br[176] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_177 bl[177] br[177] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_178 bl[178] br[178] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_179 bl[179] br[179] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_180 bl[180] br[180] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_181 bl[181] br[181] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_182 bl[182] br[182] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_183 bl[183] br[183] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_184 bl[184] br[184] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_185 bl[185] br[185] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_186 bl[186] br[186] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_187 bl[187] br[187] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_188 bl[188] br[188] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_189 bl[189] br[189] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_190 bl[190] br[190] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_191 bl[191] br[191] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_192 bl[192] br[192] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_193 bl[193] br[193] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_194 bl[194] br[194] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_195 bl[195] br[195] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_196 bl[196] br[196] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_197 bl[197] br[197] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_198 bl[198] br[198] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_199 bl[199] br[199] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_200 bl[200] br[200] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_201 bl[201] br[201] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_202 bl[202] br[202] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_203 bl[203] br[203] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_204 bl[204] br[204] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_205 bl[205] br[205] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_206 bl[206] br[206] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_207 bl[207] br[207] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_208 bl[208] br[208] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_209 bl[209] br[209] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_210 bl[210] br[210] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_211 bl[211] br[211] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_212 bl[212] br[212] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_213 bl[213] br[213] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_214 bl[214] br[214] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_215 bl[215] br[215] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_216 bl[216] br[216] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_217 bl[217] br[217] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_218 bl[218] br[218] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_219 bl[219] br[219] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_220 bl[220] br[220] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_221 bl[221] br[221] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_222 bl[222] br[222] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_223 bl[223] br[223] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_224 bl[224] br[224] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_225 bl[225] br[225] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_226 bl[226] br[226] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_227 bl[227] br[227] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_228 bl[228] br[228] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_229 bl[229] br[229] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_230 bl[230] br[230] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_231 bl[231] br[231] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_232 bl[232] br[232] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_233 bl[233] br[233] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_234 bl[234] br[234] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_235 bl[235] br[235] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_236 bl[236] br[236] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_237 bl[237] br[237] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_238 bl[238] br[238] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_239 bl[239] br[239] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_240 bl[240] br[240] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_241 bl[241] br[241] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_242 bl[242] br[242] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_243 bl[243] br[243] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_244 bl[244] br[244] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_245 bl[245] br[245] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_246 bl[246] br[246] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_247 bl[247] br[247] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_248 bl[248] br[248] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_249 bl[249] br[249] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_250 bl[250] br[250] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_251 bl[251] br[251] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_252 bl[252] br[252] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_253 bl[253] br[253] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_254 bl[254] br[254] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_255 bl[255] br[255] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_29_0 bl[0] br[0] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_1 bl[1] br[1] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_2 bl[2] br[2] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_3 bl[3] br[3] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_4 bl[4] br[4] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_5 bl[5] br[5] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_6 bl[6] br[6] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_7 bl[7] br[7] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_8 bl[8] br[8] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_9 bl[9] br[9] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_10 bl[10] br[10] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_11 bl[11] br[11] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_12 bl[12] br[12] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_13 bl[13] br[13] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_14 bl[14] br[14] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_15 bl[15] br[15] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_16 bl[16] br[16] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_17 bl[17] br[17] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_18 bl[18] br[18] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_19 bl[19] br[19] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_20 bl[20] br[20] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_21 bl[21] br[21] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_22 bl[22] br[22] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_23 bl[23] br[23] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_24 bl[24] br[24] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_25 bl[25] br[25] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_26 bl[26] br[26] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_27 bl[27] br[27] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_28 bl[28] br[28] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_29 bl[29] br[29] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_30 bl[30] br[30] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_31 bl[31] br[31] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_32 bl[32] br[32] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_33 bl[33] br[33] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_34 bl[34] br[34] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_35 bl[35] br[35] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_36 bl[36] br[36] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_37 bl[37] br[37] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_38 bl[38] br[38] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_39 bl[39] br[39] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_40 bl[40] br[40] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_41 bl[41] br[41] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_42 bl[42] br[42] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_43 bl[43] br[43] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_44 bl[44] br[44] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_45 bl[45] br[45] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_46 bl[46] br[46] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_47 bl[47] br[47] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_48 bl[48] br[48] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_49 bl[49] br[49] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_50 bl[50] br[50] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_51 bl[51] br[51] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_52 bl[52] br[52] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_53 bl[53] br[53] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_54 bl[54] br[54] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_55 bl[55] br[55] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_56 bl[56] br[56] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_57 bl[57] br[57] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_58 bl[58] br[58] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_59 bl[59] br[59] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_60 bl[60] br[60] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_61 bl[61] br[61] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_62 bl[62] br[62] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_63 bl[63] br[63] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_64 bl[64] br[64] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_65 bl[65] br[65] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_66 bl[66] br[66] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_67 bl[67] br[67] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_68 bl[68] br[68] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_69 bl[69] br[69] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_70 bl[70] br[70] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_71 bl[71] br[71] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_72 bl[72] br[72] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_73 bl[73] br[73] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_74 bl[74] br[74] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_75 bl[75] br[75] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_76 bl[76] br[76] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_77 bl[77] br[77] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_78 bl[78] br[78] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_79 bl[79] br[79] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_80 bl[80] br[80] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_81 bl[81] br[81] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_82 bl[82] br[82] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_83 bl[83] br[83] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_84 bl[84] br[84] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_85 bl[85] br[85] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_86 bl[86] br[86] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_87 bl[87] br[87] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_88 bl[88] br[88] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_89 bl[89] br[89] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_90 bl[90] br[90] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_91 bl[91] br[91] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_92 bl[92] br[92] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_93 bl[93] br[93] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_94 bl[94] br[94] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_95 bl[95] br[95] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_96 bl[96] br[96] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_97 bl[97] br[97] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_98 bl[98] br[98] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_99 bl[99] br[99] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_100 bl[100] br[100] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_101 bl[101] br[101] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_102 bl[102] br[102] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_103 bl[103] br[103] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_104 bl[104] br[104] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_105 bl[105] br[105] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_106 bl[106] br[106] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_107 bl[107] br[107] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_108 bl[108] br[108] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_109 bl[109] br[109] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_110 bl[110] br[110] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_111 bl[111] br[111] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_112 bl[112] br[112] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_113 bl[113] br[113] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_114 bl[114] br[114] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_115 bl[115] br[115] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_116 bl[116] br[116] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_117 bl[117] br[117] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_118 bl[118] br[118] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_119 bl[119] br[119] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_120 bl[120] br[120] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_121 bl[121] br[121] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_122 bl[122] br[122] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_123 bl[123] br[123] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_124 bl[124] br[124] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_125 bl[125] br[125] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_126 bl[126] br[126] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_127 bl[127] br[127] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_128 bl[128] br[128] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_129 bl[129] br[129] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_130 bl[130] br[130] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_131 bl[131] br[131] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_132 bl[132] br[132] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_133 bl[133] br[133] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_134 bl[134] br[134] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_135 bl[135] br[135] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_136 bl[136] br[136] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_137 bl[137] br[137] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_138 bl[138] br[138] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_139 bl[139] br[139] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_140 bl[140] br[140] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_141 bl[141] br[141] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_142 bl[142] br[142] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_143 bl[143] br[143] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_144 bl[144] br[144] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_145 bl[145] br[145] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_146 bl[146] br[146] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_147 bl[147] br[147] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_148 bl[148] br[148] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_149 bl[149] br[149] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_150 bl[150] br[150] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_151 bl[151] br[151] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_152 bl[152] br[152] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_153 bl[153] br[153] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_154 bl[154] br[154] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_155 bl[155] br[155] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_156 bl[156] br[156] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_157 bl[157] br[157] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_158 bl[158] br[158] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_159 bl[159] br[159] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_160 bl[160] br[160] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_161 bl[161] br[161] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_162 bl[162] br[162] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_163 bl[163] br[163] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_164 bl[164] br[164] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_165 bl[165] br[165] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_166 bl[166] br[166] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_167 bl[167] br[167] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_168 bl[168] br[168] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_169 bl[169] br[169] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_170 bl[170] br[170] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_171 bl[171] br[171] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_172 bl[172] br[172] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_173 bl[173] br[173] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_174 bl[174] br[174] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_175 bl[175] br[175] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_176 bl[176] br[176] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_177 bl[177] br[177] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_178 bl[178] br[178] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_179 bl[179] br[179] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_180 bl[180] br[180] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_181 bl[181] br[181] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_182 bl[182] br[182] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_183 bl[183] br[183] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_184 bl[184] br[184] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_185 bl[185] br[185] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_186 bl[186] br[186] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_187 bl[187] br[187] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_188 bl[188] br[188] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_189 bl[189] br[189] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_190 bl[190] br[190] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_191 bl[191] br[191] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_192 bl[192] br[192] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_193 bl[193] br[193] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_194 bl[194] br[194] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_195 bl[195] br[195] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_196 bl[196] br[196] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_197 bl[197] br[197] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_198 bl[198] br[198] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_199 bl[199] br[199] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_200 bl[200] br[200] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_201 bl[201] br[201] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_202 bl[202] br[202] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_203 bl[203] br[203] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_204 bl[204] br[204] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_205 bl[205] br[205] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_206 bl[206] br[206] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_207 bl[207] br[207] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_208 bl[208] br[208] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_209 bl[209] br[209] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_210 bl[210] br[210] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_211 bl[211] br[211] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_212 bl[212] br[212] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_213 bl[213] br[213] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_214 bl[214] br[214] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_215 bl[215] br[215] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_216 bl[216] br[216] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_217 bl[217] br[217] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_218 bl[218] br[218] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_219 bl[219] br[219] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_220 bl[220] br[220] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_221 bl[221] br[221] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_222 bl[222] br[222] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_223 bl[223] br[223] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_224 bl[224] br[224] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_225 bl[225] br[225] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_226 bl[226] br[226] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_227 bl[227] br[227] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_228 bl[228] br[228] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_229 bl[229] br[229] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_230 bl[230] br[230] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_231 bl[231] br[231] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_232 bl[232] br[232] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_233 bl[233] br[233] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_234 bl[234] br[234] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_235 bl[235] br[235] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_236 bl[236] br[236] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_237 bl[237] br[237] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_238 bl[238] br[238] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_239 bl[239] br[239] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_240 bl[240] br[240] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_241 bl[241] br[241] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_242 bl[242] br[242] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_243 bl[243] br[243] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_244 bl[244] br[244] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_245 bl[245] br[245] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_246 bl[246] br[246] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_247 bl[247] br[247] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_248 bl[248] br[248] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_249 bl[249] br[249] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_250 bl[250] br[250] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_251 bl[251] br[251] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_252 bl[252] br[252] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_253 bl[253] br[253] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_254 bl[254] br[254] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_255 bl[255] br[255] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_30_0 bl[0] br[0] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_1 bl[1] br[1] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_2 bl[2] br[2] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_3 bl[3] br[3] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_4 bl[4] br[4] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_5 bl[5] br[5] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_6 bl[6] br[6] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_7 bl[7] br[7] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_8 bl[8] br[8] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_9 bl[9] br[9] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_10 bl[10] br[10] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_11 bl[11] br[11] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_12 bl[12] br[12] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_13 bl[13] br[13] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_14 bl[14] br[14] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_15 bl[15] br[15] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_16 bl[16] br[16] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_17 bl[17] br[17] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_18 bl[18] br[18] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_19 bl[19] br[19] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_20 bl[20] br[20] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_21 bl[21] br[21] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_22 bl[22] br[22] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_23 bl[23] br[23] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_24 bl[24] br[24] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_25 bl[25] br[25] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_26 bl[26] br[26] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_27 bl[27] br[27] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_28 bl[28] br[28] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_29 bl[29] br[29] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_30 bl[30] br[30] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_31 bl[31] br[31] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_32 bl[32] br[32] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_33 bl[33] br[33] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_34 bl[34] br[34] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_35 bl[35] br[35] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_36 bl[36] br[36] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_37 bl[37] br[37] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_38 bl[38] br[38] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_39 bl[39] br[39] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_40 bl[40] br[40] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_41 bl[41] br[41] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_42 bl[42] br[42] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_43 bl[43] br[43] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_44 bl[44] br[44] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_45 bl[45] br[45] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_46 bl[46] br[46] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_47 bl[47] br[47] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_48 bl[48] br[48] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_49 bl[49] br[49] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_50 bl[50] br[50] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_51 bl[51] br[51] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_52 bl[52] br[52] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_53 bl[53] br[53] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_54 bl[54] br[54] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_55 bl[55] br[55] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_56 bl[56] br[56] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_57 bl[57] br[57] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_58 bl[58] br[58] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_59 bl[59] br[59] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_60 bl[60] br[60] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_61 bl[61] br[61] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_62 bl[62] br[62] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_63 bl[63] br[63] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_64 bl[64] br[64] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_65 bl[65] br[65] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_66 bl[66] br[66] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_67 bl[67] br[67] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_68 bl[68] br[68] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_69 bl[69] br[69] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_70 bl[70] br[70] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_71 bl[71] br[71] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_72 bl[72] br[72] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_73 bl[73] br[73] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_74 bl[74] br[74] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_75 bl[75] br[75] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_76 bl[76] br[76] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_77 bl[77] br[77] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_78 bl[78] br[78] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_79 bl[79] br[79] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_80 bl[80] br[80] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_81 bl[81] br[81] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_82 bl[82] br[82] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_83 bl[83] br[83] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_84 bl[84] br[84] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_85 bl[85] br[85] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_86 bl[86] br[86] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_87 bl[87] br[87] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_88 bl[88] br[88] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_89 bl[89] br[89] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_90 bl[90] br[90] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_91 bl[91] br[91] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_92 bl[92] br[92] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_93 bl[93] br[93] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_94 bl[94] br[94] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_95 bl[95] br[95] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_96 bl[96] br[96] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_97 bl[97] br[97] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_98 bl[98] br[98] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_99 bl[99] br[99] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_100 bl[100] br[100] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_101 bl[101] br[101] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_102 bl[102] br[102] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_103 bl[103] br[103] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_104 bl[104] br[104] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_105 bl[105] br[105] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_106 bl[106] br[106] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_107 bl[107] br[107] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_108 bl[108] br[108] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_109 bl[109] br[109] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_110 bl[110] br[110] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_111 bl[111] br[111] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_112 bl[112] br[112] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_113 bl[113] br[113] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_114 bl[114] br[114] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_115 bl[115] br[115] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_116 bl[116] br[116] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_117 bl[117] br[117] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_118 bl[118] br[118] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_119 bl[119] br[119] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_120 bl[120] br[120] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_121 bl[121] br[121] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_122 bl[122] br[122] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_123 bl[123] br[123] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_124 bl[124] br[124] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_125 bl[125] br[125] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_126 bl[126] br[126] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_127 bl[127] br[127] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_128 bl[128] br[128] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_129 bl[129] br[129] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_130 bl[130] br[130] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_131 bl[131] br[131] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_132 bl[132] br[132] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_133 bl[133] br[133] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_134 bl[134] br[134] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_135 bl[135] br[135] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_136 bl[136] br[136] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_137 bl[137] br[137] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_138 bl[138] br[138] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_139 bl[139] br[139] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_140 bl[140] br[140] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_141 bl[141] br[141] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_142 bl[142] br[142] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_143 bl[143] br[143] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_144 bl[144] br[144] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_145 bl[145] br[145] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_146 bl[146] br[146] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_147 bl[147] br[147] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_148 bl[148] br[148] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_149 bl[149] br[149] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_150 bl[150] br[150] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_151 bl[151] br[151] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_152 bl[152] br[152] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_153 bl[153] br[153] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_154 bl[154] br[154] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_155 bl[155] br[155] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_156 bl[156] br[156] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_157 bl[157] br[157] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_158 bl[158] br[158] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_159 bl[159] br[159] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_160 bl[160] br[160] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_161 bl[161] br[161] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_162 bl[162] br[162] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_163 bl[163] br[163] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_164 bl[164] br[164] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_165 bl[165] br[165] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_166 bl[166] br[166] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_167 bl[167] br[167] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_168 bl[168] br[168] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_169 bl[169] br[169] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_170 bl[170] br[170] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_171 bl[171] br[171] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_172 bl[172] br[172] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_173 bl[173] br[173] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_174 bl[174] br[174] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_175 bl[175] br[175] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_176 bl[176] br[176] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_177 bl[177] br[177] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_178 bl[178] br[178] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_179 bl[179] br[179] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_180 bl[180] br[180] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_181 bl[181] br[181] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_182 bl[182] br[182] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_183 bl[183] br[183] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_184 bl[184] br[184] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_185 bl[185] br[185] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_186 bl[186] br[186] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_187 bl[187] br[187] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_188 bl[188] br[188] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_189 bl[189] br[189] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_190 bl[190] br[190] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_191 bl[191] br[191] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_192 bl[192] br[192] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_193 bl[193] br[193] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_194 bl[194] br[194] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_195 bl[195] br[195] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_196 bl[196] br[196] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_197 bl[197] br[197] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_198 bl[198] br[198] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_199 bl[199] br[199] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_200 bl[200] br[200] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_201 bl[201] br[201] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_202 bl[202] br[202] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_203 bl[203] br[203] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_204 bl[204] br[204] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_205 bl[205] br[205] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_206 bl[206] br[206] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_207 bl[207] br[207] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_208 bl[208] br[208] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_209 bl[209] br[209] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_210 bl[210] br[210] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_211 bl[211] br[211] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_212 bl[212] br[212] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_213 bl[213] br[213] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_214 bl[214] br[214] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_215 bl[215] br[215] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_216 bl[216] br[216] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_217 bl[217] br[217] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_218 bl[218] br[218] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_219 bl[219] br[219] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_220 bl[220] br[220] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_221 bl[221] br[221] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_222 bl[222] br[222] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_223 bl[223] br[223] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_224 bl[224] br[224] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_225 bl[225] br[225] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_226 bl[226] br[226] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_227 bl[227] br[227] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_228 bl[228] br[228] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_229 bl[229] br[229] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_230 bl[230] br[230] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_231 bl[231] br[231] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_232 bl[232] br[232] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_233 bl[233] br[233] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_234 bl[234] br[234] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_235 bl[235] br[235] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_236 bl[236] br[236] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_237 bl[237] br[237] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_238 bl[238] br[238] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_239 bl[239] br[239] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_240 bl[240] br[240] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_241 bl[241] br[241] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_242 bl[242] br[242] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_243 bl[243] br[243] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_244 bl[244] br[244] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_245 bl[245] br[245] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_246 bl[246] br[246] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_247 bl[247] br[247] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_248 bl[248] br[248] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_249 bl[249] br[249] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_250 bl[250] br[250] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_251 bl[251] br[251] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_252 bl[252] br[252] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_253 bl[253] br[253] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_254 bl[254] br[254] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_255 bl[255] br[255] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_31_0 bl[0] br[0] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_1 bl[1] br[1] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_2 bl[2] br[2] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_3 bl[3] br[3] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_4 bl[4] br[4] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_5 bl[5] br[5] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_6 bl[6] br[6] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_7 bl[7] br[7] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_8 bl[8] br[8] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_9 bl[9] br[9] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_10 bl[10] br[10] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_11 bl[11] br[11] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_12 bl[12] br[12] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_13 bl[13] br[13] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_14 bl[14] br[14] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_15 bl[15] br[15] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_16 bl[16] br[16] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_17 bl[17] br[17] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_18 bl[18] br[18] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_19 bl[19] br[19] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_20 bl[20] br[20] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_21 bl[21] br[21] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_22 bl[22] br[22] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_23 bl[23] br[23] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_24 bl[24] br[24] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_25 bl[25] br[25] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_26 bl[26] br[26] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_27 bl[27] br[27] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_28 bl[28] br[28] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_29 bl[29] br[29] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_30 bl[30] br[30] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_31 bl[31] br[31] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_32 bl[32] br[32] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_33 bl[33] br[33] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_34 bl[34] br[34] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_35 bl[35] br[35] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_36 bl[36] br[36] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_37 bl[37] br[37] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_38 bl[38] br[38] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_39 bl[39] br[39] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_40 bl[40] br[40] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_41 bl[41] br[41] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_42 bl[42] br[42] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_43 bl[43] br[43] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_44 bl[44] br[44] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_45 bl[45] br[45] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_46 bl[46] br[46] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_47 bl[47] br[47] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_48 bl[48] br[48] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_49 bl[49] br[49] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_50 bl[50] br[50] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_51 bl[51] br[51] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_52 bl[52] br[52] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_53 bl[53] br[53] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_54 bl[54] br[54] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_55 bl[55] br[55] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_56 bl[56] br[56] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_57 bl[57] br[57] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_58 bl[58] br[58] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_59 bl[59] br[59] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_60 bl[60] br[60] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_61 bl[61] br[61] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_62 bl[62] br[62] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_63 bl[63] br[63] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_64 bl[64] br[64] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_65 bl[65] br[65] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_66 bl[66] br[66] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_67 bl[67] br[67] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_68 bl[68] br[68] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_69 bl[69] br[69] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_70 bl[70] br[70] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_71 bl[71] br[71] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_72 bl[72] br[72] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_73 bl[73] br[73] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_74 bl[74] br[74] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_75 bl[75] br[75] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_76 bl[76] br[76] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_77 bl[77] br[77] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_78 bl[78] br[78] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_79 bl[79] br[79] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_80 bl[80] br[80] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_81 bl[81] br[81] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_82 bl[82] br[82] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_83 bl[83] br[83] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_84 bl[84] br[84] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_85 bl[85] br[85] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_86 bl[86] br[86] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_87 bl[87] br[87] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_88 bl[88] br[88] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_89 bl[89] br[89] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_90 bl[90] br[90] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_91 bl[91] br[91] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_92 bl[92] br[92] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_93 bl[93] br[93] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_94 bl[94] br[94] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_95 bl[95] br[95] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_96 bl[96] br[96] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_97 bl[97] br[97] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_98 bl[98] br[98] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_99 bl[99] br[99] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_100 bl[100] br[100] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_101 bl[101] br[101] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_102 bl[102] br[102] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_103 bl[103] br[103] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_104 bl[104] br[104] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_105 bl[105] br[105] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_106 bl[106] br[106] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_107 bl[107] br[107] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_108 bl[108] br[108] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_109 bl[109] br[109] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_110 bl[110] br[110] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_111 bl[111] br[111] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_112 bl[112] br[112] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_113 bl[113] br[113] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_114 bl[114] br[114] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_115 bl[115] br[115] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_116 bl[116] br[116] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_117 bl[117] br[117] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_118 bl[118] br[118] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_119 bl[119] br[119] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_120 bl[120] br[120] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_121 bl[121] br[121] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_122 bl[122] br[122] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_123 bl[123] br[123] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_124 bl[124] br[124] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_125 bl[125] br[125] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_126 bl[126] br[126] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_127 bl[127] br[127] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_128 bl[128] br[128] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_129 bl[129] br[129] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_130 bl[130] br[130] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_131 bl[131] br[131] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_132 bl[132] br[132] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_133 bl[133] br[133] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_134 bl[134] br[134] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_135 bl[135] br[135] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_136 bl[136] br[136] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_137 bl[137] br[137] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_138 bl[138] br[138] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_139 bl[139] br[139] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_140 bl[140] br[140] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_141 bl[141] br[141] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_142 bl[142] br[142] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_143 bl[143] br[143] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_144 bl[144] br[144] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_145 bl[145] br[145] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_146 bl[146] br[146] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_147 bl[147] br[147] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_148 bl[148] br[148] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_149 bl[149] br[149] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_150 bl[150] br[150] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_151 bl[151] br[151] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_152 bl[152] br[152] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_153 bl[153] br[153] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_154 bl[154] br[154] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_155 bl[155] br[155] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_156 bl[156] br[156] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_157 bl[157] br[157] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_158 bl[158] br[158] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_159 bl[159] br[159] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_160 bl[160] br[160] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_161 bl[161] br[161] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_162 bl[162] br[162] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_163 bl[163] br[163] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_164 bl[164] br[164] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_165 bl[165] br[165] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_166 bl[166] br[166] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_167 bl[167] br[167] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_168 bl[168] br[168] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_169 bl[169] br[169] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_170 bl[170] br[170] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_171 bl[171] br[171] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_172 bl[172] br[172] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_173 bl[173] br[173] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_174 bl[174] br[174] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_175 bl[175] br[175] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_176 bl[176] br[176] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_177 bl[177] br[177] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_178 bl[178] br[178] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_179 bl[179] br[179] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_180 bl[180] br[180] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_181 bl[181] br[181] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_182 bl[182] br[182] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_183 bl[183] br[183] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_184 bl[184] br[184] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_185 bl[185] br[185] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_186 bl[186] br[186] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_187 bl[187] br[187] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_188 bl[188] br[188] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_189 bl[189] br[189] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_190 bl[190] br[190] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_191 bl[191] br[191] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_192 bl[192] br[192] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_193 bl[193] br[193] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_194 bl[194] br[194] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_195 bl[195] br[195] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_196 bl[196] br[196] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_197 bl[197] br[197] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_198 bl[198] br[198] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_199 bl[199] br[199] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_200 bl[200] br[200] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_201 bl[201] br[201] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_202 bl[202] br[202] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_203 bl[203] br[203] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_204 bl[204] br[204] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_205 bl[205] br[205] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_206 bl[206] br[206] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_207 bl[207] br[207] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_208 bl[208] br[208] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_209 bl[209] br[209] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_210 bl[210] br[210] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_211 bl[211] br[211] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_212 bl[212] br[212] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_213 bl[213] br[213] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_214 bl[214] br[214] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_215 bl[215] br[215] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_216 bl[216] br[216] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_217 bl[217] br[217] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_218 bl[218] br[218] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_219 bl[219] br[219] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_220 bl[220] br[220] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_221 bl[221] br[221] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_222 bl[222] br[222] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_223 bl[223] br[223] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_224 bl[224] br[224] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_225 bl[225] br[225] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_226 bl[226] br[226] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_227 bl[227] br[227] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_228 bl[228] br[228] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_229 bl[229] br[229] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_230 bl[230] br[230] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_231 bl[231] br[231] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_232 bl[232] br[232] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_233 bl[233] br[233] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_234 bl[234] br[234] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_235 bl[235] br[235] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_236 bl[236] br[236] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_237 bl[237] br[237] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_238 bl[238] br[238] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_239 bl[239] br[239] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_240 bl[240] br[240] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_241 bl[241] br[241] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_242 bl[242] br[242] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_243 bl[243] br[243] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_244 bl[244] br[244] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_245 bl[245] br[245] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_246 bl[246] br[246] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_247 bl[247] br[247] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_248 bl[248] br[248] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_249 bl[249] br[249] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_250 bl[250] br[250] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_251 bl[251] br[251] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_252 bl[252] br[252] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_253 bl[253] br[253] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_254 bl[254] br[254] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_255 bl[255] br[255] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_32_0 bl[0] br[0] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_1 bl[1] br[1] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_2 bl[2] br[2] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_3 bl[3] br[3] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_4 bl[4] br[4] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_5 bl[5] br[5] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_6 bl[6] br[6] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_7 bl[7] br[7] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_8 bl[8] br[8] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_9 bl[9] br[9] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_10 bl[10] br[10] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_11 bl[11] br[11] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_12 bl[12] br[12] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_13 bl[13] br[13] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_14 bl[14] br[14] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_15 bl[15] br[15] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_16 bl[16] br[16] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_17 bl[17] br[17] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_18 bl[18] br[18] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_19 bl[19] br[19] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_20 bl[20] br[20] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_21 bl[21] br[21] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_22 bl[22] br[22] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_23 bl[23] br[23] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_24 bl[24] br[24] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_25 bl[25] br[25] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_26 bl[26] br[26] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_27 bl[27] br[27] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_28 bl[28] br[28] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_29 bl[29] br[29] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_30 bl[30] br[30] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_31 bl[31] br[31] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_32 bl[32] br[32] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_33 bl[33] br[33] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_34 bl[34] br[34] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_35 bl[35] br[35] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_36 bl[36] br[36] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_37 bl[37] br[37] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_38 bl[38] br[38] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_39 bl[39] br[39] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_40 bl[40] br[40] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_41 bl[41] br[41] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_42 bl[42] br[42] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_43 bl[43] br[43] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_44 bl[44] br[44] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_45 bl[45] br[45] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_46 bl[46] br[46] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_47 bl[47] br[47] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_48 bl[48] br[48] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_49 bl[49] br[49] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_50 bl[50] br[50] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_51 bl[51] br[51] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_52 bl[52] br[52] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_53 bl[53] br[53] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_54 bl[54] br[54] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_55 bl[55] br[55] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_56 bl[56] br[56] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_57 bl[57] br[57] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_58 bl[58] br[58] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_59 bl[59] br[59] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_60 bl[60] br[60] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_61 bl[61] br[61] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_62 bl[62] br[62] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_63 bl[63] br[63] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_64 bl[64] br[64] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_65 bl[65] br[65] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_66 bl[66] br[66] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_67 bl[67] br[67] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_68 bl[68] br[68] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_69 bl[69] br[69] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_70 bl[70] br[70] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_71 bl[71] br[71] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_72 bl[72] br[72] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_73 bl[73] br[73] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_74 bl[74] br[74] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_75 bl[75] br[75] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_76 bl[76] br[76] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_77 bl[77] br[77] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_78 bl[78] br[78] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_79 bl[79] br[79] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_80 bl[80] br[80] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_81 bl[81] br[81] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_82 bl[82] br[82] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_83 bl[83] br[83] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_84 bl[84] br[84] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_85 bl[85] br[85] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_86 bl[86] br[86] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_87 bl[87] br[87] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_88 bl[88] br[88] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_89 bl[89] br[89] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_90 bl[90] br[90] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_91 bl[91] br[91] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_92 bl[92] br[92] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_93 bl[93] br[93] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_94 bl[94] br[94] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_95 bl[95] br[95] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_96 bl[96] br[96] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_97 bl[97] br[97] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_98 bl[98] br[98] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_99 bl[99] br[99] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_100 bl[100] br[100] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_101 bl[101] br[101] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_102 bl[102] br[102] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_103 bl[103] br[103] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_104 bl[104] br[104] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_105 bl[105] br[105] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_106 bl[106] br[106] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_107 bl[107] br[107] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_108 bl[108] br[108] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_109 bl[109] br[109] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_110 bl[110] br[110] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_111 bl[111] br[111] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_112 bl[112] br[112] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_113 bl[113] br[113] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_114 bl[114] br[114] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_115 bl[115] br[115] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_116 bl[116] br[116] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_117 bl[117] br[117] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_118 bl[118] br[118] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_119 bl[119] br[119] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_120 bl[120] br[120] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_121 bl[121] br[121] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_122 bl[122] br[122] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_123 bl[123] br[123] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_124 bl[124] br[124] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_125 bl[125] br[125] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_126 bl[126] br[126] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_127 bl[127] br[127] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_128 bl[128] br[128] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_129 bl[129] br[129] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_130 bl[130] br[130] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_131 bl[131] br[131] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_132 bl[132] br[132] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_133 bl[133] br[133] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_134 bl[134] br[134] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_135 bl[135] br[135] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_136 bl[136] br[136] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_137 bl[137] br[137] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_138 bl[138] br[138] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_139 bl[139] br[139] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_140 bl[140] br[140] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_141 bl[141] br[141] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_142 bl[142] br[142] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_143 bl[143] br[143] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_144 bl[144] br[144] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_145 bl[145] br[145] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_146 bl[146] br[146] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_147 bl[147] br[147] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_148 bl[148] br[148] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_149 bl[149] br[149] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_150 bl[150] br[150] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_151 bl[151] br[151] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_152 bl[152] br[152] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_153 bl[153] br[153] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_154 bl[154] br[154] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_155 bl[155] br[155] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_156 bl[156] br[156] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_157 bl[157] br[157] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_158 bl[158] br[158] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_159 bl[159] br[159] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_160 bl[160] br[160] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_161 bl[161] br[161] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_162 bl[162] br[162] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_163 bl[163] br[163] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_164 bl[164] br[164] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_165 bl[165] br[165] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_166 bl[166] br[166] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_167 bl[167] br[167] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_168 bl[168] br[168] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_169 bl[169] br[169] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_170 bl[170] br[170] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_171 bl[171] br[171] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_172 bl[172] br[172] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_173 bl[173] br[173] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_174 bl[174] br[174] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_175 bl[175] br[175] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_176 bl[176] br[176] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_177 bl[177] br[177] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_178 bl[178] br[178] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_179 bl[179] br[179] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_180 bl[180] br[180] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_181 bl[181] br[181] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_182 bl[182] br[182] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_183 bl[183] br[183] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_184 bl[184] br[184] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_185 bl[185] br[185] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_186 bl[186] br[186] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_187 bl[187] br[187] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_188 bl[188] br[188] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_189 bl[189] br[189] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_190 bl[190] br[190] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_191 bl[191] br[191] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_192 bl[192] br[192] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_193 bl[193] br[193] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_194 bl[194] br[194] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_195 bl[195] br[195] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_196 bl[196] br[196] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_197 bl[197] br[197] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_198 bl[198] br[198] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_199 bl[199] br[199] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_200 bl[200] br[200] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_201 bl[201] br[201] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_202 bl[202] br[202] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_203 bl[203] br[203] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_204 bl[204] br[204] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_205 bl[205] br[205] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_206 bl[206] br[206] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_207 bl[207] br[207] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_208 bl[208] br[208] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_209 bl[209] br[209] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_210 bl[210] br[210] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_211 bl[211] br[211] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_212 bl[212] br[212] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_213 bl[213] br[213] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_214 bl[214] br[214] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_215 bl[215] br[215] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_216 bl[216] br[216] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_217 bl[217] br[217] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_218 bl[218] br[218] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_219 bl[219] br[219] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_220 bl[220] br[220] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_221 bl[221] br[221] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_222 bl[222] br[222] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_223 bl[223] br[223] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_224 bl[224] br[224] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_225 bl[225] br[225] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_226 bl[226] br[226] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_227 bl[227] br[227] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_228 bl[228] br[228] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_229 bl[229] br[229] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_230 bl[230] br[230] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_231 bl[231] br[231] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_232 bl[232] br[232] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_233 bl[233] br[233] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_234 bl[234] br[234] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_235 bl[235] br[235] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_236 bl[236] br[236] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_237 bl[237] br[237] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_238 bl[238] br[238] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_239 bl[239] br[239] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_240 bl[240] br[240] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_241 bl[241] br[241] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_242 bl[242] br[242] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_243 bl[243] br[243] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_244 bl[244] br[244] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_245 bl[245] br[245] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_246 bl[246] br[246] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_247 bl[247] br[247] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_248 bl[248] br[248] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_249 bl[249] br[249] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_250 bl[250] br[250] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_251 bl[251] br[251] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_252 bl[252] br[252] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_253 bl[253] br[253] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_254 bl[254] br[254] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_255 bl[255] br[255] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_33_0 bl[0] br[0] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_1 bl[1] br[1] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_2 bl[2] br[2] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_3 bl[3] br[3] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_4 bl[4] br[4] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_5 bl[5] br[5] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_6 bl[6] br[6] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_7 bl[7] br[7] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_8 bl[8] br[8] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_9 bl[9] br[9] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_10 bl[10] br[10] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_11 bl[11] br[11] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_12 bl[12] br[12] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_13 bl[13] br[13] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_14 bl[14] br[14] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_15 bl[15] br[15] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_16 bl[16] br[16] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_17 bl[17] br[17] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_18 bl[18] br[18] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_19 bl[19] br[19] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_20 bl[20] br[20] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_21 bl[21] br[21] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_22 bl[22] br[22] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_23 bl[23] br[23] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_24 bl[24] br[24] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_25 bl[25] br[25] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_26 bl[26] br[26] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_27 bl[27] br[27] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_28 bl[28] br[28] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_29 bl[29] br[29] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_30 bl[30] br[30] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_31 bl[31] br[31] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_32 bl[32] br[32] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_33 bl[33] br[33] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_34 bl[34] br[34] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_35 bl[35] br[35] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_36 bl[36] br[36] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_37 bl[37] br[37] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_38 bl[38] br[38] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_39 bl[39] br[39] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_40 bl[40] br[40] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_41 bl[41] br[41] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_42 bl[42] br[42] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_43 bl[43] br[43] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_44 bl[44] br[44] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_45 bl[45] br[45] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_46 bl[46] br[46] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_47 bl[47] br[47] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_48 bl[48] br[48] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_49 bl[49] br[49] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_50 bl[50] br[50] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_51 bl[51] br[51] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_52 bl[52] br[52] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_53 bl[53] br[53] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_54 bl[54] br[54] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_55 bl[55] br[55] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_56 bl[56] br[56] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_57 bl[57] br[57] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_58 bl[58] br[58] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_59 bl[59] br[59] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_60 bl[60] br[60] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_61 bl[61] br[61] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_62 bl[62] br[62] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_63 bl[63] br[63] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_64 bl[64] br[64] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_65 bl[65] br[65] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_66 bl[66] br[66] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_67 bl[67] br[67] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_68 bl[68] br[68] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_69 bl[69] br[69] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_70 bl[70] br[70] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_71 bl[71] br[71] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_72 bl[72] br[72] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_73 bl[73] br[73] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_74 bl[74] br[74] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_75 bl[75] br[75] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_76 bl[76] br[76] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_77 bl[77] br[77] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_78 bl[78] br[78] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_79 bl[79] br[79] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_80 bl[80] br[80] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_81 bl[81] br[81] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_82 bl[82] br[82] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_83 bl[83] br[83] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_84 bl[84] br[84] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_85 bl[85] br[85] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_86 bl[86] br[86] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_87 bl[87] br[87] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_88 bl[88] br[88] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_89 bl[89] br[89] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_90 bl[90] br[90] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_91 bl[91] br[91] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_92 bl[92] br[92] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_93 bl[93] br[93] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_94 bl[94] br[94] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_95 bl[95] br[95] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_96 bl[96] br[96] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_97 bl[97] br[97] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_98 bl[98] br[98] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_99 bl[99] br[99] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_100 bl[100] br[100] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_101 bl[101] br[101] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_102 bl[102] br[102] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_103 bl[103] br[103] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_104 bl[104] br[104] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_105 bl[105] br[105] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_106 bl[106] br[106] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_107 bl[107] br[107] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_108 bl[108] br[108] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_109 bl[109] br[109] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_110 bl[110] br[110] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_111 bl[111] br[111] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_112 bl[112] br[112] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_113 bl[113] br[113] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_114 bl[114] br[114] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_115 bl[115] br[115] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_116 bl[116] br[116] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_117 bl[117] br[117] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_118 bl[118] br[118] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_119 bl[119] br[119] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_120 bl[120] br[120] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_121 bl[121] br[121] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_122 bl[122] br[122] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_123 bl[123] br[123] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_124 bl[124] br[124] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_125 bl[125] br[125] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_126 bl[126] br[126] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_127 bl[127] br[127] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_128 bl[128] br[128] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_129 bl[129] br[129] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_130 bl[130] br[130] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_131 bl[131] br[131] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_132 bl[132] br[132] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_133 bl[133] br[133] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_134 bl[134] br[134] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_135 bl[135] br[135] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_136 bl[136] br[136] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_137 bl[137] br[137] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_138 bl[138] br[138] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_139 bl[139] br[139] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_140 bl[140] br[140] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_141 bl[141] br[141] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_142 bl[142] br[142] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_143 bl[143] br[143] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_144 bl[144] br[144] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_145 bl[145] br[145] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_146 bl[146] br[146] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_147 bl[147] br[147] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_148 bl[148] br[148] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_149 bl[149] br[149] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_150 bl[150] br[150] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_151 bl[151] br[151] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_152 bl[152] br[152] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_153 bl[153] br[153] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_154 bl[154] br[154] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_155 bl[155] br[155] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_156 bl[156] br[156] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_157 bl[157] br[157] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_158 bl[158] br[158] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_159 bl[159] br[159] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_160 bl[160] br[160] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_161 bl[161] br[161] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_162 bl[162] br[162] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_163 bl[163] br[163] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_164 bl[164] br[164] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_165 bl[165] br[165] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_166 bl[166] br[166] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_167 bl[167] br[167] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_168 bl[168] br[168] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_169 bl[169] br[169] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_170 bl[170] br[170] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_171 bl[171] br[171] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_172 bl[172] br[172] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_173 bl[173] br[173] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_174 bl[174] br[174] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_175 bl[175] br[175] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_176 bl[176] br[176] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_177 bl[177] br[177] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_178 bl[178] br[178] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_179 bl[179] br[179] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_180 bl[180] br[180] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_181 bl[181] br[181] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_182 bl[182] br[182] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_183 bl[183] br[183] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_184 bl[184] br[184] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_185 bl[185] br[185] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_186 bl[186] br[186] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_187 bl[187] br[187] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_188 bl[188] br[188] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_189 bl[189] br[189] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_190 bl[190] br[190] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_191 bl[191] br[191] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_192 bl[192] br[192] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_193 bl[193] br[193] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_194 bl[194] br[194] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_195 bl[195] br[195] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_196 bl[196] br[196] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_197 bl[197] br[197] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_198 bl[198] br[198] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_199 bl[199] br[199] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_200 bl[200] br[200] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_201 bl[201] br[201] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_202 bl[202] br[202] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_203 bl[203] br[203] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_204 bl[204] br[204] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_205 bl[205] br[205] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_206 bl[206] br[206] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_207 bl[207] br[207] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_208 bl[208] br[208] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_209 bl[209] br[209] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_210 bl[210] br[210] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_211 bl[211] br[211] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_212 bl[212] br[212] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_213 bl[213] br[213] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_214 bl[214] br[214] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_215 bl[215] br[215] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_216 bl[216] br[216] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_217 bl[217] br[217] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_218 bl[218] br[218] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_219 bl[219] br[219] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_220 bl[220] br[220] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_221 bl[221] br[221] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_222 bl[222] br[222] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_223 bl[223] br[223] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_224 bl[224] br[224] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_225 bl[225] br[225] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_226 bl[226] br[226] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_227 bl[227] br[227] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_228 bl[228] br[228] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_229 bl[229] br[229] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_230 bl[230] br[230] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_231 bl[231] br[231] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_232 bl[232] br[232] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_233 bl[233] br[233] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_234 bl[234] br[234] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_235 bl[235] br[235] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_236 bl[236] br[236] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_237 bl[237] br[237] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_238 bl[238] br[238] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_239 bl[239] br[239] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_240 bl[240] br[240] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_241 bl[241] br[241] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_242 bl[242] br[242] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_243 bl[243] br[243] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_244 bl[244] br[244] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_245 bl[245] br[245] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_246 bl[246] br[246] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_247 bl[247] br[247] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_248 bl[248] br[248] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_249 bl[249] br[249] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_250 bl[250] br[250] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_251 bl[251] br[251] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_252 bl[252] br[252] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_253 bl[253] br[253] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_254 bl[254] br[254] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_255 bl[255] br[255] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_34_0 bl[0] br[0] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_1 bl[1] br[1] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_2 bl[2] br[2] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_3 bl[3] br[3] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_4 bl[4] br[4] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_5 bl[5] br[5] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_6 bl[6] br[6] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_7 bl[7] br[7] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_8 bl[8] br[8] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_9 bl[9] br[9] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_10 bl[10] br[10] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_11 bl[11] br[11] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_12 bl[12] br[12] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_13 bl[13] br[13] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_14 bl[14] br[14] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_15 bl[15] br[15] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_16 bl[16] br[16] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_17 bl[17] br[17] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_18 bl[18] br[18] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_19 bl[19] br[19] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_20 bl[20] br[20] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_21 bl[21] br[21] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_22 bl[22] br[22] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_23 bl[23] br[23] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_24 bl[24] br[24] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_25 bl[25] br[25] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_26 bl[26] br[26] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_27 bl[27] br[27] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_28 bl[28] br[28] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_29 bl[29] br[29] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_30 bl[30] br[30] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_31 bl[31] br[31] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_32 bl[32] br[32] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_33 bl[33] br[33] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_34 bl[34] br[34] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_35 bl[35] br[35] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_36 bl[36] br[36] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_37 bl[37] br[37] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_38 bl[38] br[38] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_39 bl[39] br[39] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_40 bl[40] br[40] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_41 bl[41] br[41] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_42 bl[42] br[42] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_43 bl[43] br[43] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_44 bl[44] br[44] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_45 bl[45] br[45] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_46 bl[46] br[46] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_47 bl[47] br[47] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_48 bl[48] br[48] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_49 bl[49] br[49] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_50 bl[50] br[50] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_51 bl[51] br[51] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_52 bl[52] br[52] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_53 bl[53] br[53] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_54 bl[54] br[54] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_55 bl[55] br[55] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_56 bl[56] br[56] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_57 bl[57] br[57] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_58 bl[58] br[58] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_59 bl[59] br[59] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_60 bl[60] br[60] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_61 bl[61] br[61] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_62 bl[62] br[62] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_63 bl[63] br[63] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_64 bl[64] br[64] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_65 bl[65] br[65] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_66 bl[66] br[66] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_67 bl[67] br[67] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_68 bl[68] br[68] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_69 bl[69] br[69] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_70 bl[70] br[70] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_71 bl[71] br[71] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_72 bl[72] br[72] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_73 bl[73] br[73] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_74 bl[74] br[74] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_75 bl[75] br[75] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_76 bl[76] br[76] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_77 bl[77] br[77] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_78 bl[78] br[78] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_79 bl[79] br[79] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_80 bl[80] br[80] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_81 bl[81] br[81] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_82 bl[82] br[82] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_83 bl[83] br[83] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_84 bl[84] br[84] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_85 bl[85] br[85] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_86 bl[86] br[86] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_87 bl[87] br[87] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_88 bl[88] br[88] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_89 bl[89] br[89] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_90 bl[90] br[90] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_91 bl[91] br[91] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_92 bl[92] br[92] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_93 bl[93] br[93] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_94 bl[94] br[94] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_95 bl[95] br[95] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_96 bl[96] br[96] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_97 bl[97] br[97] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_98 bl[98] br[98] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_99 bl[99] br[99] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_100 bl[100] br[100] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_101 bl[101] br[101] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_102 bl[102] br[102] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_103 bl[103] br[103] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_104 bl[104] br[104] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_105 bl[105] br[105] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_106 bl[106] br[106] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_107 bl[107] br[107] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_108 bl[108] br[108] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_109 bl[109] br[109] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_110 bl[110] br[110] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_111 bl[111] br[111] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_112 bl[112] br[112] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_113 bl[113] br[113] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_114 bl[114] br[114] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_115 bl[115] br[115] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_116 bl[116] br[116] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_117 bl[117] br[117] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_118 bl[118] br[118] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_119 bl[119] br[119] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_120 bl[120] br[120] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_121 bl[121] br[121] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_122 bl[122] br[122] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_123 bl[123] br[123] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_124 bl[124] br[124] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_125 bl[125] br[125] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_126 bl[126] br[126] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_127 bl[127] br[127] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_128 bl[128] br[128] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_129 bl[129] br[129] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_130 bl[130] br[130] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_131 bl[131] br[131] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_132 bl[132] br[132] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_133 bl[133] br[133] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_134 bl[134] br[134] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_135 bl[135] br[135] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_136 bl[136] br[136] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_137 bl[137] br[137] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_138 bl[138] br[138] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_139 bl[139] br[139] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_140 bl[140] br[140] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_141 bl[141] br[141] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_142 bl[142] br[142] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_143 bl[143] br[143] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_144 bl[144] br[144] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_145 bl[145] br[145] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_146 bl[146] br[146] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_147 bl[147] br[147] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_148 bl[148] br[148] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_149 bl[149] br[149] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_150 bl[150] br[150] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_151 bl[151] br[151] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_152 bl[152] br[152] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_153 bl[153] br[153] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_154 bl[154] br[154] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_155 bl[155] br[155] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_156 bl[156] br[156] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_157 bl[157] br[157] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_158 bl[158] br[158] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_159 bl[159] br[159] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_160 bl[160] br[160] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_161 bl[161] br[161] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_162 bl[162] br[162] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_163 bl[163] br[163] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_164 bl[164] br[164] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_165 bl[165] br[165] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_166 bl[166] br[166] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_167 bl[167] br[167] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_168 bl[168] br[168] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_169 bl[169] br[169] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_170 bl[170] br[170] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_171 bl[171] br[171] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_172 bl[172] br[172] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_173 bl[173] br[173] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_174 bl[174] br[174] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_175 bl[175] br[175] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_176 bl[176] br[176] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_177 bl[177] br[177] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_178 bl[178] br[178] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_179 bl[179] br[179] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_180 bl[180] br[180] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_181 bl[181] br[181] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_182 bl[182] br[182] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_183 bl[183] br[183] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_184 bl[184] br[184] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_185 bl[185] br[185] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_186 bl[186] br[186] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_187 bl[187] br[187] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_188 bl[188] br[188] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_189 bl[189] br[189] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_190 bl[190] br[190] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_191 bl[191] br[191] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_192 bl[192] br[192] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_193 bl[193] br[193] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_194 bl[194] br[194] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_195 bl[195] br[195] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_196 bl[196] br[196] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_197 bl[197] br[197] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_198 bl[198] br[198] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_199 bl[199] br[199] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_200 bl[200] br[200] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_201 bl[201] br[201] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_202 bl[202] br[202] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_203 bl[203] br[203] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_204 bl[204] br[204] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_205 bl[205] br[205] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_206 bl[206] br[206] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_207 bl[207] br[207] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_208 bl[208] br[208] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_209 bl[209] br[209] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_210 bl[210] br[210] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_211 bl[211] br[211] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_212 bl[212] br[212] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_213 bl[213] br[213] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_214 bl[214] br[214] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_215 bl[215] br[215] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_216 bl[216] br[216] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_217 bl[217] br[217] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_218 bl[218] br[218] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_219 bl[219] br[219] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_220 bl[220] br[220] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_221 bl[221] br[221] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_222 bl[222] br[222] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_223 bl[223] br[223] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_224 bl[224] br[224] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_225 bl[225] br[225] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_226 bl[226] br[226] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_227 bl[227] br[227] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_228 bl[228] br[228] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_229 bl[229] br[229] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_230 bl[230] br[230] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_231 bl[231] br[231] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_232 bl[232] br[232] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_233 bl[233] br[233] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_234 bl[234] br[234] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_235 bl[235] br[235] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_236 bl[236] br[236] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_237 bl[237] br[237] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_238 bl[238] br[238] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_239 bl[239] br[239] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_240 bl[240] br[240] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_241 bl[241] br[241] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_242 bl[242] br[242] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_243 bl[243] br[243] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_244 bl[244] br[244] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_245 bl[245] br[245] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_246 bl[246] br[246] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_247 bl[247] br[247] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_248 bl[248] br[248] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_249 bl[249] br[249] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_250 bl[250] br[250] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_251 bl[251] br[251] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_252 bl[252] br[252] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_253 bl[253] br[253] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_254 bl[254] br[254] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_255 bl[255] br[255] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_35_0 bl[0] br[0] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_1 bl[1] br[1] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_2 bl[2] br[2] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_3 bl[3] br[3] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_4 bl[4] br[4] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_5 bl[5] br[5] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_6 bl[6] br[6] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_7 bl[7] br[7] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_8 bl[8] br[8] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_9 bl[9] br[9] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_10 bl[10] br[10] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_11 bl[11] br[11] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_12 bl[12] br[12] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_13 bl[13] br[13] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_14 bl[14] br[14] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_15 bl[15] br[15] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_16 bl[16] br[16] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_17 bl[17] br[17] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_18 bl[18] br[18] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_19 bl[19] br[19] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_20 bl[20] br[20] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_21 bl[21] br[21] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_22 bl[22] br[22] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_23 bl[23] br[23] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_24 bl[24] br[24] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_25 bl[25] br[25] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_26 bl[26] br[26] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_27 bl[27] br[27] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_28 bl[28] br[28] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_29 bl[29] br[29] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_30 bl[30] br[30] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_31 bl[31] br[31] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_32 bl[32] br[32] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_33 bl[33] br[33] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_34 bl[34] br[34] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_35 bl[35] br[35] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_36 bl[36] br[36] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_37 bl[37] br[37] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_38 bl[38] br[38] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_39 bl[39] br[39] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_40 bl[40] br[40] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_41 bl[41] br[41] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_42 bl[42] br[42] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_43 bl[43] br[43] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_44 bl[44] br[44] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_45 bl[45] br[45] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_46 bl[46] br[46] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_47 bl[47] br[47] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_48 bl[48] br[48] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_49 bl[49] br[49] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_50 bl[50] br[50] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_51 bl[51] br[51] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_52 bl[52] br[52] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_53 bl[53] br[53] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_54 bl[54] br[54] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_55 bl[55] br[55] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_56 bl[56] br[56] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_57 bl[57] br[57] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_58 bl[58] br[58] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_59 bl[59] br[59] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_60 bl[60] br[60] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_61 bl[61] br[61] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_62 bl[62] br[62] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_63 bl[63] br[63] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_64 bl[64] br[64] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_65 bl[65] br[65] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_66 bl[66] br[66] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_67 bl[67] br[67] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_68 bl[68] br[68] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_69 bl[69] br[69] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_70 bl[70] br[70] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_71 bl[71] br[71] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_72 bl[72] br[72] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_73 bl[73] br[73] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_74 bl[74] br[74] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_75 bl[75] br[75] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_76 bl[76] br[76] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_77 bl[77] br[77] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_78 bl[78] br[78] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_79 bl[79] br[79] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_80 bl[80] br[80] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_81 bl[81] br[81] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_82 bl[82] br[82] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_83 bl[83] br[83] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_84 bl[84] br[84] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_85 bl[85] br[85] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_86 bl[86] br[86] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_87 bl[87] br[87] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_88 bl[88] br[88] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_89 bl[89] br[89] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_90 bl[90] br[90] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_91 bl[91] br[91] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_92 bl[92] br[92] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_93 bl[93] br[93] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_94 bl[94] br[94] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_95 bl[95] br[95] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_96 bl[96] br[96] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_97 bl[97] br[97] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_98 bl[98] br[98] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_99 bl[99] br[99] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_100 bl[100] br[100] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_101 bl[101] br[101] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_102 bl[102] br[102] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_103 bl[103] br[103] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_104 bl[104] br[104] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_105 bl[105] br[105] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_106 bl[106] br[106] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_107 bl[107] br[107] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_108 bl[108] br[108] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_109 bl[109] br[109] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_110 bl[110] br[110] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_111 bl[111] br[111] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_112 bl[112] br[112] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_113 bl[113] br[113] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_114 bl[114] br[114] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_115 bl[115] br[115] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_116 bl[116] br[116] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_117 bl[117] br[117] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_118 bl[118] br[118] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_119 bl[119] br[119] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_120 bl[120] br[120] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_121 bl[121] br[121] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_122 bl[122] br[122] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_123 bl[123] br[123] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_124 bl[124] br[124] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_125 bl[125] br[125] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_126 bl[126] br[126] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_127 bl[127] br[127] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_128 bl[128] br[128] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_129 bl[129] br[129] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_130 bl[130] br[130] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_131 bl[131] br[131] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_132 bl[132] br[132] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_133 bl[133] br[133] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_134 bl[134] br[134] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_135 bl[135] br[135] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_136 bl[136] br[136] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_137 bl[137] br[137] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_138 bl[138] br[138] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_139 bl[139] br[139] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_140 bl[140] br[140] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_141 bl[141] br[141] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_142 bl[142] br[142] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_143 bl[143] br[143] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_144 bl[144] br[144] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_145 bl[145] br[145] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_146 bl[146] br[146] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_147 bl[147] br[147] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_148 bl[148] br[148] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_149 bl[149] br[149] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_150 bl[150] br[150] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_151 bl[151] br[151] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_152 bl[152] br[152] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_153 bl[153] br[153] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_154 bl[154] br[154] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_155 bl[155] br[155] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_156 bl[156] br[156] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_157 bl[157] br[157] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_158 bl[158] br[158] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_159 bl[159] br[159] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_160 bl[160] br[160] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_161 bl[161] br[161] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_162 bl[162] br[162] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_163 bl[163] br[163] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_164 bl[164] br[164] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_165 bl[165] br[165] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_166 bl[166] br[166] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_167 bl[167] br[167] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_168 bl[168] br[168] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_169 bl[169] br[169] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_170 bl[170] br[170] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_171 bl[171] br[171] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_172 bl[172] br[172] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_173 bl[173] br[173] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_174 bl[174] br[174] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_175 bl[175] br[175] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_176 bl[176] br[176] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_177 bl[177] br[177] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_178 bl[178] br[178] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_179 bl[179] br[179] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_180 bl[180] br[180] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_181 bl[181] br[181] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_182 bl[182] br[182] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_183 bl[183] br[183] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_184 bl[184] br[184] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_185 bl[185] br[185] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_186 bl[186] br[186] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_187 bl[187] br[187] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_188 bl[188] br[188] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_189 bl[189] br[189] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_190 bl[190] br[190] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_191 bl[191] br[191] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_192 bl[192] br[192] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_193 bl[193] br[193] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_194 bl[194] br[194] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_195 bl[195] br[195] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_196 bl[196] br[196] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_197 bl[197] br[197] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_198 bl[198] br[198] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_199 bl[199] br[199] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_200 bl[200] br[200] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_201 bl[201] br[201] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_202 bl[202] br[202] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_203 bl[203] br[203] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_204 bl[204] br[204] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_205 bl[205] br[205] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_206 bl[206] br[206] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_207 bl[207] br[207] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_208 bl[208] br[208] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_209 bl[209] br[209] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_210 bl[210] br[210] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_211 bl[211] br[211] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_212 bl[212] br[212] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_213 bl[213] br[213] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_214 bl[214] br[214] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_215 bl[215] br[215] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_216 bl[216] br[216] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_217 bl[217] br[217] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_218 bl[218] br[218] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_219 bl[219] br[219] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_220 bl[220] br[220] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_221 bl[221] br[221] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_222 bl[222] br[222] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_223 bl[223] br[223] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_224 bl[224] br[224] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_225 bl[225] br[225] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_226 bl[226] br[226] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_227 bl[227] br[227] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_228 bl[228] br[228] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_229 bl[229] br[229] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_230 bl[230] br[230] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_231 bl[231] br[231] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_232 bl[232] br[232] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_233 bl[233] br[233] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_234 bl[234] br[234] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_235 bl[235] br[235] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_236 bl[236] br[236] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_237 bl[237] br[237] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_238 bl[238] br[238] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_239 bl[239] br[239] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_240 bl[240] br[240] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_241 bl[241] br[241] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_242 bl[242] br[242] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_243 bl[243] br[243] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_244 bl[244] br[244] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_245 bl[245] br[245] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_246 bl[246] br[246] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_247 bl[247] br[247] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_248 bl[248] br[248] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_249 bl[249] br[249] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_250 bl[250] br[250] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_251 bl[251] br[251] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_252 bl[252] br[252] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_253 bl[253] br[253] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_254 bl[254] br[254] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_255 bl[255] br[255] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_36_0 bl[0] br[0] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_1 bl[1] br[1] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_2 bl[2] br[2] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_3 bl[3] br[3] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_4 bl[4] br[4] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_5 bl[5] br[5] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_6 bl[6] br[6] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_7 bl[7] br[7] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_8 bl[8] br[8] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_9 bl[9] br[9] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_10 bl[10] br[10] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_11 bl[11] br[11] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_12 bl[12] br[12] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_13 bl[13] br[13] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_14 bl[14] br[14] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_15 bl[15] br[15] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_16 bl[16] br[16] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_17 bl[17] br[17] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_18 bl[18] br[18] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_19 bl[19] br[19] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_20 bl[20] br[20] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_21 bl[21] br[21] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_22 bl[22] br[22] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_23 bl[23] br[23] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_24 bl[24] br[24] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_25 bl[25] br[25] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_26 bl[26] br[26] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_27 bl[27] br[27] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_28 bl[28] br[28] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_29 bl[29] br[29] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_30 bl[30] br[30] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_31 bl[31] br[31] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_32 bl[32] br[32] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_33 bl[33] br[33] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_34 bl[34] br[34] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_35 bl[35] br[35] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_36 bl[36] br[36] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_37 bl[37] br[37] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_38 bl[38] br[38] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_39 bl[39] br[39] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_40 bl[40] br[40] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_41 bl[41] br[41] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_42 bl[42] br[42] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_43 bl[43] br[43] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_44 bl[44] br[44] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_45 bl[45] br[45] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_46 bl[46] br[46] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_47 bl[47] br[47] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_48 bl[48] br[48] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_49 bl[49] br[49] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_50 bl[50] br[50] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_51 bl[51] br[51] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_52 bl[52] br[52] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_53 bl[53] br[53] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_54 bl[54] br[54] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_55 bl[55] br[55] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_56 bl[56] br[56] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_57 bl[57] br[57] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_58 bl[58] br[58] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_59 bl[59] br[59] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_60 bl[60] br[60] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_61 bl[61] br[61] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_62 bl[62] br[62] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_63 bl[63] br[63] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_64 bl[64] br[64] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_65 bl[65] br[65] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_66 bl[66] br[66] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_67 bl[67] br[67] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_68 bl[68] br[68] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_69 bl[69] br[69] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_70 bl[70] br[70] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_71 bl[71] br[71] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_72 bl[72] br[72] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_73 bl[73] br[73] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_74 bl[74] br[74] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_75 bl[75] br[75] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_76 bl[76] br[76] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_77 bl[77] br[77] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_78 bl[78] br[78] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_79 bl[79] br[79] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_80 bl[80] br[80] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_81 bl[81] br[81] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_82 bl[82] br[82] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_83 bl[83] br[83] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_84 bl[84] br[84] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_85 bl[85] br[85] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_86 bl[86] br[86] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_87 bl[87] br[87] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_88 bl[88] br[88] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_89 bl[89] br[89] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_90 bl[90] br[90] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_91 bl[91] br[91] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_92 bl[92] br[92] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_93 bl[93] br[93] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_94 bl[94] br[94] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_95 bl[95] br[95] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_96 bl[96] br[96] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_97 bl[97] br[97] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_98 bl[98] br[98] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_99 bl[99] br[99] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_100 bl[100] br[100] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_101 bl[101] br[101] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_102 bl[102] br[102] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_103 bl[103] br[103] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_104 bl[104] br[104] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_105 bl[105] br[105] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_106 bl[106] br[106] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_107 bl[107] br[107] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_108 bl[108] br[108] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_109 bl[109] br[109] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_110 bl[110] br[110] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_111 bl[111] br[111] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_112 bl[112] br[112] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_113 bl[113] br[113] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_114 bl[114] br[114] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_115 bl[115] br[115] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_116 bl[116] br[116] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_117 bl[117] br[117] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_118 bl[118] br[118] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_119 bl[119] br[119] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_120 bl[120] br[120] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_121 bl[121] br[121] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_122 bl[122] br[122] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_123 bl[123] br[123] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_124 bl[124] br[124] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_125 bl[125] br[125] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_126 bl[126] br[126] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_127 bl[127] br[127] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_128 bl[128] br[128] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_129 bl[129] br[129] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_130 bl[130] br[130] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_131 bl[131] br[131] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_132 bl[132] br[132] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_133 bl[133] br[133] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_134 bl[134] br[134] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_135 bl[135] br[135] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_136 bl[136] br[136] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_137 bl[137] br[137] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_138 bl[138] br[138] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_139 bl[139] br[139] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_140 bl[140] br[140] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_141 bl[141] br[141] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_142 bl[142] br[142] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_143 bl[143] br[143] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_144 bl[144] br[144] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_145 bl[145] br[145] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_146 bl[146] br[146] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_147 bl[147] br[147] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_148 bl[148] br[148] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_149 bl[149] br[149] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_150 bl[150] br[150] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_151 bl[151] br[151] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_152 bl[152] br[152] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_153 bl[153] br[153] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_154 bl[154] br[154] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_155 bl[155] br[155] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_156 bl[156] br[156] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_157 bl[157] br[157] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_158 bl[158] br[158] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_159 bl[159] br[159] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_160 bl[160] br[160] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_161 bl[161] br[161] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_162 bl[162] br[162] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_163 bl[163] br[163] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_164 bl[164] br[164] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_165 bl[165] br[165] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_166 bl[166] br[166] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_167 bl[167] br[167] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_168 bl[168] br[168] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_169 bl[169] br[169] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_170 bl[170] br[170] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_171 bl[171] br[171] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_172 bl[172] br[172] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_173 bl[173] br[173] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_174 bl[174] br[174] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_175 bl[175] br[175] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_176 bl[176] br[176] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_177 bl[177] br[177] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_178 bl[178] br[178] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_179 bl[179] br[179] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_180 bl[180] br[180] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_181 bl[181] br[181] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_182 bl[182] br[182] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_183 bl[183] br[183] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_184 bl[184] br[184] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_185 bl[185] br[185] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_186 bl[186] br[186] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_187 bl[187] br[187] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_188 bl[188] br[188] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_189 bl[189] br[189] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_190 bl[190] br[190] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_191 bl[191] br[191] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_192 bl[192] br[192] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_193 bl[193] br[193] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_194 bl[194] br[194] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_195 bl[195] br[195] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_196 bl[196] br[196] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_197 bl[197] br[197] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_198 bl[198] br[198] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_199 bl[199] br[199] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_200 bl[200] br[200] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_201 bl[201] br[201] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_202 bl[202] br[202] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_203 bl[203] br[203] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_204 bl[204] br[204] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_205 bl[205] br[205] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_206 bl[206] br[206] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_207 bl[207] br[207] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_208 bl[208] br[208] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_209 bl[209] br[209] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_210 bl[210] br[210] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_211 bl[211] br[211] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_212 bl[212] br[212] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_213 bl[213] br[213] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_214 bl[214] br[214] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_215 bl[215] br[215] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_216 bl[216] br[216] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_217 bl[217] br[217] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_218 bl[218] br[218] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_219 bl[219] br[219] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_220 bl[220] br[220] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_221 bl[221] br[221] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_222 bl[222] br[222] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_223 bl[223] br[223] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_224 bl[224] br[224] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_225 bl[225] br[225] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_226 bl[226] br[226] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_227 bl[227] br[227] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_228 bl[228] br[228] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_229 bl[229] br[229] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_230 bl[230] br[230] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_231 bl[231] br[231] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_232 bl[232] br[232] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_233 bl[233] br[233] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_234 bl[234] br[234] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_235 bl[235] br[235] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_236 bl[236] br[236] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_237 bl[237] br[237] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_238 bl[238] br[238] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_239 bl[239] br[239] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_240 bl[240] br[240] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_241 bl[241] br[241] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_242 bl[242] br[242] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_243 bl[243] br[243] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_244 bl[244] br[244] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_245 bl[245] br[245] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_246 bl[246] br[246] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_247 bl[247] br[247] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_248 bl[248] br[248] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_249 bl[249] br[249] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_250 bl[250] br[250] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_251 bl[251] br[251] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_252 bl[252] br[252] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_253 bl[253] br[253] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_254 bl[254] br[254] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_255 bl[255] br[255] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_37_0 bl[0] br[0] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_1 bl[1] br[1] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_2 bl[2] br[2] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_3 bl[3] br[3] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_4 bl[4] br[4] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_5 bl[5] br[5] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_6 bl[6] br[6] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_7 bl[7] br[7] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_8 bl[8] br[8] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_9 bl[9] br[9] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_10 bl[10] br[10] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_11 bl[11] br[11] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_12 bl[12] br[12] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_13 bl[13] br[13] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_14 bl[14] br[14] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_15 bl[15] br[15] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_16 bl[16] br[16] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_17 bl[17] br[17] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_18 bl[18] br[18] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_19 bl[19] br[19] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_20 bl[20] br[20] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_21 bl[21] br[21] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_22 bl[22] br[22] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_23 bl[23] br[23] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_24 bl[24] br[24] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_25 bl[25] br[25] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_26 bl[26] br[26] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_27 bl[27] br[27] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_28 bl[28] br[28] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_29 bl[29] br[29] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_30 bl[30] br[30] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_31 bl[31] br[31] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_32 bl[32] br[32] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_33 bl[33] br[33] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_34 bl[34] br[34] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_35 bl[35] br[35] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_36 bl[36] br[36] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_37 bl[37] br[37] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_38 bl[38] br[38] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_39 bl[39] br[39] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_40 bl[40] br[40] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_41 bl[41] br[41] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_42 bl[42] br[42] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_43 bl[43] br[43] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_44 bl[44] br[44] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_45 bl[45] br[45] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_46 bl[46] br[46] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_47 bl[47] br[47] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_48 bl[48] br[48] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_49 bl[49] br[49] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_50 bl[50] br[50] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_51 bl[51] br[51] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_52 bl[52] br[52] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_53 bl[53] br[53] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_54 bl[54] br[54] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_55 bl[55] br[55] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_56 bl[56] br[56] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_57 bl[57] br[57] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_58 bl[58] br[58] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_59 bl[59] br[59] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_60 bl[60] br[60] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_61 bl[61] br[61] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_62 bl[62] br[62] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_63 bl[63] br[63] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_64 bl[64] br[64] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_65 bl[65] br[65] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_66 bl[66] br[66] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_67 bl[67] br[67] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_68 bl[68] br[68] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_69 bl[69] br[69] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_70 bl[70] br[70] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_71 bl[71] br[71] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_72 bl[72] br[72] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_73 bl[73] br[73] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_74 bl[74] br[74] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_75 bl[75] br[75] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_76 bl[76] br[76] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_77 bl[77] br[77] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_78 bl[78] br[78] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_79 bl[79] br[79] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_80 bl[80] br[80] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_81 bl[81] br[81] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_82 bl[82] br[82] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_83 bl[83] br[83] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_84 bl[84] br[84] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_85 bl[85] br[85] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_86 bl[86] br[86] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_87 bl[87] br[87] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_88 bl[88] br[88] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_89 bl[89] br[89] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_90 bl[90] br[90] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_91 bl[91] br[91] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_92 bl[92] br[92] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_93 bl[93] br[93] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_94 bl[94] br[94] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_95 bl[95] br[95] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_96 bl[96] br[96] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_97 bl[97] br[97] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_98 bl[98] br[98] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_99 bl[99] br[99] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_100 bl[100] br[100] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_101 bl[101] br[101] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_102 bl[102] br[102] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_103 bl[103] br[103] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_104 bl[104] br[104] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_105 bl[105] br[105] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_106 bl[106] br[106] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_107 bl[107] br[107] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_108 bl[108] br[108] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_109 bl[109] br[109] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_110 bl[110] br[110] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_111 bl[111] br[111] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_112 bl[112] br[112] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_113 bl[113] br[113] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_114 bl[114] br[114] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_115 bl[115] br[115] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_116 bl[116] br[116] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_117 bl[117] br[117] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_118 bl[118] br[118] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_119 bl[119] br[119] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_120 bl[120] br[120] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_121 bl[121] br[121] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_122 bl[122] br[122] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_123 bl[123] br[123] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_124 bl[124] br[124] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_125 bl[125] br[125] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_126 bl[126] br[126] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_127 bl[127] br[127] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_128 bl[128] br[128] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_129 bl[129] br[129] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_130 bl[130] br[130] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_131 bl[131] br[131] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_132 bl[132] br[132] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_133 bl[133] br[133] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_134 bl[134] br[134] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_135 bl[135] br[135] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_136 bl[136] br[136] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_137 bl[137] br[137] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_138 bl[138] br[138] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_139 bl[139] br[139] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_140 bl[140] br[140] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_141 bl[141] br[141] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_142 bl[142] br[142] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_143 bl[143] br[143] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_144 bl[144] br[144] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_145 bl[145] br[145] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_146 bl[146] br[146] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_147 bl[147] br[147] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_148 bl[148] br[148] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_149 bl[149] br[149] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_150 bl[150] br[150] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_151 bl[151] br[151] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_152 bl[152] br[152] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_153 bl[153] br[153] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_154 bl[154] br[154] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_155 bl[155] br[155] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_156 bl[156] br[156] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_157 bl[157] br[157] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_158 bl[158] br[158] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_159 bl[159] br[159] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_160 bl[160] br[160] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_161 bl[161] br[161] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_162 bl[162] br[162] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_163 bl[163] br[163] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_164 bl[164] br[164] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_165 bl[165] br[165] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_166 bl[166] br[166] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_167 bl[167] br[167] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_168 bl[168] br[168] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_169 bl[169] br[169] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_170 bl[170] br[170] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_171 bl[171] br[171] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_172 bl[172] br[172] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_173 bl[173] br[173] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_174 bl[174] br[174] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_175 bl[175] br[175] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_176 bl[176] br[176] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_177 bl[177] br[177] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_178 bl[178] br[178] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_179 bl[179] br[179] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_180 bl[180] br[180] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_181 bl[181] br[181] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_182 bl[182] br[182] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_183 bl[183] br[183] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_184 bl[184] br[184] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_185 bl[185] br[185] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_186 bl[186] br[186] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_187 bl[187] br[187] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_188 bl[188] br[188] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_189 bl[189] br[189] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_190 bl[190] br[190] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_191 bl[191] br[191] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_192 bl[192] br[192] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_193 bl[193] br[193] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_194 bl[194] br[194] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_195 bl[195] br[195] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_196 bl[196] br[196] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_197 bl[197] br[197] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_198 bl[198] br[198] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_199 bl[199] br[199] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_200 bl[200] br[200] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_201 bl[201] br[201] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_202 bl[202] br[202] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_203 bl[203] br[203] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_204 bl[204] br[204] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_205 bl[205] br[205] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_206 bl[206] br[206] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_207 bl[207] br[207] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_208 bl[208] br[208] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_209 bl[209] br[209] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_210 bl[210] br[210] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_211 bl[211] br[211] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_212 bl[212] br[212] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_213 bl[213] br[213] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_214 bl[214] br[214] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_215 bl[215] br[215] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_216 bl[216] br[216] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_217 bl[217] br[217] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_218 bl[218] br[218] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_219 bl[219] br[219] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_220 bl[220] br[220] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_221 bl[221] br[221] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_222 bl[222] br[222] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_223 bl[223] br[223] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_224 bl[224] br[224] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_225 bl[225] br[225] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_226 bl[226] br[226] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_227 bl[227] br[227] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_228 bl[228] br[228] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_229 bl[229] br[229] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_230 bl[230] br[230] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_231 bl[231] br[231] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_232 bl[232] br[232] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_233 bl[233] br[233] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_234 bl[234] br[234] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_235 bl[235] br[235] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_236 bl[236] br[236] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_237 bl[237] br[237] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_238 bl[238] br[238] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_239 bl[239] br[239] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_240 bl[240] br[240] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_241 bl[241] br[241] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_242 bl[242] br[242] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_243 bl[243] br[243] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_244 bl[244] br[244] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_245 bl[245] br[245] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_246 bl[246] br[246] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_247 bl[247] br[247] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_248 bl[248] br[248] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_249 bl[249] br[249] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_250 bl[250] br[250] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_251 bl[251] br[251] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_252 bl[252] br[252] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_253 bl[253] br[253] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_254 bl[254] br[254] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_255 bl[255] br[255] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_38_0 bl[0] br[0] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_1 bl[1] br[1] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_2 bl[2] br[2] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_3 bl[3] br[3] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_4 bl[4] br[4] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_5 bl[5] br[5] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_6 bl[6] br[6] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_7 bl[7] br[7] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_8 bl[8] br[8] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_9 bl[9] br[9] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_10 bl[10] br[10] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_11 bl[11] br[11] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_12 bl[12] br[12] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_13 bl[13] br[13] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_14 bl[14] br[14] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_15 bl[15] br[15] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_16 bl[16] br[16] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_17 bl[17] br[17] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_18 bl[18] br[18] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_19 bl[19] br[19] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_20 bl[20] br[20] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_21 bl[21] br[21] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_22 bl[22] br[22] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_23 bl[23] br[23] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_24 bl[24] br[24] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_25 bl[25] br[25] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_26 bl[26] br[26] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_27 bl[27] br[27] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_28 bl[28] br[28] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_29 bl[29] br[29] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_30 bl[30] br[30] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_31 bl[31] br[31] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_32 bl[32] br[32] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_33 bl[33] br[33] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_34 bl[34] br[34] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_35 bl[35] br[35] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_36 bl[36] br[36] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_37 bl[37] br[37] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_38 bl[38] br[38] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_39 bl[39] br[39] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_40 bl[40] br[40] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_41 bl[41] br[41] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_42 bl[42] br[42] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_43 bl[43] br[43] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_44 bl[44] br[44] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_45 bl[45] br[45] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_46 bl[46] br[46] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_47 bl[47] br[47] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_48 bl[48] br[48] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_49 bl[49] br[49] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_50 bl[50] br[50] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_51 bl[51] br[51] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_52 bl[52] br[52] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_53 bl[53] br[53] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_54 bl[54] br[54] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_55 bl[55] br[55] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_56 bl[56] br[56] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_57 bl[57] br[57] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_58 bl[58] br[58] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_59 bl[59] br[59] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_60 bl[60] br[60] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_61 bl[61] br[61] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_62 bl[62] br[62] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_63 bl[63] br[63] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_64 bl[64] br[64] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_65 bl[65] br[65] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_66 bl[66] br[66] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_67 bl[67] br[67] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_68 bl[68] br[68] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_69 bl[69] br[69] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_70 bl[70] br[70] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_71 bl[71] br[71] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_72 bl[72] br[72] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_73 bl[73] br[73] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_74 bl[74] br[74] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_75 bl[75] br[75] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_76 bl[76] br[76] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_77 bl[77] br[77] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_78 bl[78] br[78] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_79 bl[79] br[79] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_80 bl[80] br[80] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_81 bl[81] br[81] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_82 bl[82] br[82] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_83 bl[83] br[83] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_84 bl[84] br[84] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_85 bl[85] br[85] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_86 bl[86] br[86] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_87 bl[87] br[87] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_88 bl[88] br[88] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_89 bl[89] br[89] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_90 bl[90] br[90] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_91 bl[91] br[91] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_92 bl[92] br[92] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_93 bl[93] br[93] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_94 bl[94] br[94] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_95 bl[95] br[95] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_96 bl[96] br[96] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_97 bl[97] br[97] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_98 bl[98] br[98] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_99 bl[99] br[99] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_100 bl[100] br[100] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_101 bl[101] br[101] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_102 bl[102] br[102] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_103 bl[103] br[103] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_104 bl[104] br[104] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_105 bl[105] br[105] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_106 bl[106] br[106] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_107 bl[107] br[107] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_108 bl[108] br[108] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_109 bl[109] br[109] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_110 bl[110] br[110] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_111 bl[111] br[111] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_112 bl[112] br[112] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_113 bl[113] br[113] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_114 bl[114] br[114] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_115 bl[115] br[115] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_116 bl[116] br[116] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_117 bl[117] br[117] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_118 bl[118] br[118] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_119 bl[119] br[119] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_120 bl[120] br[120] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_121 bl[121] br[121] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_122 bl[122] br[122] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_123 bl[123] br[123] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_124 bl[124] br[124] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_125 bl[125] br[125] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_126 bl[126] br[126] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_127 bl[127] br[127] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_128 bl[128] br[128] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_129 bl[129] br[129] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_130 bl[130] br[130] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_131 bl[131] br[131] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_132 bl[132] br[132] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_133 bl[133] br[133] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_134 bl[134] br[134] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_135 bl[135] br[135] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_136 bl[136] br[136] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_137 bl[137] br[137] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_138 bl[138] br[138] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_139 bl[139] br[139] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_140 bl[140] br[140] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_141 bl[141] br[141] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_142 bl[142] br[142] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_143 bl[143] br[143] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_144 bl[144] br[144] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_145 bl[145] br[145] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_146 bl[146] br[146] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_147 bl[147] br[147] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_148 bl[148] br[148] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_149 bl[149] br[149] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_150 bl[150] br[150] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_151 bl[151] br[151] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_152 bl[152] br[152] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_153 bl[153] br[153] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_154 bl[154] br[154] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_155 bl[155] br[155] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_156 bl[156] br[156] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_157 bl[157] br[157] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_158 bl[158] br[158] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_159 bl[159] br[159] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_160 bl[160] br[160] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_161 bl[161] br[161] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_162 bl[162] br[162] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_163 bl[163] br[163] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_164 bl[164] br[164] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_165 bl[165] br[165] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_166 bl[166] br[166] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_167 bl[167] br[167] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_168 bl[168] br[168] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_169 bl[169] br[169] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_170 bl[170] br[170] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_171 bl[171] br[171] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_172 bl[172] br[172] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_173 bl[173] br[173] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_174 bl[174] br[174] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_175 bl[175] br[175] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_176 bl[176] br[176] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_177 bl[177] br[177] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_178 bl[178] br[178] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_179 bl[179] br[179] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_180 bl[180] br[180] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_181 bl[181] br[181] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_182 bl[182] br[182] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_183 bl[183] br[183] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_184 bl[184] br[184] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_185 bl[185] br[185] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_186 bl[186] br[186] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_187 bl[187] br[187] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_188 bl[188] br[188] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_189 bl[189] br[189] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_190 bl[190] br[190] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_191 bl[191] br[191] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_192 bl[192] br[192] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_193 bl[193] br[193] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_194 bl[194] br[194] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_195 bl[195] br[195] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_196 bl[196] br[196] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_197 bl[197] br[197] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_198 bl[198] br[198] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_199 bl[199] br[199] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_200 bl[200] br[200] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_201 bl[201] br[201] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_202 bl[202] br[202] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_203 bl[203] br[203] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_204 bl[204] br[204] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_205 bl[205] br[205] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_206 bl[206] br[206] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_207 bl[207] br[207] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_208 bl[208] br[208] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_209 bl[209] br[209] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_210 bl[210] br[210] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_211 bl[211] br[211] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_212 bl[212] br[212] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_213 bl[213] br[213] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_214 bl[214] br[214] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_215 bl[215] br[215] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_216 bl[216] br[216] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_217 bl[217] br[217] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_218 bl[218] br[218] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_219 bl[219] br[219] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_220 bl[220] br[220] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_221 bl[221] br[221] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_222 bl[222] br[222] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_223 bl[223] br[223] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_224 bl[224] br[224] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_225 bl[225] br[225] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_226 bl[226] br[226] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_227 bl[227] br[227] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_228 bl[228] br[228] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_229 bl[229] br[229] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_230 bl[230] br[230] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_231 bl[231] br[231] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_232 bl[232] br[232] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_233 bl[233] br[233] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_234 bl[234] br[234] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_235 bl[235] br[235] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_236 bl[236] br[236] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_237 bl[237] br[237] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_238 bl[238] br[238] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_239 bl[239] br[239] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_240 bl[240] br[240] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_241 bl[241] br[241] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_242 bl[242] br[242] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_243 bl[243] br[243] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_244 bl[244] br[244] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_245 bl[245] br[245] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_246 bl[246] br[246] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_247 bl[247] br[247] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_248 bl[248] br[248] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_249 bl[249] br[249] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_250 bl[250] br[250] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_251 bl[251] br[251] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_252 bl[252] br[252] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_253 bl[253] br[253] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_254 bl[254] br[254] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_255 bl[255] br[255] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_39_0 bl[0] br[0] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_1 bl[1] br[1] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_2 bl[2] br[2] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_3 bl[3] br[3] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_4 bl[4] br[4] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_5 bl[5] br[5] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_6 bl[6] br[6] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_7 bl[7] br[7] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_8 bl[8] br[8] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_9 bl[9] br[9] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_10 bl[10] br[10] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_11 bl[11] br[11] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_12 bl[12] br[12] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_13 bl[13] br[13] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_14 bl[14] br[14] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_15 bl[15] br[15] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_16 bl[16] br[16] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_17 bl[17] br[17] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_18 bl[18] br[18] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_19 bl[19] br[19] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_20 bl[20] br[20] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_21 bl[21] br[21] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_22 bl[22] br[22] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_23 bl[23] br[23] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_24 bl[24] br[24] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_25 bl[25] br[25] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_26 bl[26] br[26] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_27 bl[27] br[27] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_28 bl[28] br[28] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_29 bl[29] br[29] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_30 bl[30] br[30] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_31 bl[31] br[31] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_32 bl[32] br[32] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_33 bl[33] br[33] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_34 bl[34] br[34] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_35 bl[35] br[35] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_36 bl[36] br[36] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_37 bl[37] br[37] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_38 bl[38] br[38] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_39 bl[39] br[39] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_40 bl[40] br[40] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_41 bl[41] br[41] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_42 bl[42] br[42] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_43 bl[43] br[43] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_44 bl[44] br[44] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_45 bl[45] br[45] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_46 bl[46] br[46] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_47 bl[47] br[47] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_48 bl[48] br[48] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_49 bl[49] br[49] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_50 bl[50] br[50] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_51 bl[51] br[51] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_52 bl[52] br[52] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_53 bl[53] br[53] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_54 bl[54] br[54] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_55 bl[55] br[55] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_56 bl[56] br[56] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_57 bl[57] br[57] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_58 bl[58] br[58] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_59 bl[59] br[59] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_60 bl[60] br[60] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_61 bl[61] br[61] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_62 bl[62] br[62] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_63 bl[63] br[63] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_64 bl[64] br[64] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_65 bl[65] br[65] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_66 bl[66] br[66] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_67 bl[67] br[67] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_68 bl[68] br[68] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_69 bl[69] br[69] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_70 bl[70] br[70] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_71 bl[71] br[71] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_72 bl[72] br[72] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_73 bl[73] br[73] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_74 bl[74] br[74] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_75 bl[75] br[75] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_76 bl[76] br[76] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_77 bl[77] br[77] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_78 bl[78] br[78] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_79 bl[79] br[79] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_80 bl[80] br[80] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_81 bl[81] br[81] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_82 bl[82] br[82] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_83 bl[83] br[83] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_84 bl[84] br[84] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_85 bl[85] br[85] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_86 bl[86] br[86] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_87 bl[87] br[87] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_88 bl[88] br[88] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_89 bl[89] br[89] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_90 bl[90] br[90] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_91 bl[91] br[91] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_92 bl[92] br[92] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_93 bl[93] br[93] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_94 bl[94] br[94] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_95 bl[95] br[95] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_96 bl[96] br[96] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_97 bl[97] br[97] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_98 bl[98] br[98] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_99 bl[99] br[99] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_100 bl[100] br[100] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_101 bl[101] br[101] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_102 bl[102] br[102] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_103 bl[103] br[103] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_104 bl[104] br[104] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_105 bl[105] br[105] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_106 bl[106] br[106] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_107 bl[107] br[107] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_108 bl[108] br[108] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_109 bl[109] br[109] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_110 bl[110] br[110] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_111 bl[111] br[111] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_112 bl[112] br[112] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_113 bl[113] br[113] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_114 bl[114] br[114] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_115 bl[115] br[115] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_116 bl[116] br[116] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_117 bl[117] br[117] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_118 bl[118] br[118] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_119 bl[119] br[119] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_120 bl[120] br[120] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_121 bl[121] br[121] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_122 bl[122] br[122] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_123 bl[123] br[123] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_124 bl[124] br[124] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_125 bl[125] br[125] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_126 bl[126] br[126] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_127 bl[127] br[127] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_128 bl[128] br[128] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_129 bl[129] br[129] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_130 bl[130] br[130] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_131 bl[131] br[131] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_132 bl[132] br[132] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_133 bl[133] br[133] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_134 bl[134] br[134] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_135 bl[135] br[135] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_136 bl[136] br[136] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_137 bl[137] br[137] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_138 bl[138] br[138] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_139 bl[139] br[139] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_140 bl[140] br[140] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_141 bl[141] br[141] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_142 bl[142] br[142] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_143 bl[143] br[143] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_144 bl[144] br[144] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_145 bl[145] br[145] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_146 bl[146] br[146] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_147 bl[147] br[147] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_148 bl[148] br[148] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_149 bl[149] br[149] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_150 bl[150] br[150] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_151 bl[151] br[151] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_152 bl[152] br[152] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_153 bl[153] br[153] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_154 bl[154] br[154] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_155 bl[155] br[155] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_156 bl[156] br[156] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_157 bl[157] br[157] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_158 bl[158] br[158] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_159 bl[159] br[159] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_160 bl[160] br[160] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_161 bl[161] br[161] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_162 bl[162] br[162] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_163 bl[163] br[163] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_164 bl[164] br[164] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_165 bl[165] br[165] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_166 bl[166] br[166] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_167 bl[167] br[167] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_168 bl[168] br[168] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_169 bl[169] br[169] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_170 bl[170] br[170] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_171 bl[171] br[171] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_172 bl[172] br[172] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_173 bl[173] br[173] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_174 bl[174] br[174] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_175 bl[175] br[175] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_176 bl[176] br[176] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_177 bl[177] br[177] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_178 bl[178] br[178] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_179 bl[179] br[179] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_180 bl[180] br[180] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_181 bl[181] br[181] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_182 bl[182] br[182] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_183 bl[183] br[183] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_184 bl[184] br[184] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_185 bl[185] br[185] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_186 bl[186] br[186] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_187 bl[187] br[187] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_188 bl[188] br[188] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_189 bl[189] br[189] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_190 bl[190] br[190] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_191 bl[191] br[191] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_192 bl[192] br[192] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_193 bl[193] br[193] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_194 bl[194] br[194] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_195 bl[195] br[195] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_196 bl[196] br[196] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_197 bl[197] br[197] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_198 bl[198] br[198] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_199 bl[199] br[199] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_200 bl[200] br[200] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_201 bl[201] br[201] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_202 bl[202] br[202] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_203 bl[203] br[203] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_204 bl[204] br[204] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_205 bl[205] br[205] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_206 bl[206] br[206] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_207 bl[207] br[207] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_208 bl[208] br[208] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_209 bl[209] br[209] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_210 bl[210] br[210] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_211 bl[211] br[211] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_212 bl[212] br[212] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_213 bl[213] br[213] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_214 bl[214] br[214] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_215 bl[215] br[215] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_216 bl[216] br[216] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_217 bl[217] br[217] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_218 bl[218] br[218] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_219 bl[219] br[219] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_220 bl[220] br[220] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_221 bl[221] br[221] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_222 bl[222] br[222] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_223 bl[223] br[223] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_224 bl[224] br[224] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_225 bl[225] br[225] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_226 bl[226] br[226] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_227 bl[227] br[227] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_228 bl[228] br[228] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_229 bl[229] br[229] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_230 bl[230] br[230] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_231 bl[231] br[231] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_232 bl[232] br[232] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_233 bl[233] br[233] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_234 bl[234] br[234] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_235 bl[235] br[235] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_236 bl[236] br[236] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_237 bl[237] br[237] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_238 bl[238] br[238] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_239 bl[239] br[239] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_240 bl[240] br[240] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_241 bl[241] br[241] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_242 bl[242] br[242] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_243 bl[243] br[243] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_244 bl[244] br[244] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_245 bl[245] br[245] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_246 bl[246] br[246] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_247 bl[247] br[247] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_248 bl[248] br[248] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_249 bl[249] br[249] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_250 bl[250] br[250] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_251 bl[251] br[251] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_252 bl[252] br[252] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_253 bl[253] br[253] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_254 bl[254] br[254] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_255 bl[255] br[255] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_40_0 bl[0] br[0] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_1 bl[1] br[1] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_2 bl[2] br[2] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_3 bl[3] br[3] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_4 bl[4] br[4] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_5 bl[5] br[5] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_6 bl[6] br[6] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_7 bl[7] br[7] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_8 bl[8] br[8] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_9 bl[9] br[9] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_10 bl[10] br[10] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_11 bl[11] br[11] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_12 bl[12] br[12] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_13 bl[13] br[13] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_14 bl[14] br[14] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_15 bl[15] br[15] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_16 bl[16] br[16] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_17 bl[17] br[17] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_18 bl[18] br[18] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_19 bl[19] br[19] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_20 bl[20] br[20] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_21 bl[21] br[21] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_22 bl[22] br[22] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_23 bl[23] br[23] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_24 bl[24] br[24] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_25 bl[25] br[25] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_26 bl[26] br[26] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_27 bl[27] br[27] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_28 bl[28] br[28] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_29 bl[29] br[29] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_30 bl[30] br[30] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_31 bl[31] br[31] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_32 bl[32] br[32] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_33 bl[33] br[33] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_34 bl[34] br[34] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_35 bl[35] br[35] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_36 bl[36] br[36] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_37 bl[37] br[37] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_38 bl[38] br[38] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_39 bl[39] br[39] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_40 bl[40] br[40] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_41 bl[41] br[41] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_42 bl[42] br[42] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_43 bl[43] br[43] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_44 bl[44] br[44] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_45 bl[45] br[45] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_46 bl[46] br[46] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_47 bl[47] br[47] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_48 bl[48] br[48] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_49 bl[49] br[49] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_50 bl[50] br[50] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_51 bl[51] br[51] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_52 bl[52] br[52] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_53 bl[53] br[53] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_54 bl[54] br[54] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_55 bl[55] br[55] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_56 bl[56] br[56] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_57 bl[57] br[57] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_58 bl[58] br[58] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_59 bl[59] br[59] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_60 bl[60] br[60] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_61 bl[61] br[61] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_62 bl[62] br[62] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_63 bl[63] br[63] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_64 bl[64] br[64] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_65 bl[65] br[65] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_66 bl[66] br[66] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_67 bl[67] br[67] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_68 bl[68] br[68] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_69 bl[69] br[69] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_70 bl[70] br[70] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_71 bl[71] br[71] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_72 bl[72] br[72] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_73 bl[73] br[73] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_74 bl[74] br[74] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_75 bl[75] br[75] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_76 bl[76] br[76] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_77 bl[77] br[77] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_78 bl[78] br[78] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_79 bl[79] br[79] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_80 bl[80] br[80] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_81 bl[81] br[81] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_82 bl[82] br[82] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_83 bl[83] br[83] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_84 bl[84] br[84] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_85 bl[85] br[85] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_86 bl[86] br[86] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_87 bl[87] br[87] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_88 bl[88] br[88] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_89 bl[89] br[89] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_90 bl[90] br[90] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_91 bl[91] br[91] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_92 bl[92] br[92] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_93 bl[93] br[93] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_94 bl[94] br[94] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_95 bl[95] br[95] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_96 bl[96] br[96] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_97 bl[97] br[97] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_98 bl[98] br[98] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_99 bl[99] br[99] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_100 bl[100] br[100] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_101 bl[101] br[101] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_102 bl[102] br[102] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_103 bl[103] br[103] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_104 bl[104] br[104] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_105 bl[105] br[105] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_106 bl[106] br[106] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_107 bl[107] br[107] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_108 bl[108] br[108] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_109 bl[109] br[109] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_110 bl[110] br[110] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_111 bl[111] br[111] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_112 bl[112] br[112] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_113 bl[113] br[113] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_114 bl[114] br[114] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_115 bl[115] br[115] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_116 bl[116] br[116] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_117 bl[117] br[117] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_118 bl[118] br[118] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_119 bl[119] br[119] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_120 bl[120] br[120] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_121 bl[121] br[121] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_122 bl[122] br[122] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_123 bl[123] br[123] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_124 bl[124] br[124] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_125 bl[125] br[125] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_126 bl[126] br[126] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_127 bl[127] br[127] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_128 bl[128] br[128] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_129 bl[129] br[129] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_130 bl[130] br[130] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_131 bl[131] br[131] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_132 bl[132] br[132] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_133 bl[133] br[133] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_134 bl[134] br[134] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_135 bl[135] br[135] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_136 bl[136] br[136] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_137 bl[137] br[137] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_138 bl[138] br[138] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_139 bl[139] br[139] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_140 bl[140] br[140] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_141 bl[141] br[141] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_142 bl[142] br[142] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_143 bl[143] br[143] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_144 bl[144] br[144] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_145 bl[145] br[145] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_146 bl[146] br[146] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_147 bl[147] br[147] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_148 bl[148] br[148] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_149 bl[149] br[149] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_150 bl[150] br[150] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_151 bl[151] br[151] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_152 bl[152] br[152] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_153 bl[153] br[153] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_154 bl[154] br[154] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_155 bl[155] br[155] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_156 bl[156] br[156] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_157 bl[157] br[157] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_158 bl[158] br[158] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_159 bl[159] br[159] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_160 bl[160] br[160] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_161 bl[161] br[161] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_162 bl[162] br[162] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_163 bl[163] br[163] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_164 bl[164] br[164] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_165 bl[165] br[165] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_166 bl[166] br[166] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_167 bl[167] br[167] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_168 bl[168] br[168] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_169 bl[169] br[169] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_170 bl[170] br[170] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_171 bl[171] br[171] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_172 bl[172] br[172] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_173 bl[173] br[173] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_174 bl[174] br[174] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_175 bl[175] br[175] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_176 bl[176] br[176] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_177 bl[177] br[177] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_178 bl[178] br[178] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_179 bl[179] br[179] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_180 bl[180] br[180] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_181 bl[181] br[181] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_182 bl[182] br[182] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_183 bl[183] br[183] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_184 bl[184] br[184] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_185 bl[185] br[185] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_186 bl[186] br[186] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_187 bl[187] br[187] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_188 bl[188] br[188] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_189 bl[189] br[189] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_190 bl[190] br[190] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_191 bl[191] br[191] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_192 bl[192] br[192] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_193 bl[193] br[193] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_194 bl[194] br[194] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_195 bl[195] br[195] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_196 bl[196] br[196] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_197 bl[197] br[197] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_198 bl[198] br[198] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_199 bl[199] br[199] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_200 bl[200] br[200] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_201 bl[201] br[201] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_202 bl[202] br[202] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_203 bl[203] br[203] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_204 bl[204] br[204] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_205 bl[205] br[205] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_206 bl[206] br[206] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_207 bl[207] br[207] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_208 bl[208] br[208] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_209 bl[209] br[209] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_210 bl[210] br[210] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_211 bl[211] br[211] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_212 bl[212] br[212] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_213 bl[213] br[213] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_214 bl[214] br[214] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_215 bl[215] br[215] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_216 bl[216] br[216] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_217 bl[217] br[217] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_218 bl[218] br[218] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_219 bl[219] br[219] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_220 bl[220] br[220] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_221 bl[221] br[221] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_222 bl[222] br[222] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_223 bl[223] br[223] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_224 bl[224] br[224] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_225 bl[225] br[225] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_226 bl[226] br[226] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_227 bl[227] br[227] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_228 bl[228] br[228] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_229 bl[229] br[229] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_230 bl[230] br[230] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_231 bl[231] br[231] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_232 bl[232] br[232] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_233 bl[233] br[233] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_234 bl[234] br[234] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_235 bl[235] br[235] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_236 bl[236] br[236] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_237 bl[237] br[237] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_238 bl[238] br[238] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_239 bl[239] br[239] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_240 bl[240] br[240] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_241 bl[241] br[241] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_242 bl[242] br[242] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_243 bl[243] br[243] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_244 bl[244] br[244] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_245 bl[245] br[245] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_246 bl[246] br[246] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_247 bl[247] br[247] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_248 bl[248] br[248] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_249 bl[249] br[249] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_250 bl[250] br[250] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_251 bl[251] br[251] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_252 bl[252] br[252] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_253 bl[253] br[253] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_254 bl[254] br[254] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_255 bl[255] br[255] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_41_0 bl[0] br[0] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_1 bl[1] br[1] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_2 bl[2] br[2] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_3 bl[3] br[3] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_4 bl[4] br[4] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_5 bl[5] br[5] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_6 bl[6] br[6] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_7 bl[7] br[7] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_8 bl[8] br[8] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_9 bl[9] br[9] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_10 bl[10] br[10] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_11 bl[11] br[11] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_12 bl[12] br[12] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_13 bl[13] br[13] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_14 bl[14] br[14] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_15 bl[15] br[15] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_16 bl[16] br[16] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_17 bl[17] br[17] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_18 bl[18] br[18] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_19 bl[19] br[19] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_20 bl[20] br[20] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_21 bl[21] br[21] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_22 bl[22] br[22] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_23 bl[23] br[23] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_24 bl[24] br[24] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_25 bl[25] br[25] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_26 bl[26] br[26] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_27 bl[27] br[27] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_28 bl[28] br[28] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_29 bl[29] br[29] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_30 bl[30] br[30] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_31 bl[31] br[31] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_32 bl[32] br[32] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_33 bl[33] br[33] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_34 bl[34] br[34] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_35 bl[35] br[35] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_36 bl[36] br[36] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_37 bl[37] br[37] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_38 bl[38] br[38] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_39 bl[39] br[39] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_40 bl[40] br[40] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_41 bl[41] br[41] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_42 bl[42] br[42] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_43 bl[43] br[43] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_44 bl[44] br[44] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_45 bl[45] br[45] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_46 bl[46] br[46] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_47 bl[47] br[47] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_48 bl[48] br[48] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_49 bl[49] br[49] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_50 bl[50] br[50] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_51 bl[51] br[51] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_52 bl[52] br[52] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_53 bl[53] br[53] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_54 bl[54] br[54] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_55 bl[55] br[55] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_56 bl[56] br[56] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_57 bl[57] br[57] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_58 bl[58] br[58] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_59 bl[59] br[59] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_60 bl[60] br[60] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_61 bl[61] br[61] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_62 bl[62] br[62] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_63 bl[63] br[63] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_64 bl[64] br[64] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_65 bl[65] br[65] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_66 bl[66] br[66] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_67 bl[67] br[67] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_68 bl[68] br[68] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_69 bl[69] br[69] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_70 bl[70] br[70] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_71 bl[71] br[71] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_72 bl[72] br[72] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_73 bl[73] br[73] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_74 bl[74] br[74] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_75 bl[75] br[75] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_76 bl[76] br[76] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_77 bl[77] br[77] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_78 bl[78] br[78] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_79 bl[79] br[79] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_80 bl[80] br[80] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_81 bl[81] br[81] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_82 bl[82] br[82] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_83 bl[83] br[83] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_84 bl[84] br[84] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_85 bl[85] br[85] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_86 bl[86] br[86] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_87 bl[87] br[87] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_88 bl[88] br[88] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_89 bl[89] br[89] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_90 bl[90] br[90] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_91 bl[91] br[91] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_92 bl[92] br[92] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_93 bl[93] br[93] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_94 bl[94] br[94] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_95 bl[95] br[95] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_96 bl[96] br[96] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_97 bl[97] br[97] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_98 bl[98] br[98] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_99 bl[99] br[99] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_100 bl[100] br[100] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_101 bl[101] br[101] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_102 bl[102] br[102] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_103 bl[103] br[103] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_104 bl[104] br[104] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_105 bl[105] br[105] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_106 bl[106] br[106] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_107 bl[107] br[107] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_108 bl[108] br[108] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_109 bl[109] br[109] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_110 bl[110] br[110] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_111 bl[111] br[111] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_112 bl[112] br[112] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_113 bl[113] br[113] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_114 bl[114] br[114] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_115 bl[115] br[115] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_116 bl[116] br[116] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_117 bl[117] br[117] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_118 bl[118] br[118] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_119 bl[119] br[119] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_120 bl[120] br[120] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_121 bl[121] br[121] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_122 bl[122] br[122] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_123 bl[123] br[123] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_124 bl[124] br[124] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_125 bl[125] br[125] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_126 bl[126] br[126] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_127 bl[127] br[127] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_128 bl[128] br[128] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_129 bl[129] br[129] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_130 bl[130] br[130] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_131 bl[131] br[131] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_132 bl[132] br[132] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_133 bl[133] br[133] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_134 bl[134] br[134] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_135 bl[135] br[135] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_136 bl[136] br[136] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_137 bl[137] br[137] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_138 bl[138] br[138] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_139 bl[139] br[139] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_140 bl[140] br[140] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_141 bl[141] br[141] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_142 bl[142] br[142] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_143 bl[143] br[143] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_144 bl[144] br[144] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_145 bl[145] br[145] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_146 bl[146] br[146] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_147 bl[147] br[147] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_148 bl[148] br[148] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_149 bl[149] br[149] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_150 bl[150] br[150] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_151 bl[151] br[151] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_152 bl[152] br[152] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_153 bl[153] br[153] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_154 bl[154] br[154] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_155 bl[155] br[155] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_156 bl[156] br[156] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_157 bl[157] br[157] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_158 bl[158] br[158] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_159 bl[159] br[159] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_160 bl[160] br[160] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_161 bl[161] br[161] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_162 bl[162] br[162] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_163 bl[163] br[163] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_164 bl[164] br[164] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_165 bl[165] br[165] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_166 bl[166] br[166] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_167 bl[167] br[167] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_168 bl[168] br[168] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_169 bl[169] br[169] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_170 bl[170] br[170] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_171 bl[171] br[171] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_172 bl[172] br[172] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_173 bl[173] br[173] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_174 bl[174] br[174] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_175 bl[175] br[175] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_176 bl[176] br[176] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_177 bl[177] br[177] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_178 bl[178] br[178] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_179 bl[179] br[179] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_180 bl[180] br[180] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_181 bl[181] br[181] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_182 bl[182] br[182] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_183 bl[183] br[183] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_184 bl[184] br[184] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_185 bl[185] br[185] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_186 bl[186] br[186] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_187 bl[187] br[187] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_188 bl[188] br[188] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_189 bl[189] br[189] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_190 bl[190] br[190] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_191 bl[191] br[191] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_192 bl[192] br[192] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_193 bl[193] br[193] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_194 bl[194] br[194] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_195 bl[195] br[195] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_196 bl[196] br[196] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_197 bl[197] br[197] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_198 bl[198] br[198] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_199 bl[199] br[199] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_200 bl[200] br[200] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_201 bl[201] br[201] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_202 bl[202] br[202] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_203 bl[203] br[203] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_204 bl[204] br[204] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_205 bl[205] br[205] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_206 bl[206] br[206] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_207 bl[207] br[207] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_208 bl[208] br[208] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_209 bl[209] br[209] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_210 bl[210] br[210] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_211 bl[211] br[211] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_212 bl[212] br[212] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_213 bl[213] br[213] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_214 bl[214] br[214] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_215 bl[215] br[215] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_216 bl[216] br[216] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_217 bl[217] br[217] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_218 bl[218] br[218] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_219 bl[219] br[219] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_220 bl[220] br[220] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_221 bl[221] br[221] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_222 bl[222] br[222] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_223 bl[223] br[223] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_224 bl[224] br[224] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_225 bl[225] br[225] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_226 bl[226] br[226] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_227 bl[227] br[227] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_228 bl[228] br[228] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_229 bl[229] br[229] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_230 bl[230] br[230] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_231 bl[231] br[231] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_232 bl[232] br[232] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_233 bl[233] br[233] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_234 bl[234] br[234] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_235 bl[235] br[235] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_236 bl[236] br[236] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_237 bl[237] br[237] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_238 bl[238] br[238] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_239 bl[239] br[239] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_240 bl[240] br[240] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_241 bl[241] br[241] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_242 bl[242] br[242] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_243 bl[243] br[243] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_244 bl[244] br[244] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_245 bl[245] br[245] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_246 bl[246] br[246] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_247 bl[247] br[247] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_248 bl[248] br[248] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_249 bl[249] br[249] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_250 bl[250] br[250] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_251 bl[251] br[251] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_252 bl[252] br[252] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_253 bl[253] br[253] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_254 bl[254] br[254] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_255 bl[255] br[255] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_42_0 bl[0] br[0] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_1 bl[1] br[1] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_2 bl[2] br[2] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_3 bl[3] br[3] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_4 bl[4] br[4] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_5 bl[5] br[5] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_6 bl[6] br[6] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_7 bl[7] br[7] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_8 bl[8] br[8] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_9 bl[9] br[9] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_10 bl[10] br[10] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_11 bl[11] br[11] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_12 bl[12] br[12] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_13 bl[13] br[13] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_14 bl[14] br[14] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_15 bl[15] br[15] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_16 bl[16] br[16] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_17 bl[17] br[17] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_18 bl[18] br[18] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_19 bl[19] br[19] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_20 bl[20] br[20] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_21 bl[21] br[21] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_22 bl[22] br[22] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_23 bl[23] br[23] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_24 bl[24] br[24] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_25 bl[25] br[25] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_26 bl[26] br[26] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_27 bl[27] br[27] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_28 bl[28] br[28] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_29 bl[29] br[29] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_30 bl[30] br[30] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_31 bl[31] br[31] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_32 bl[32] br[32] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_33 bl[33] br[33] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_34 bl[34] br[34] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_35 bl[35] br[35] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_36 bl[36] br[36] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_37 bl[37] br[37] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_38 bl[38] br[38] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_39 bl[39] br[39] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_40 bl[40] br[40] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_41 bl[41] br[41] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_42 bl[42] br[42] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_43 bl[43] br[43] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_44 bl[44] br[44] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_45 bl[45] br[45] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_46 bl[46] br[46] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_47 bl[47] br[47] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_48 bl[48] br[48] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_49 bl[49] br[49] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_50 bl[50] br[50] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_51 bl[51] br[51] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_52 bl[52] br[52] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_53 bl[53] br[53] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_54 bl[54] br[54] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_55 bl[55] br[55] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_56 bl[56] br[56] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_57 bl[57] br[57] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_58 bl[58] br[58] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_59 bl[59] br[59] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_60 bl[60] br[60] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_61 bl[61] br[61] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_62 bl[62] br[62] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_63 bl[63] br[63] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_64 bl[64] br[64] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_65 bl[65] br[65] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_66 bl[66] br[66] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_67 bl[67] br[67] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_68 bl[68] br[68] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_69 bl[69] br[69] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_70 bl[70] br[70] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_71 bl[71] br[71] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_72 bl[72] br[72] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_73 bl[73] br[73] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_74 bl[74] br[74] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_75 bl[75] br[75] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_76 bl[76] br[76] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_77 bl[77] br[77] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_78 bl[78] br[78] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_79 bl[79] br[79] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_80 bl[80] br[80] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_81 bl[81] br[81] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_82 bl[82] br[82] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_83 bl[83] br[83] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_84 bl[84] br[84] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_85 bl[85] br[85] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_86 bl[86] br[86] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_87 bl[87] br[87] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_88 bl[88] br[88] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_89 bl[89] br[89] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_90 bl[90] br[90] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_91 bl[91] br[91] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_92 bl[92] br[92] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_93 bl[93] br[93] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_94 bl[94] br[94] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_95 bl[95] br[95] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_96 bl[96] br[96] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_97 bl[97] br[97] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_98 bl[98] br[98] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_99 bl[99] br[99] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_100 bl[100] br[100] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_101 bl[101] br[101] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_102 bl[102] br[102] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_103 bl[103] br[103] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_104 bl[104] br[104] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_105 bl[105] br[105] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_106 bl[106] br[106] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_107 bl[107] br[107] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_108 bl[108] br[108] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_109 bl[109] br[109] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_110 bl[110] br[110] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_111 bl[111] br[111] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_112 bl[112] br[112] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_113 bl[113] br[113] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_114 bl[114] br[114] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_115 bl[115] br[115] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_116 bl[116] br[116] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_117 bl[117] br[117] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_118 bl[118] br[118] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_119 bl[119] br[119] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_120 bl[120] br[120] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_121 bl[121] br[121] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_122 bl[122] br[122] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_123 bl[123] br[123] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_124 bl[124] br[124] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_125 bl[125] br[125] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_126 bl[126] br[126] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_127 bl[127] br[127] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_128 bl[128] br[128] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_129 bl[129] br[129] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_130 bl[130] br[130] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_131 bl[131] br[131] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_132 bl[132] br[132] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_133 bl[133] br[133] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_134 bl[134] br[134] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_135 bl[135] br[135] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_136 bl[136] br[136] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_137 bl[137] br[137] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_138 bl[138] br[138] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_139 bl[139] br[139] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_140 bl[140] br[140] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_141 bl[141] br[141] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_142 bl[142] br[142] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_143 bl[143] br[143] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_144 bl[144] br[144] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_145 bl[145] br[145] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_146 bl[146] br[146] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_147 bl[147] br[147] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_148 bl[148] br[148] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_149 bl[149] br[149] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_150 bl[150] br[150] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_151 bl[151] br[151] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_152 bl[152] br[152] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_153 bl[153] br[153] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_154 bl[154] br[154] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_155 bl[155] br[155] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_156 bl[156] br[156] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_157 bl[157] br[157] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_158 bl[158] br[158] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_159 bl[159] br[159] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_160 bl[160] br[160] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_161 bl[161] br[161] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_162 bl[162] br[162] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_163 bl[163] br[163] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_164 bl[164] br[164] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_165 bl[165] br[165] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_166 bl[166] br[166] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_167 bl[167] br[167] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_168 bl[168] br[168] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_169 bl[169] br[169] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_170 bl[170] br[170] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_171 bl[171] br[171] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_172 bl[172] br[172] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_173 bl[173] br[173] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_174 bl[174] br[174] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_175 bl[175] br[175] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_176 bl[176] br[176] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_177 bl[177] br[177] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_178 bl[178] br[178] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_179 bl[179] br[179] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_180 bl[180] br[180] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_181 bl[181] br[181] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_182 bl[182] br[182] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_183 bl[183] br[183] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_184 bl[184] br[184] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_185 bl[185] br[185] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_186 bl[186] br[186] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_187 bl[187] br[187] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_188 bl[188] br[188] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_189 bl[189] br[189] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_190 bl[190] br[190] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_191 bl[191] br[191] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_192 bl[192] br[192] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_193 bl[193] br[193] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_194 bl[194] br[194] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_195 bl[195] br[195] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_196 bl[196] br[196] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_197 bl[197] br[197] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_198 bl[198] br[198] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_199 bl[199] br[199] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_200 bl[200] br[200] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_201 bl[201] br[201] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_202 bl[202] br[202] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_203 bl[203] br[203] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_204 bl[204] br[204] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_205 bl[205] br[205] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_206 bl[206] br[206] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_207 bl[207] br[207] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_208 bl[208] br[208] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_209 bl[209] br[209] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_210 bl[210] br[210] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_211 bl[211] br[211] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_212 bl[212] br[212] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_213 bl[213] br[213] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_214 bl[214] br[214] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_215 bl[215] br[215] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_216 bl[216] br[216] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_217 bl[217] br[217] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_218 bl[218] br[218] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_219 bl[219] br[219] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_220 bl[220] br[220] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_221 bl[221] br[221] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_222 bl[222] br[222] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_223 bl[223] br[223] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_224 bl[224] br[224] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_225 bl[225] br[225] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_226 bl[226] br[226] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_227 bl[227] br[227] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_228 bl[228] br[228] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_229 bl[229] br[229] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_230 bl[230] br[230] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_231 bl[231] br[231] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_232 bl[232] br[232] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_233 bl[233] br[233] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_234 bl[234] br[234] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_235 bl[235] br[235] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_236 bl[236] br[236] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_237 bl[237] br[237] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_238 bl[238] br[238] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_239 bl[239] br[239] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_240 bl[240] br[240] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_241 bl[241] br[241] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_242 bl[242] br[242] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_243 bl[243] br[243] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_244 bl[244] br[244] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_245 bl[245] br[245] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_246 bl[246] br[246] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_247 bl[247] br[247] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_248 bl[248] br[248] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_249 bl[249] br[249] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_250 bl[250] br[250] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_251 bl[251] br[251] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_252 bl[252] br[252] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_253 bl[253] br[253] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_254 bl[254] br[254] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_255 bl[255] br[255] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_43_0 bl[0] br[0] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_1 bl[1] br[1] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_2 bl[2] br[2] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_3 bl[3] br[3] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_4 bl[4] br[4] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_5 bl[5] br[5] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_6 bl[6] br[6] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_7 bl[7] br[7] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_8 bl[8] br[8] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_9 bl[9] br[9] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_10 bl[10] br[10] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_11 bl[11] br[11] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_12 bl[12] br[12] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_13 bl[13] br[13] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_14 bl[14] br[14] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_15 bl[15] br[15] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_16 bl[16] br[16] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_17 bl[17] br[17] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_18 bl[18] br[18] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_19 bl[19] br[19] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_20 bl[20] br[20] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_21 bl[21] br[21] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_22 bl[22] br[22] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_23 bl[23] br[23] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_24 bl[24] br[24] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_25 bl[25] br[25] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_26 bl[26] br[26] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_27 bl[27] br[27] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_28 bl[28] br[28] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_29 bl[29] br[29] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_30 bl[30] br[30] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_31 bl[31] br[31] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_32 bl[32] br[32] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_33 bl[33] br[33] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_34 bl[34] br[34] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_35 bl[35] br[35] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_36 bl[36] br[36] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_37 bl[37] br[37] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_38 bl[38] br[38] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_39 bl[39] br[39] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_40 bl[40] br[40] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_41 bl[41] br[41] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_42 bl[42] br[42] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_43 bl[43] br[43] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_44 bl[44] br[44] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_45 bl[45] br[45] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_46 bl[46] br[46] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_47 bl[47] br[47] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_48 bl[48] br[48] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_49 bl[49] br[49] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_50 bl[50] br[50] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_51 bl[51] br[51] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_52 bl[52] br[52] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_53 bl[53] br[53] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_54 bl[54] br[54] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_55 bl[55] br[55] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_56 bl[56] br[56] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_57 bl[57] br[57] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_58 bl[58] br[58] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_59 bl[59] br[59] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_60 bl[60] br[60] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_61 bl[61] br[61] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_62 bl[62] br[62] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_63 bl[63] br[63] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_64 bl[64] br[64] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_65 bl[65] br[65] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_66 bl[66] br[66] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_67 bl[67] br[67] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_68 bl[68] br[68] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_69 bl[69] br[69] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_70 bl[70] br[70] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_71 bl[71] br[71] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_72 bl[72] br[72] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_73 bl[73] br[73] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_74 bl[74] br[74] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_75 bl[75] br[75] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_76 bl[76] br[76] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_77 bl[77] br[77] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_78 bl[78] br[78] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_79 bl[79] br[79] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_80 bl[80] br[80] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_81 bl[81] br[81] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_82 bl[82] br[82] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_83 bl[83] br[83] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_84 bl[84] br[84] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_85 bl[85] br[85] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_86 bl[86] br[86] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_87 bl[87] br[87] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_88 bl[88] br[88] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_89 bl[89] br[89] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_90 bl[90] br[90] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_91 bl[91] br[91] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_92 bl[92] br[92] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_93 bl[93] br[93] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_94 bl[94] br[94] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_95 bl[95] br[95] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_96 bl[96] br[96] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_97 bl[97] br[97] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_98 bl[98] br[98] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_99 bl[99] br[99] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_100 bl[100] br[100] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_101 bl[101] br[101] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_102 bl[102] br[102] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_103 bl[103] br[103] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_104 bl[104] br[104] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_105 bl[105] br[105] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_106 bl[106] br[106] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_107 bl[107] br[107] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_108 bl[108] br[108] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_109 bl[109] br[109] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_110 bl[110] br[110] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_111 bl[111] br[111] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_112 bl[112] br[112] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_113 bl[113] br[113] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_114 bl[114] br[114] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_115 bl[115] br[115] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_116 bl[116] br[116] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_117 bl[117] br[117] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_118 bl[118] br[118] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_119 bl[119] br[119] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_120 bl[120] br[120] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_121 bl[121] br[121] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_122 bl[122] br[122] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_123 bl[123] br[123] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_124 bl[124] br[124] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_125 bl[125] br[125] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_126 bl[126] br[126] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_127 bl[127] br[127] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_128 bl[128] br[128] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_129 bl[129] br[129] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_130 bl[130] br[130] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_131 bl[131] br[131] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_132 bl[132] br[132] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_133 bl[133] br[133] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_134 bl[134] br[134] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_135 bl[135] br[135] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_136 bl[136] br[136] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_137 bl[137] br[137] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_138 bl[138] br[138] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_139 bl[139] br[139] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_140 bl[140] br[140] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_141 bl[141] br[141] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_142 bl[142] br[142] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_143 bl[143] br[143] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_144 bl[144] br[144] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_145 bl[145] br[145] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_146 bl[146] br[146] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_147 bl[147] br[147] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_148 bl[148] br[148] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_149 bl[149] br[149] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_150 bl[150] br[150] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_151 bl[151] br[151] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_152 bl[152] br[152] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_153 bl[153] br[153] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_154 bl[154] br[154] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_155 bl[155] br[155] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_156 bl[156] br[156] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_157 bl[157] br[157] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_158 bl[158] br[158] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_159 bl[159] br[159] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_160 bl[160] br[160] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_161 bl[161] br[161] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_162 bl[162] br[162] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_163 bl[163] br[163] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_164 bl[164] br[164] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_165 bl[165] br[165] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_166 bl[166] br[166] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_167 bl[167] br[167] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_168 bl[168] br[168] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_169 bl[169] br[169] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_170 bl[170] br[170] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_171 bl[171] br[171] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_172 bl[172] br[172] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_173 bl[173] br[173] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_174 bl[174] br[174] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_175 bl[175] br[175] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_176 bl[176] br[176] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_177 bl[177] br[177] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_178 bl[178] br[178] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_179 bl[179] br[179] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_180 bl[180] br[180] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_181 bl[181] br[181] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_182 bl[182] br[182] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_183 bl[183] br[183] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_184 bl[184] br[184] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_185 bl[185] br[185] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_186 bl[186] br[186] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_187 bl[187] br[187] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_188 bl[188] br[188] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_189 bl[189] br[189] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_190 bl[190] br[190] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_191 bl[191] br[191] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_192 bl[192] br[192] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_193 bl[193] br[193] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_194 bl[194] br[194] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_195 bl[195] br[195] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_196 bl[196] br[196] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_197 bl[197] br[197] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_198 bl[198] br[198] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_199 bl[199] br[199] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_200 bl[200] br[200] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_201 bl[201] br[201] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_202 bl[202] br[202] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_203 bl[203] br[203] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_204 bl[204] br[204] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_205 bl[205] br[205] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_206 bl[206] br[206] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_207 bl[207] br[207] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_208 bl[208] br[208] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_209 bl[209] br[209] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_210 bl[210] br[210] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_211 bl[211] br[211] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_212 bl[212] br[212] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_213 bl[213] br[213] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_214 bl[214] br[214] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_215 bl[215] br[215] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_216 bl[216] br[216] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_217 bl[217] br[217] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_218 bl[218] br[218] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_219 bl[219] br[219] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_220 bl[220] br[220] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_221 bl[221] br[221] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_222 bl[222] br[222] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_223 bl[223] br[223] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_224 bl[224] br[224] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_225 bl[225] br[225] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_226 bl[226] br[226] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_227 bl[227] br[227] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_228 bl[228] br[228] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_229 bl[229] br[229] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_230 bl[230] br[230] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_231 bl[231] br[231] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_232 bl[232] br[232] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_233 bl[233] br[233] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_234 bl[234] br[234] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_235 bl[235] br[235] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_236 bl[236] br[236] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_237 bl[237] br[237] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_238 bl[238] br[238] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_239 bl[239] br[239] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_240 bl[240] br[240] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_241 bl[241] br[241] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_242 bl[242] br[242] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_243 bl[243] br[243] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_244 bl[244] br[244] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_245 bl[245] br[245] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_246 bl[246] br[246] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_247 bl[247] br[247] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_248 bl[248] br[248] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_249 bl[249] br[249] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_250 bl[250] br[250] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_251 bl[251] br[251] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_252 bl[252] br[252] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_253 bl[253] br[253] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_254 bl[254] br[254] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_255 bl[255] br[255] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_44_0 bl[0] br[0] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_1 bl[1] br[1] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_2 bl[2] br[2] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_3 bl[3] br[3] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_4 bl[4] br[4] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_5 bl[5] br[5] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_6 bl[6] br[6] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_7 bl[7] br[7] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_8 bl[8] br[8] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_9 bl[9] br[9] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_10 bl[10] br[10] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_11 bl[11] br[11] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_12 bl[12] br[12] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_13 bl[13] br[13] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_14 bl[14] br[14] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_15 bl[15] br[15] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_16 bl[16] br[16] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_17 bl[17] br[17] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_18 bl[18] br[18] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_19 bl[19] br[19] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_20 bl[20] br[20] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_21 bl[21] br[21] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_22 bl[22] br[22] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_23 bl[23] br[23] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_24 bl[24] br[24] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_25 bl[25] br[25] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_26 bl[26] br[26] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_27 bl[27] br[27] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_28 bl[28] br[28] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_29 bl[29] br[29] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_30 bl[30] br[30] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_31 bl[31] br[31] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_32 bl[32] br[32] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_33 bl[33] br[33] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_34 bl[34] br[34] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_35 bl[35] br[35] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_36 bl[36] br[36] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_37 bl[37] br[37] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_38 bl[38] br[38] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_39 bl[39] br[39] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_40 bl[40] br[40] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_41 bl[41] br[41] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_42 bl[42] br[42] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_43 bl[43] br[43] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_44 bl[44] br[44] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_45 bl[45] br[45] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_46 bl[46] br[46] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_47 bl[47] br[47] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_48 bl[48] br[48] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_49 bl[49] br[49] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_50 bl[50] br[50] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_51 bl[51] br[51] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_52 bl[52] br[52] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_53 bl[53] br[53] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_54 bl[54] br[54] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_55 bl[55] br[55] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_56 bl[56] br[56] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_57 bl[57] br[57] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_58 bl[58] br[58] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_59 bl[59] br[59] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_60 bl[60] br[60] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_61 bl[61] br[61] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_62 bl[62] br[62] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_63 bl[63] br[63] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_64 bl[64] br[64] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_65 bl[65] br[65] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_66 bl[66] br[66] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_67 bl[67] br[67] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_68 bl[68] br[68] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_69 bl[69] br[69] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_70 bl[70] br[70] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_71 bl[71] br[71] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_72 bl[72] br[72] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_73 bl[73] br[73] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_74 bl[74] br[74] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_75 bl[75] br[75] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_76 bl[76] br[76] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_77 bl[77] br[77] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_78 bl[78] br[78] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_79 bl[79] br[79] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_80 bl[80] br[80] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_81 bl[81] br[81] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_82 bl[82] br[82] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_83 bl[83] br[83] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_84 bl[84] br[84] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_85 bl[85] br[85] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_86 bl[86] br[86] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_87 bl[87] br[87] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_88 bl[88] br[88] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_89 bl[89] br[89] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_90 bl[90] br[90] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_91 bl[91] br[91] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_92 bl[92] br[92] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_93 bl[93] br[93] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_94 bl[94] br[94] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_95 bl[95] br[95] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_96 bl[96] br[96] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_97 bl[97] br[97] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_98 bl[98] br[98] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_99 bl[99] br[99] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_100 bl[100] br[100] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_101 bl[101] br[101] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_102 bl[102] br[102] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_103 bl[103] br[103] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_104 bl[104] br[104] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_105 bl[105] br[105] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_106 bl[106] br[106] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_107 bl[107] br[107] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_108 bl[108] br[108] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_109 bl[109] br[109] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_110 bl[110] br[110] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_111 bl[111] br[111] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_112 bl[112] br[112] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_113 bl[113] br[113] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_114 bl[114] br[114] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_115 bl[115] br[115] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_116 bl[116] br[116] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_117 bl[117] br[117] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_118 bl[118] br[118] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_119 bl[119] br[119] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_120 bl[120] br[120] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_121 bl[121] br[121] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_122 bl[122] br[122] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_123 bl[123] br[123] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_124 bl[124] br[124] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_125 bl[125] br[125] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_126 bl[126] br[126] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_127 bl[127] br[127] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_128 bl[128] br[128] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_129 bl[129] br[129] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_130 bl[130] br[130] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_131 bl[131] br[131] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_132 bl[132] br[132] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_133 bl[133] br[133] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_134 bl[134] br[134] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_135 bl[135] br[135] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_136 bl[136] br[136] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_137 bl[137] br[137] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_138 bl[138] br[138] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_139 bl[139] br[139] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_140 bl[140] br[140] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_141 bl[141] br[141] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_142 bl[142] br[142] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_143 bl[143] br[143] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_144 bl[144] br[144] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_145 bl[145] br[145] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_146 bl[146] br[146] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_147 bl[147] br[147] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_148 bl[148] br[148] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_149 bl[149] br[149] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_150 bl[150] br[150] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_151 bl[151] br[151] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_152 bl[152] br[152] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_153 bl[153] br[153] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_154 bl[154] br[154] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_155 bl[155] br[155] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_156 bl[156] br[156] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_157 bl[157] br[157] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_158 bl[158] br[158] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_159 bl[159] br[159] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_160 bl[160] br[160] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_161 bl[161] br[161] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_162 bl[162] br[162] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_163 bl[163] br[163] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_164 bl[164] br[164] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_165 bl[165] br[165] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_166 bl[166] br[166] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_167 bl[167] br[167] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_168 bl[168] br[168] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_169 bl[169] br[169] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_170 bl[170] br[170] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_171 bl[171] br[171] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_172 bl[172] br[172] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_173 bl[173] br[173] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_174 bl[174] br[174] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_175 bl[175] br[175] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_176 bl[176] br[176] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_177 bl[177] br[177] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_178 bl[178] br[178] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_179 bl[179] br[179] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_180 bl[180] br[180] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_181 bl[181] br[181] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_182 bl[182] br[182] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_183 bl[183] br[183] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_184 bl[184] br[184] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_185 bl[185] br[185] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_186 bl[186] br[186] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_187 bl[187] br[187] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_188 bl[188] br[188] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_189 bl[189] br[189] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_190 bl[190] br[190] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_191 bl[191] br[191] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_192 bl[192] br[192] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_193 bl[193] br[193] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_194 bl[194] br[194] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_195 bl[195] br[195] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_196 bl[196] br[196] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_197 bl[197] br[197] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_198 bl[198] br[198] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_199 bl[199] br[199] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_200 bl[200] br[200] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_201 bl[201] br[201] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_202 bl[202] br[202] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_203 bl[203] br[203] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_204 bl[204] br[204] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_205 bl[205] br[205] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_206 bl[206] br[206] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_207 bl[207] br[207] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_208 bl[208] br[208] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_209 bl[209] br[209] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_210 bl[210] br[210] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_211 bl[211] br[211] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_212 bl[212] br[212] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_213 bl[213] br[213] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_214 bl[214] br[214] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_215 bl[215] br[215] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_216 bl[216] br[216] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_217 bl[217] br[217] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_218 bl[218] br[218] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_219 bl[219] br[219] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_220 bl[220] br[220] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_221 bl[221] br[221] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_222 bl[222] br[222] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_223 bl[223] br[223] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_224 bl[224] br[224] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_225 bl[225] br[225] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_226 bl[226] br[226] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_227 bl[227] br[227] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_228 bl[228] br[228] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_229 bl[229] br[229] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_230 bl[230] br[230] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_231 bl[231] br[231] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_232 bl[232] br[232] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_233 bl[233] br[233] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_234 bl[234] br[234] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_235 bl[235] br[235] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_236 bl[236] br[236] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_237 bl[237] br[237] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_238 bl[238] br[238] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_239 bl[239] br[239] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_240 bl[240] br[240] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_241 bl[241] br[241] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_242 bl[242] br[242] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_243 bl[243] br[243] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_244 bl[244] br[244] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_245 bl[245] br[245] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_246 bl[246] br[246] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_247 bl[247] br[247] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_248 bl[248] br[248] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_249 bl[249] br[249] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_250 bl[250] br[250] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_251 bl[251] br[251] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_252 bl[252] br[252] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_253 bl[253] br[253] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_254 bl[254] br[254] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_255 bl[255] br[255] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_45_0 bl[0] br[0] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_1 bl[1] br[1] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_2 bl[2] br[2] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_3 bl[3] br[3] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_4 bl[4] br[4] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_5 bl[5] br[5] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_6 bl[6] br[6] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_7 bl[7] br[7] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_8 bl[8] br[8] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_9 bl[9] br[9] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_10 bl[10] br[10] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_11 bl[11] br[11] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_12 bl[12] br[12] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_13 bl[13] br[13] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_14 bl[14] br[14] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_15 bl[15] br[15] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_16 bl[16] br[16] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_17 bl[17] br[17] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_18 bl[18] br[18] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_19 bl[19] br[19] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_20 bl[20] br[20] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_21 bl[21] br[21] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_22 bl[22] br[22] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_23 bl[23] br[23] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_24 bl[24] br[24] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_25 bl[25] br[25] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_26 bl[26] br[26] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_27 bl[27] br[27] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_28 bl[28] br[28] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_29 bl[29] br[29] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_30 bl[30] br[30] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_31 bl[31] br[31] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_32 bl[32] br[32] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_33 bl[33] br[33] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_34 bl[34] br[34] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_35 bl[35] br[35] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_36 bl[36] br[36] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_37 bl[37] br[37] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_38 bl[38] br[38] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_39 bl[39] br[39] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_40 bl[40] br[40] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_41 bl[41] br[41] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_42 bl[42] br[42] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_43 bl[43] br[43] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_44 bl[44] br[44] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_45 bl[45] br[45] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_46 bl[46] br[46] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_47 bl[47] br[47] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_48 bl[48] br[48] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_49 bl[49] br[49] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_50 bl[50] br[50] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_51 bl[51] br[51] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_52 bl[52] br[52] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_53 bl[53] br[53] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_54 bl[54] br[54] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_55 bl[55] br[55] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_56 bl[56] br[56] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_57 bl[57] br[57] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_58 bl[58] br[58] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_59 bl[59] br[59] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_60 bl[60] br[60] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_61 bl[61] br[61] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_62 bl[62] br[62] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_63 bl[63] br[63] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_64 bl[64] br[64] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_65 bl[65] br[65] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_66 bl[66] br[66] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_67 bl[67] br[67] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_68 bl[68] br[68] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_69 bl[69] br[69] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_70 bl[70] br[70] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_71 bl[71] br[71] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_72 bl[72] br[72] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_73 bl[73] br[73] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_74 bl[74] br[74] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_75 bl[75] br[75] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_76 bl[76] br[76] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_77 bl[77] br[77] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_78 bl[78] br[78] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_79 bl[79] br[79] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_80 bl[80] br[80] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_81 bl[81] br[81] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_82 bl[82] br[82] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_83 bl[83] br[83] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_84 bl[84] br[84] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_85 bl[85] br[85] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_86 bl[86] br[86] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_87 bl[87] br[87] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_88 bl[88] br[88] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_89 bl[89] br[89] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_90 bl[90] br[90] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_91 bl[91] br[91] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_92 bl[92] br[92] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_93 bl[93] br[93] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_94 bl[94] br[94] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_95 bl[95] br[95] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_96 bl[96] br[96] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_97 bl[97] br[97] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_98 bl[98] br[98] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_99 bl[99] br[99] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_100 bl[100] br[100] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_101 bl[101] br[101] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_102 bl[102] br[102] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_103 bl[103] br[103] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_104 bl[104] br[104] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_105 bl[105] br[105] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_106 bl[106] br[106] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_107 bl[107] br[107] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_108 bl[108] br[108] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_109 bl[109] br[109] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_110 bl[110] br[110] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_111 bl[111] br[111] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_112 bl[112] br[112] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_113 bl[113] br[113] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_114 bl[114] br[114] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_115 bl[115] br[115] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_116 bl[116] br[116] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_117 bl[117] br[117] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_118 bl[118] br[118] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_119 bl[119] br[119] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_120 bl[120] br[120] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_121 bl[121] br[121] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_122 bl[122] br[122] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_123 bl[123] br[123] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_124 bl[124] br[124] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_125 bl[125] br[125] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_126 bl[126] br[126] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_127 bl[127] br[127] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_128 bl[128] br[128] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_129 bl[129] br[129] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_130 bl[130] br[130] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_131 bl[131] br[131] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_132 bl[132] br[132] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_133 bl[133] br[133] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_134 bl[134] br[134] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_135 bl[135] br[135] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_136 bl[136] br[136] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_137 bl[137] br[137] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_138 bl[138] br[138] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_139 bl[139] br[139] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_140 bl[140] br[140] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_141 bl[141] br[141] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_142 bl[142] br[142] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_143 bl[143] br[143] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_144 bl[144] br[144] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_145 bl[145] br[145] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_146 bl[146] br[146] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_147 bl[147] br[147] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_148 bl[148] br[148] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_149 bl[149] br[149] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_150 bl[150] br[150] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_151 bl[151] br[151] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_152 bl[152] br[152] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_153 bl[153] br[153] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_154 bl[154] br[154] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_155 bl[155] br[155] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_156 bl[156] br[156] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_157 bl[157] br[157] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_158 bl[158] br[158] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_159 bl[159] br[159] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_160 bl[160] br[160] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_161 bl[161] br[161] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_162 bl[162] br[162] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_163 bl[163] br[163] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_164 bl[164] br[164] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_165 bl[165] br[165] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_166 bl[166] br[166] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_167 bl[167] br[167] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_168 bl[168] br[168] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_169 bl[169] br[169] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_170 bl[170] br[170] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_171 bl[171] br[171] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_172 bl[172] br[172] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_173 bl[173] br[173] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_174 bl[174] br[174] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_175 bl[175] br[175] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_176 bl[176] br[176] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_177 bl[177] br[177] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_178 bl[178] br[178] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_179 bl[179] br[179] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_180 bl[180] br[180] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_181 bl[181] br[181] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_182 bl[182] br[182] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_183 bl[183] br[183] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_184 bl[184] br[184] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_185 bl[185] br[185] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_186 bl[186] br[186] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_187 bl[187] br[187] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_188 bl[188] br[188] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_189 bl[189] br[189] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_190 bl[190] br[190] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_191 bl[191] br[191] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_192 bl[192] br[192] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_193 bl[193] br[193] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_194 bl[194] br[194] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_195 bl[195] br[195] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_196 bl[196] br[196] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_197 bl[197] br[197] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_198 bl[198] br[198] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_199 bl[199] br[199] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_200 bl[200] br[200] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_201 bl[201] br[201] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_202 bl[202] br[202] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_203 bl[203] br[203] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_204 bl[204] br[204] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_205 bl[205] br[205] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_206 bl[206] br[206] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_207 bl[207] br[207] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_208 bl[208] br[208] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_209 bl[209] br[209] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_210 bl[210] br[210] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_211 bl[211] br[211] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_212 bl[212] br[212] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_213 bl[213] br[213] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_214 bl[214] br[214] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_215 bl[215] br[215] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_216 bl[216] br[216] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_217 bl[217] br[217] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_218 bl[218] br[218] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_219 bl[219] br[219] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_220 bl[220] br[220] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_221 bl[221] br[221] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_222 bl[222] br[222] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_223 bl[223] br[223] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_224 bl[224] br[224] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_225 bl[225] br[225] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_226 bl[226] br[226] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_227 bl[227] br[227] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_228 bl[228] br[228] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_229 bl[229] br[229] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_230 bl[230] br[230] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_231 bl[231] br[231] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_232 bl[232] br[232] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_233 bl[233] br[233] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_234 bl[234] br[234] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_235 bl[235] br[235] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_236 bl[236] br[236] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_237 bl[237] br[237] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_238 bl[238] br[238] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_239 bl[239] br[239] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_240 bl[240] br[240] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_241 bl[241] br[241] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_242 bl[242] br[242] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_243 bl[243] br[243] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_244 bl[244] br[244] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_245 bl[245] br[245] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_246 bl[246] br[246] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_247 bl[247] br[247] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_248 bl[248] br[248] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_249 bl[249] br[249] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_250 bl[250] br[250] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_251 bl[251] br[251] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_252 bl[252] br[252] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_253 bl[253] br[253] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_254 bl[254] br[254] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_255 bl[255] br[255] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_46_0 bl[0] br[0] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_1 bl[1] br[1] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_2 bl[2] br[2] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_3 bl[3] br[3] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_4 bl[4] br[4] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_5 bl[5] br[5] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_6 bl[6] br[6] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_7 bl[7] br[7] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_8 bl[8] br[8] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_9 bl[9] br[9] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_10 bl[10] br[10] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_11 bl[11] br[11] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_12 bl[12] br[12] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_13 bl[13] br[13] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_14 bl[14] br[14] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_15 bl[15] br[15] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_16 bl[16] br[16] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_17 bl[17] br[17] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_18 bl[18] br[18] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_19 bl[19] br[19] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_20 bl[20] br[20] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_21 bl[21] br[21] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_22 bl[22] br[22] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_23 bl[23] br[23] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_24 bl[24] br[24] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_25 bl[25] br[25] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_26 bl[26] br[26] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_27 bl[27] br[27] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_28 bl[28] br[28] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_29 bl[29] br[29] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_30 bl[30] br[30] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_31 bl[31] br[31] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_32 bl[32] br[32] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_33 bl[33] br[33] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_34 bl[34] br[34] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_35 bl[35] br[35] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_36 bl[36] br[36] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_37 bl[37] br[37] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_38 bl[38] br[38] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_39 bl[39] br[39] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_40 bl[40] br[40] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_41 bl[41] br[41] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_42 bl[42] br[42] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_43 bl[43] br[43] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_44 bl[44] br[44] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_45 bl[45] br[45] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_46 bl[46] br[46] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_47 bl[47] br[47] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_48 bl[48] br[48] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_49 bl[49] br[49] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_50 bl[50] br[50] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_51 bl[51] br[51] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_52 bl[52] br[52] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_53 bl[53] br[53] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_54 bl[54] br[54] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_55 bl[55] br[55] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_56 bl[56] br[56] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_57 bl[57] br[57] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_58 bl[58] br[58] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_59 bl[59] br[59] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_60 bl[60] br[60] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_61 bl[61] br[61] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_62 bl[62] br[62] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_63 bl[63] br[63] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_64 bl[64] br[64] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_65 bl[65] br[65] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_66 bl[66] br[66] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_67 bl[67] br[67] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_68 bl[68] br[68] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_69 bl[69] br[69] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_70 bl[70] br[70] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_71 bl[71] br[71] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_72 bl[72] br[72] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_73 bl[73] br[73] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_74 bl[74] br[74] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_75 bl[75] br[75] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_76 bl[76] br[76] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_77 bl[77] br[77] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_78 bl[78] br[78] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_79 bl[79] br[79] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_80 bl[80] br[80] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_81 bl[81] br[81] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_82 bl[82] br[82] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_83 bl[83] br[83] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_84 bl[84] br[84] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_85 bl[85] br[85] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_86 bl[86] br[86] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_87 bl[87] br[87] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_88 bl[88] br[88] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_89 bl[89] br[89] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_90 bl[90] br[90] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_91 bl[91] br[91] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_92 bl[92] br[92] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_93 bl[93] br[93] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_94 bl[94] br[94] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_95 bl[95] br[95] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_96 bl[96] br[96] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_97 bl[97] br[97] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_98 bl[98] br[98] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_99 bl[99] br[99] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_100 bl[100] br[100] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_101 bl[101] br[101] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_102 bl[102] br[102] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_103 bl[103] br[103] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_104 bl[104] br[104] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_105 bl[105] br[105] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_106 bl[106] br[106] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_107 bl[107] br[107] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_108 bl[108] br[108] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_109 bl[109] br[109] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_110 bl[110] br[110] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_111 bl[111] br[111] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_112 bl[112] br[112] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_113 bl[113] br[113] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_114 bl[114] br[114] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_115 bl[115] br[115] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_116 bl[116] br[116] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_117 bl[117] br[117] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_118 bl[118] br[118] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_119 bl[119] br[119] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_120 bl[120] br[120] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_121 bl[121] br[121] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_122 bl[122] br[122] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_123 bl[123] br[123] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_124 bl[124] br[124] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_125 bl[125] br[125] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_126 bl[126] br[126] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_127 bl[127] br[127] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_128 bl[128] br[128] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_129 bl[129] br[129] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_130 bl[130] br[130] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_131 bl[131] br[131] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_132 bl[132] br[132] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_133 bl[133] br[133] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_134 bl[134] br[134] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_135 bl[135] br[135] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_136 bl[136] br[136] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_137 bl[137] br[137] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_138 bl[138] br[138] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_139 bl[139] br[139] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_140 bl[140] br[140] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_141 bl[141] br[141] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_142 bl[142] br[142] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_143 bl[143] br[143] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_144 bl[144] br[144] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_145 bl[145] br[145] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_146 bl[146] br[146] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_147 bl[147] br[147] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_148 bl[148] br[148] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_149 bl[149] br[149] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_150 bl[150] br[150] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_151 bl[151] br[151] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_152 bl[152] br[152] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_153 bl[153] br[153] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_154 bl[154] br[154] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_155 bl[155] br[155] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_156 bl[156] br[156] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_157 bl[157] br[157] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_158 bl[158] br[158] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_159 bl[159] br[159] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_160 bl[160] br[160] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_161 bl[161] br[161] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_162 bl[162] br[162] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_163 bl[163] br[163] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_164 bl[164] br[164] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_165 bl[165] br[165] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_166 bl[166] br[166] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_167 bl[167] br[167] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_168 bl[168] br[168] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_169 bl[169] br[169] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_170 bl[170] br[170] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_171 bl[171] br[171] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_172 bl[172] br[172] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_173 bl[173] br[173] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_174 bl[174] br[174] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_175 bl[175] br[175] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_176 bl[176] br[176] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_177 bl[177] br[177] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_178 bl[178] br[178] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_179 bl[179] br[179] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_180 bl[180] br[180] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_181 bl[181] br[181] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_182 bl[182] br[182] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_183 bl[183] br[183] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_184 bl[184] br[184] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_185 bl[185] br[185] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_186 bl[186] br[186] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_187 bl[187] br[187] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_188 bl[188] br[188] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_189 bl[189] br[189] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_190 bl[190] br[190] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_191 bl[191] br[191] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_192 bl[192] br[192] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_193 bl[193] br[193] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_194 bl[194] br[194] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_195 bl[195] br[195] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_196 bl[196] br[196] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_197 bl[197] br[197] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_198 bl[198] br[198] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_199 bl[199] br[199] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_200 bl[200] br[200] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_201 bl[201] br[201] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_202 bl[202] br[202] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_203 bl[203] br[203] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_204 bl[204] br[204] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_205 bl[205] br[205] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_206 bl[206] br[206] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_207 bl[207] br[207] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_208 bl[208] br[208] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_209 bl[209] br[209] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_210 bl[210] br[210] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_211 bl[211] br[211] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_212 bl[212] br[212] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_213 bl[213] br[213] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_214 bl[214] br[214] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_215 bl[215] br[215] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_216 bl[216] br[216] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_217 bl[217] br[217] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_218 bl[218] br[218] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_219 bl[219] br[219] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_220 bl[220] br[220] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_221 bl[221] br[221] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_222 bl[222] br[222] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_223 bl[223] br[223] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_224 bl[224] br[224] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_225 bl[225] br[225] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_226 bl[226] br[226] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_227 bl[227] br[227] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_228 bl[228] br[228] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_229 bl[229] br[229] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_230 bl[230] br[230] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_231 bl[231] br[231] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_232 bl[232] br[232] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_233 bl[233] br[233] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_234 bl[234] br[234] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_235 bl[235] br[235] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_236 bl[236] br[236] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_237 bl[237] br[237] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_238 bl[238] br[238] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_239 bl[239] br[239] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_240 bl[240] br[240] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_241 bl[241] br[241] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_242 bl[242] br[242] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_243 bl[243] br[243] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_244 bl[244] br[244] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_245 bl[245] br[245] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_246 bl[246] br[246] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_247 bl[247] br[247] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_248 bl[248] br[248] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_249 bl[249] br[249] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_250 bl[250] br[250] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_251 bl[251] br[251] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_252 bl[252] br[252] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_253 bl[253] br[253] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_254 bl[254] br[254] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_255 bl[255] br[255] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_47_0 bl[0] br[0] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_1 bl[1] br[1] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_2 bl[2] br[2] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_3 bl[3] br[3] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_4 bl[4] br[4] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_5 bl[5] br[5] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_6 bl[6] br[6] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_7 bl[7] br[7] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_8 bl[8] br[8] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_9 bl[9] br[9] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_10 bl[10] br[10] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_11 bl[11] br[11] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_12 bl[12] br[12] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_13 bl[13] br[13] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_14 bl[14] br[14] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_15 bl[15] br[15] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_16 bl[16] br[16] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_17 bl[17] br[17] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_18 bl[18] br[18] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_19 bl[19] br[19] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_20 bl[20] br[20] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_21 bl[21] br[21] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_22 bl[22] br[22] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_23 bl[23] br[23] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_24 bl[24] br[24] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_25 bl[25] br[25] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_26 bl[26] br[26] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_27 bl[27] br[27] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_28 bl[28] br[28] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_29 bl[29] br[29] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_30 bl[30] br[30] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_31 bl[31] br[31] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_32 bl[32] br[32] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_33 bl[33] br[33] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_34 bl[34] br[34] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_35 bl[35] br[35] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_36 bl[36] br[36] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_37 bl[37] br[37] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_38 bl[38] br[38] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_39 bl[39] br[39] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_40 bl[40] br[40] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_41 bl[41] br[41] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_42 bl[42] br[42] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_43 bl[43] br[43] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_44 bl[44] br[44] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_45 bl[45] br[45] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_46 bl[46] br[46] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_47 bl[47] br[47] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_48 bl[48] br[48] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_49 bl[49] br[49] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_50 bl[50] br[50] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_51 bl[51] br[51] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_52 bl[52] br[52] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_53 bl[53] br[53] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_54 bl[54] br[54] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_55 bl[55] br[55] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_56 bl[56] br[56] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_57 bl[57] br[57] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_58 bl[58] br[58] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_59 bl[59] br[59] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_60 bl[60] br[60] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_61 bl[61] br[61] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_62 bl[62] br[62] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_63 bl[63] br[63] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_64 bl[64] br[64] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_65 bl[65] br[65] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_66 bl[66] br[66] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_67 bl[67] br[67] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_68 bl[68] br[68] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_69 bl[69] br[69] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_70 bl[70] br[70] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_71 bl[71] br[71] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_72 bl[72] br[72] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_73 bl[73] br[73] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_74 bl[74] br[74] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_75 bl[75] br[75] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_76 bl[76] br[76] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_77 bl[77] br[77] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_78 bl[78] br[78] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_79 bl[79] br[79] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_80 bl[80] br[80] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_81 bl[81] br[81] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_82 bl[82] br[82] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_83 bl[83] br[83] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_84 bl[84] br[84] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_85 bl[85] br[85] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_86 bl[86] br[86] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_87 bl[87] br[87] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_88 bl[88] br[88] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_89 bl[89] br[89] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_90 bl[90] br[90] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_91 bl[91] br[91] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_92 bl[92] br[92] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_93 bl[93] br[93] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_94 bl[94] br[94] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_95 bl[95] br[95] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_96 bl[96] br[96] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_97 bl[97] br[97] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_98 bl[98] br[98] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_99 bl[99] br[99] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_100 bl[100] br[100] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_101 bl[101] br[101] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_102 bl[102] br[102] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_103 bl[103] br[103] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_104 bl[104] br[104] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_105 bl[105] br[105] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_106 bl[106] br[106] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_107 bl[107] br[107] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_108 bl[108] br[108] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_109 bl[109] br[109] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_110 bl[110] br[110] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_111 bl[111] br[111] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_112 bl[112] br[112] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_113 bl[113] br[113] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_114 bl[114] br[114] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_115 bl[115] br[115] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_116 bl[116] br[116] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_117 bl[117] br[117] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_118 bl[118] br[118] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_119 bl[119] br[119] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_120 bl[120] br[120] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_121 bl[121] br[121] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_122 bl[122] br[122] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_123 bl[123] br[123] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_124 bl[124] br[124] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_125 bl[125] br[125] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_126 bl[126] br[126] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_127 bl[127] br[127] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_128 bl[128] br[128] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_129 bl[129] br[129] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_130 bl[130] br[130] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_131 bl[131] br[131] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_132 bl[132] br[132] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_133 bl[133] br[133] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_134 bl[134] br[134] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_135 bl[135] br[135] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_136 bl[136] br[136] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_137 bl[137] br[137] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_138 bl[138] br[138] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_139 bl[139] br[139] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_140 bl[140] br[140] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_141 bl[141] br[141] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_142 bl[142] br[142] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_143 bl[143] br[143] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_144 bl[144] br[144] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_145 bl[145] br[145] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_146 bl[146] br[146] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_147 bl[147] br[147] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_148 bl[148] br[148] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_149 bl[149] br[149] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_150 bl[150] br[150] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_151 bl[151] br[151] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_152 bl[152] br[152] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_153 bl[153] br[153] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_154 bl[154] br[154] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_155 bl[155] br[155] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_156 bl[156] br[156] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_157 bl[157] br[157] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_158 bl[158] br[158] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_159 bl[159] br[159] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_160 bl[160] br[160] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_161 bl[161] br[161] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_162 bl[162] br[162] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_163 bl[163] br[163] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_164 bl[164] br[164] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_165 bl[165] br[165] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_166 bl[166] br[166] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_167 bl[167] br[167] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_168 bl[168] br[168] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_169 bl[169] br[169] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_170 bl[170] br[170] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_171 bl[171] br[171] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_172 bl[172] br[172] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_173 bl[173] br[173] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_174 bl[174] br[174] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_175 bl[175] br[175] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_176 bl[176] br[176] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_177 bl[177] br[177] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_178 bl[178] br[178] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_179 bl[179] br[179] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_180 bl[180] br[180] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_181 bl[181] br[181] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_182 bl[182] br[182] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_183 bl[183] br[183] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_184 bl[184] br[184] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_185 bl[185] br[185] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_186 bl[186] br[186] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_187 bl[187] br[187] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_188 bl[188] br[188] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_189 bl[189] br[189] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_190 bl[190] br[190] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_191 bl[191] br[191] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_192 bl[192] br[192] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_193 bl[193] br[193] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_194 bl[194] br[194] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_195 bl[195] br[195] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_196 bl[196] br[196] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_197 bl[197] br[197] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_198 bl[198] br[198] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_199 bl[199] br[199] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_200 bl[200] br[200] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_201 bl[201] br[201] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_202 bl[202] br[202] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_203 bl[203] br[203] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_204 bl[204] br[204] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_205 bl[205] br[205] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_206 bl[206] br[206] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_207 bl[207] br[207] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_208 bl[208] br[208] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_209 bl[209] br[209] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_210 bl[210] br[210] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_211 bl[211] br[211] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_212 bl[212] br[212] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_213 bl[213] br[213] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_214 bl[214] br[214] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_215 bl[215] br[215] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_216 bl[216] br[216] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_217 bl[217] br[217] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_218 bl[218] br[218] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_219 bl[219] br[219] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_220 bl[220] br[220] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_221 bl[221] br[221] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_222 bl[222] br[222] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_223 bl[223] br[223] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_224 bl[224] br[224] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_225 bl[225] br[225] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_226 bl[226] br[226] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_227 bl[227] br[227] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_228 bl[228] br[228] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_229 bl[229] br[229] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_230 bl[230] br[230] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_231 bl[231] br[231] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_232 bl[232] br[232] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_233 bl[233] br[233] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_234 bl[234] br[234] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_235 bl[235] br[235] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_236 bl[236] br[236] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_237 bl[237] br[237] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_238 bl[238] br[238] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_239 bl[239] br[239] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_240 bl[240] br[240] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_241 bl[241] br[241] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_242 bl[242] br[242] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_243 bl[243] br[243] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_244 bl[244] br[244] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_245 bl[245] br[245] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_246 bl[246] br[246] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_247 bl[247] br[247] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_248 bl[248] br[248] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_249 bl[249] br[249] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_250 bl[250] br[250] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_251 bl[251] br[251] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_252 bl[252] br[252] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_253 bl[253] br[253] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_254 bl[254] br[254] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_255 bl[255] br[255] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_48_0 bl[0] br[0] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_1 bl[1] br[1] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_2 bl[2] br[2] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_3 bl[3] br[3] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_4 bl[4] br[4] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_5 bl[5] br[5] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_6 bl[6] br[6] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_7 bl[7] br[7] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_8 bl[8] br[8] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_9 bl[9] br[9] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_10 bl[10] br[10] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_11 bl[11] br[11] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_12 bl[12] br[12] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_13 bl[13] br[13] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_14 bl[14] br[14] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_15 bl[15] br[15] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_16 bl[16] br[16] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_17 bl[17] br[17] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_18 bl[18] br[18] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_19 bl[19] br[19] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_20 bl[20] br[20] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_21 bl[21] br[21] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_22 bl[22] br[22] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_23 bl[23] br[23] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_24 bl[24] br[24] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_25 bl[25] br[25] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_26 bl[26] br[26] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_27 bl[27] br[27] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_28 bl[28] br[28] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_29 bl[29] br[29] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_30 bl[30] br[30] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_31 bl[31] br[31] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_32 bl[32] br[32] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_33 bl[33] br[33] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_34 bl[34] br[34] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_35 bl[35] br[35] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_36 bl[36] br[36] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_37 bl[37] br[37] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_38 bl[38] br[38] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_39 bl[39] br[39] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_40 bl[40] br[40] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_41 bl[41] br[41] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_42 bl[42] br[42] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_43 bl[43] br[43] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_44 bl[44] br[44] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_45 bl[45] br[45] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_46 bl[46] br[46] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_47 bl[47] br[47] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_48 bl[48] br[48] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_49 bl[49] br[49] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_50 bl[50] br[50] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_51 bl[51] br[51] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_52 bl[52] br[52] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_53 bl[53] br[53] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_54 bl[54] br[54] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_55 bl[55] br[55] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_56 bl[56] br[56] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_57 bl[57] br[57] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_58 bl[58] br[58] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_59 bl[59] br[59] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_60 bl[60] br[60] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_61 bl[61] br[61] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_62 bl[62] br[62] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_63 bl[63] br[63] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_64 bl[64] br[64] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_65 bl[65] br[65] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_66 bl[66] br[66] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_67 bl[67] br[67] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_68 bl[68] br[68] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_69 bl[69] br[69] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_70 bl[70] br[70] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_71 bl[71] br[71] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_72 bl[72] br[72] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_73 bl[73] br[73] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_74 bl[74] br[74] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_75 bl[75] br[75] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_76 bl[76] br[76] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_77 bl[77] br[77] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_78 bl[78] br[78] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_79 bl[79] br[79] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_80 bl[80] br[80] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_81 bl[81] br[81] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_82 bl[82] br[82] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_83 bl[83] br[83] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_84 bl[84] br[84] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_85 bl[85] br[85] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_86 bl[86] br[86] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_87 bl[87] br[87] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_88 bl[88] br[88] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_89 bl[89] br[89] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_90 bl[90] br[90] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_91 bl[91] br[91] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_92 bl[92] br[92] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_93 bl[93] br[93] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_94 bl[94] br[94] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_95 bl[95] br[95] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_96 bl[96] br[96] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_97 bl[97] br[97] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_98 bl[98] br[98] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_99 bl[99] br[99] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_100 bl[100] br[100] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_101 bl[101] br[101] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_102 bl[102] br[102] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_103 bl[103] br[103] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_104 bl[104] br[104] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_105 bl[105] br[105] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_106 bl[106] br[106] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_107 bl[107] br[107] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_108 bl[108] br[108] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_109 bl[109] br[109] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_110 bl[110] br[110] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_111 bl[111] br[111] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_112 bl[112] br[112] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_113 bl[113] br[113] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_114 bl[114] br[114] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_115 bl[115] br[115] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_116 bl[116] br[116] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_117 bl[117] br[117] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_118 bl[118] br[118] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_119 bl[119] br[119] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_120 bl[120] br[120] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_121 bl[121] br[121] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_122 bl[122] br[122] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_123 bl[123] br[123] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_124 bl[124] br[124] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_125 bl[125] br[125] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_126 bl[126] br[126] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_127 bl[127] br[127] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_128 bl[128] br[128] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_129 bl[129] br[129] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_130 bl[130] br[130] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_131 bl[131] br[131] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_132 bl[132] br[132] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_133 bl[133] br[133] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_134 bl[134] br[134] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_135 bl[135] br[135] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_136 bl[136] br[136] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_137 bl[137] br[137] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_138 bl[138] br[138] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_139 bl[139] br[139] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_140 bl[140] br[140] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_141 bl[141] br[141] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_142 bl[142] br[142] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_143 bl[143] br[143] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_144 bl[144] br[144] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_145 bl[145] br[145] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_146 bl[146] br[146] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_147 bl[147] br[147] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_148 bl[148] br[148] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_149 bl[149] br[149] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_150 bl[150] br[150] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_151 bl[151] br[151] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_152 bl[152] br[152] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_153 bl[153] br[153] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_154 bl[154] br[154] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_155 bl[155] br[155] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_156 bl[156] br[156] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_157 bl[157] br[157] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_158 bl[158] br[158] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_159 bl[159] br[159] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_160 bl[160] br[160] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_161 bl[161] br[161] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_162 bl[162] br[162] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_163 bl[163] br[163] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_164 bl[164] br[164] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_165 bl[165] br[165] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_166 bl[166] br[166] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_167 bl[167] br[167] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_168 bl[168] br[168] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_169 bl[169] br[169] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_170 bl[170] br[170] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_171 bl[171] br[171] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_172 bl[172] br[172] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_173 bl[173] br[173] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_174 bl[174] br[174] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_175 bl[175] br[175] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_176 bl[176] br[176] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_177 bl[177] br[177] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_178 bl[178] br[178] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_179 bl[179] br[179] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_180 bl[180] br[180] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_181 bl[181] br[181] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_182 bl[182] br[182] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_183 bl[183] br[183] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_184 bl[184] br[184] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_185 bl[185] br[185] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_186 bl[186] br[186] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_187 bl[187] br[187] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_188 bl[188] br[188] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_189 bl[189] br[189] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_190 bl[190] br[190] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_191 bl[191] br[191] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_192 bl[192] br[192] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_193 bl[193] br[193] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_194 bl[194] br[194] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_195 bl[195] br[195] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_196 bl[196] br[196] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_197 bl[197] br[197] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_198 bl[198] br[198] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_199 bl[199] br[199] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_200 bl[200] br[200] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_201 bl[201] br[201] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_202 bl[202] br[202] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_203 bl[203] br[203] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_204 bl[204] br[204] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_205 bl[205] br[205] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_206 bl[206] br[206] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_207 bl[207] br[207] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_208 bl[208] br[208] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_209 bl[209] br[209] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_210 bl[210] br[210] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_211 bl[211] br[211] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_212 bl[212] br[212] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_213 bl[213] br[213] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_214 bl[214] br[214] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_215 bl[215] br[215] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_216 bl[216] br[216] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_217 bl[217] br[217] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_218 bl[218] br[218] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_219 bl[219] br[219] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_220 bl[220] br[220] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_221 bl[221] br[221] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_222 bl[222] br[222] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_223 bl[223] br[223] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_224 bl[224] br[224] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_225 bl[225] br[225] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_226 bl[226] br[226] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_227 bl[227] br[227] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_228 bl[228] br[228] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_229 bl[229] br[229] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_230 bl[230] br[230] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_231 bl[231] br[231] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_232 bl[232] br[232] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_233 bl[233] br[233] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_234 bl[234] br[234] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_235 bl[235] br[235] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_236 bl[236] br[236] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_237 bl[237] br[237] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_238 bl[238] br[238] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_239 bl[239] br[239] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_240 bl[240] br[240] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_241 bl[241] br[241] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_242 bl[242] br[242] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_243 bl[243] br[243] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_244 bl[244] br[244] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_245 bl[245] br[245] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_246 bl[246] br[246] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_247 bl[247] br[247] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_248 bl[248] br[248] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_249 bl[249] br[249] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_250 bl[250] br[250] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_251 bl[251] br[251] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_252 bl[252] br[252] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_253 bl[253] br[253] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_254 bl[254] br[254] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_255 bl[255] br[255] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_49_0 bl[0] br[0] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_1 bl[1] br[1] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_2 bl[2] br[2] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_3 bl[3] br[3] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_4 bl[4] br[4] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_5 bl[5] br[5] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_6 bl[6] br[6] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_7 bl[7] br[7] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_8 bl[8] br[8] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_9 bl[9] br[9] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_10 bl[10] br[10] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_11 bl[11] br[11] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_12 bl[12] br[12] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_13 bl[13] br[13] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_14 bl[14] br[14] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_15 bl[15] br[15] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_16 bl[16] br[16] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_17 bl[17] br[17] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_18 bl[18] br[18] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_19 bl[19] br[19] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_20 bl[20] br[20] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_21 bl[21] br[21] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_22 bl[22] br[22] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_23 bl[23] br[23] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_24 bl[24] br[24] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_25 bl[25] br[25] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_26 bl[26] br[26] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_27 bl[27] br[27] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_28 bl[28] br[28] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_29 bl[29] br[29] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_30 bl[30] br[30] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_31 bl[31] br[31] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_32 bl[32] br[32] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_33 bl[33] br[33] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_34 bl[34] br[34] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_35 bl[35] br[35] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_36 bl[36] br[36] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_37 bl[37] br[37] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_38 bl[38] br[38] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_39 bl[39] br[39] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_40 bl[40] br[40] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_41 bl[41] br[41] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_42 bl[42] br[42] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_43 bl[43] br[43] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_44 bl[44] br[44] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_45 bl[45] br[45] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_46 bl[46] br[46] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_47 bl[47] br[47] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_48 bl[48] br[48] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_49 bl[49] br[49] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_50 bl[50] br[50] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_51 bl[51] br[51] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_52 bl[52] br[52] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_53 bl[53] br[53] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_54 bl[54] br[54] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_55 bl[55] br[55] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_56 bl[56] br[56] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_57 bl[57] br[57] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_58 bl[58] br[58] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_59 bl[59] br[59] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_60 bl[60] br[60] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_61 bl[61] br[61] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_62 bl[62] br[62] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_63 bl[63] br[63] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_64 bl[64] br[64] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_65 bl[65] br[65] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_66 bl[66] br[66] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_67 bl[67] br[67] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_68 bl[68] br[68] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_69 bl[69] br[69] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_70 bl[70] br[70] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_71 bl[71] br[71] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_72 bl[72] br[72] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_73 bl[73] br[73] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_74 bl[74] br[74] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_75 bl[75] br[75] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_76 bl[76] br[76] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_77 bl[77] br[77] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_78 bl[78] br[78] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_79 bl[79] br[79] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_80 bl[80] br[80] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_81 bl[81] br[81] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_82 bl[82] br[82] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_83 bl[83] br[83] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_84 bl[84] br[84] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_85 bl[85] br[85] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_86 bl[86] br[86] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_87 bl[87] br[87] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_88 bl[88] br[88] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_89 bl[89] br[89] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_90 bl[90] br[90] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_91 bl[91] br[91] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_92 bl[92] br[92] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_93 bl[93] br[93] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_94 bl[94] br[94] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_95 bl[95] br[95] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_96 bl[96] br[96] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_97 bl[97] br[97] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_98 bl[98] br[98] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_99 bl[99] br[99] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_100 bl[100] br[100] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_101 bl[101] br[101] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_102 bl[102] br[102] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_103 bl[103] br[103] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_104 bl[104] br[104] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_105 bl[105] br[105] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_106 bl[106] br[106] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_107 bl[107] br[107] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_108 bl[108] br[108] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_109 bl[109] br[109] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_110 bl[110] br[110] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_111 bl[111] br[111] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_112 bl[112] br[112] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_113 bl[113] br[113] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_114 bl[114] br[114] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_115 bl[115] br[115] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_116 bl[116] br[116] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_117 bl[117] br[117] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_118 bl[118] br[118] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_119 bl[119] br[119] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_120 bl[120] br[120] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_121 bl[121] br[121] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_122 bl[122] br[122] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_123 bl[123] br[123] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_124 bl[124] br[124] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_125 bl[125] br[125] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_126 bl[126] br[126] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_127 bl[127] br[127] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_128 bl[128] br[128] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_129 bl[129] br[129] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_130 bl[130] br[130] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_131 bl[131] br[131] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_132 bl[132] br[132] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_133 bl[133] br[133] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_134 bl[134] br[134] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_135 bl[135] br[135] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_136 bl[136] br[136] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_137 bl[137] br[137] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_138 bl[138] br[138] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_139 bl[139] br[139] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_140 bl[140] br[140] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_141 bl[141] br[141] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_142 bl[142] br[142] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_143 bl[143] br[143] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_144 bl[144] br[144] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_145 bl[145] br[145] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_146 bl[146] br[146] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_147 bl[147] br[147] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_148 bl[148] br[148] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_149 bl[149] br[149] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_150 bl[150] br[150] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_151 bl[151] br[151] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_152 bl[152] br[152] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_153 bl[153] br[153] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_154 bl[154] br[154] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_155 bl[155] br[155] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_156 bl[156] br[156] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_157 bl[157] br[157] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_158 bl[158] br[158] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_159 bl[159] br[159] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_160 bl[160] br[160] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_161 bl[161] br[161] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_162 bl[162] br[162] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_163 bl[163] br[163] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_164 bl[164] br[164] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_165 bl[165] br[165] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_166 bl[166] br[166] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_167 bl[167] br[167] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_168 bl[168] br[168] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_169 bl[169] br[169] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_170 bl[170] br[170] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_171 bl[171] br[171] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_172 bl[172] br[172] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_173 bl[173] br[173] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_174 bl[174] br[174] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_175 bl[175] br[175] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_176 bl[176] br[176] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_177 bl[177] br[177] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_178 bl[178] br[178] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_179 bl[179] br[179] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_180 bl[180] br[180] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_181 bl[181] br[181] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_182 bl[182] br[182] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_183 bl[183] br[183] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_184 bl[184] br[184] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_185 bl[185] br[185] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_186 bl[186] br[186] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_187 bl[187] br[187] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_188 bl[188] br[188] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_189 bl[189] br[189] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_190 bl[190] br[190] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_191 bl[191] br[191] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_192 bl[192] br[192] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_193 bl[193] br[193] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_194 bl[194] br[194] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_195 bl[195] br[195] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_196 bl[196] br[196] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_197 bl[197] br[197] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_198 bl[198] br[198] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_199 bl[199] br[199] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_200 bl[200] br[200] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_201 bl[201] br[201] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_202 bl[202] br[202] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_203 bl[203] br[203] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_204 bl[204] br[204] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_205 bl[205] br[205] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_206 bl[206] br[206] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_207 bl[207] br[207] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_208 bl[208] br[208] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_209 bl[209] br[209] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_210 bl[210] br[210] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_211 bl[211] br[211] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_212 bl[212] br[212] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_213 bl[213] br[213] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_214 bl[214] br[214] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_215 bl[215] br[215] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_216 bl[216] br[216] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_217 bl[217] br[217] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_218 bl[218] br[218] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_219 bl[219] br[219] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_220 bl[220] br[220] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_221 bl[221] br[221] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_222 bl[222] br[222] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_223 bl[223] br[223] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_224 bl[224] br[224] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_225 bl[225] br[225] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_226 bl[226] br[226] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_227 bl[227] br[227] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_228 bl[228] br[228] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_229 bl[229] br[229] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_230 bl[230] br[230] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_231 bl[231] br[231] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_232 bl[232] br[232] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_233 bl[233] br[233] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_234 bl[234] br[234] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_235 bl[235] br[235] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_236 bl[236] br[236] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_237 bl[237] br[237] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_238 bl[238] br[238] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_239 bl[239] br[239] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_240 bl[240] br[240] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_241 bl[241] br[241] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_242 bl[242] br[242] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_243 bl[243] br[243] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_244 bl[244] br[244] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_245 bl[245] br[245] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_246 bl[246] br[246] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_247 bl[247] br[247] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_248 bl[248] br[248] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_249 bl[249] br[249] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_250 bl[250] br[250] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_251 bl[251] br[251] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_252 bl[252] br[252] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_253 bl[253] br[253] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_254 bl[254] br[254] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_255 bl[255] br[255] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_50_0 bl[0] br[0] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_1 bl[1] br[1] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_2 bl[2] br[2] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_3 bl[3] br[3] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_4 bl[4] br[4] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_5 bl[5] br[5] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_6 bl[6] br[6] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_7 bl[7] br[7] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_8 bl[8] br[8] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_9 bl[9] br[9] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_10 bl[10] br[10] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_11 bl[11] br[11] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_12 bl[12] br[12] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_13 bl[13] br[13] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_14 bl[14] br[14] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_15 bl[15] br[15] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_16 bl[16] br[16] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_17 bl[17] br[17] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_18 bl[18] br[18] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_19 bl[19] br[19] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_20 bl[20] br[20] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_21 bl[21] br[21] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_22 bl[22] br[22] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_23 bl[23] br[23] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_24 bl[24] br[24] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_25 bl[25] br[25] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_26 bl[26] br[26] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_27 bl[27] br[27] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_28 bl[28] br[28] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_29 bl[29] br[29] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_30 bl[30] br[30] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_31 bl[31] br[31] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_32 bl[32] br[32] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_33 bl[33] br[33] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_34 bl[34] br[34] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_35 bl[35] br[35] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_36 bl[36] br[36] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_37 bl[37] br[37] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_38 bl[38] br[38] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_39 bl[39] br[39] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_40 bl[40] br[40] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_41 bl[41] br[41] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_42 bl[42] br[42] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_43 bl[43] br[43] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_44 bl[44] br[44] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_45 bl[45] br[45] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_46 bl[46] br[46] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_47 bl[47] br[47] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_48 bl[48] br[48] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_49 bl[49] br[49] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_50 bl[50] br[50] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_51 bl[51] br[51] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_52 bl[52] br[52] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_53 bl[53] br[53] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_54 bl[54] br[54] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_55 bl[55] br[55] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_56 bl[56] br[56] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_57 bl[57] br[57] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_58 bl[58] br[58] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_59 bl[59] br[59] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_60 bl[60] br[60] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_61 bl[61] br[61] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_62 bl[62] br[62] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_63 bl[63] br[63] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_64 bl[64] br[64] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_65 bl[65] br[65] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_66 bl[66] br[66] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_67 bl[67] br[67] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_68 bl[68] br[68] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_69 bl[69] br[69] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_70 bl[70] br[70] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_71 bl[71] br[71] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_72 bl[72] br[72] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_73 bl[73] br[73] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_74 bl[74] br[74] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_75 bl[75] br[75] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_76 bl[76] br[76] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_77 bl[77] br[77] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_78 bl[78] br[78] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_79 bl[79] br[79] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_80 bl[80] br[80] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_81 bl[81] br[81] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_82 bl[82] br[82] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_83 bl[83] br[83] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_84 bl[84] br[84] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_85 bl[85] br[85] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_86 bl[86] br[86] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_87 bl[87] br[87] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_88 bl[88] br[88] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_89 bl[89] br[89] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_90 bl[90] br[90] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_91 bl[91] br[91] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_92 bl[92] br[92] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_93 bl[93] br[93] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_94 bl[94] br[94] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_95 bl[95] br[95] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_96 bl[96] br[96] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_97 bl[97] br[97] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_98 bl[98] br[98] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_99 bl[99] br[99] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_100 bl[100] br[100] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_101 bl[101] br[101] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_102 bl[102] br[102] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_103 bl[103] br[103] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_104 bl[104] br[104] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_105 bl[105] br[105] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_106 bl[106] br[106] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_107 bl[107] br[107] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_108 bl[108] br[108] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_109 bl[109] br[109] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_110 bl[110] br[110] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_111 bl[111] br[111] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_112 bl[112] br[112] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_113 bl[113] br[113] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_114 bl[114] br[114] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_115 bl[115] br[115] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_116 bl[116] br[116] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_117 bl[117] br[117] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_118 bl[118] br[118] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_119 bl[119] br[119] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_120 bl[120] br[120] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_121 bl[121] br[121] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_122 bl[122] br[122] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_123 bl[123] br[123] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_124 bl[124] br[124] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_125 bl[125] br[125] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_126 bl[126] br[126] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_127 bl[127] br[127] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_128 bl[128] br[128] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_129 bl[129] br[129] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_130 bl[130] br[130] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_131 bl[131] br[131] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_132 bl[132] br[132] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_133 bl[133] br[133] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_134 bl[134] br[134] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_135 bl[135] br[135] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_136 bl[136] br[136] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_137 bl[137] br[137] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_138 bl[138] br[138] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_139 bl[139] br[139] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_140 bl[140] br[140] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_141 bl[141] br[141] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_142 bl[142] br[142] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_143 bl[143] br[143] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_144 bl[144] br[144] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_145 bl[145] br[145] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_146 bl[146] br[146] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_147 bl[147] br[147] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_148 bl[148] br[148] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_149 bl[149] br[149] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_150 bl[150] br[150] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_151 bl[151] br[151] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_152 bl[152] br[152] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_153 bl[153] br[153] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_154 bl[154] br[154] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_155 bl[155] br[155] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_156 bl[156] br[156] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_157 bl[157] br[157] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_158 bl[158] br[158] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_159 bl[159] br[159] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_160 bl[160] br[160] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_161 bl[161] br[161] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_162 bl[162] br[162] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_163 bl[163] br[163] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_164 bl[164] br[164] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_165 bl[165] br[165] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_166 bl[166] br[166] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_167 bl[167] br[167] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_168 bl[168] br[168] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_169 bl[169] br[169] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_170 bl[170] br[170] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_171 bl[171] br[171] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_172 bl[172] br[172] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_173 bl[173] br[173] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_174 bl[174] br[174] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_175 bl[175] br[175] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_176 bl[176] br[176] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_177 bl[177] br[177] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_178 bl[178] br[178] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_179 bl[179] br[179] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_180 bl[180] br[180] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_181 bl[181] br[181] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_182 bl[182] br[182] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_183 bl[183] br[183] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_184 bl[184] br[184] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_185 bl[185] br[185] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_186 bl[186] br[186] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_187 bl[187] br[187] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_188 bl[188] br[188] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_189 bl[189] br[189] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_190 bl[190] br[190] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_191 bl[191] br[191] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_192 bl[192] br[192] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_193 bl[193] br[193] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_194 bl[194] br[194] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_195 bl[195] br[195] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_196 bl[196] br[196] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_197 bl[197] br[197] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_198 bl[198] br[198] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_199 bl[199] br[199] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_200 bl[200] br[200] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_201 bl[201] br[201] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_202 bl[202] br[202] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_203 bl[203] br[203] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_204 bl[204] br[204] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_205 bl[205] br[205] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_206 bl[206] br[206] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_207 bl[207] br[207] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_208 bl[208] br[208] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_209 bl[209] br[209] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_210 bl[210] br[210] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_211 bl[211] br[211] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_212 bl[212] br[212] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_213 bl[213] br[213] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_214 bl[214] br[214] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_215 bl[215] br[215] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_216 bl[216] br[216] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_217 bl[217] br[217] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_218 bl[218] br[218] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_219 bl[219] br[219] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_220 bl[220] br[220] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_221 bl[221] br[221] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_222 bl[222] br[222] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_223 bl[223] br[223] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_224 bl[224] br[224] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_225 bl[225] br[225] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_226 bl[226] br[226] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_227 bl[227] br[227] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_228 bl[228] br[228] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_229 bl[229] br[229] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_230 bl[230] br[230] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_231 bl[231] br[231] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_232 bl[232] br[232] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_233 bl[233] br[233] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_234 bl[234] br[234] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_235 bl[235] br[235] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_236 bl[236] br[236] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_237 bl[237] br[237] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_238 bl[238] br[238] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_239 bl[239] br[239] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_240 bl[240] br[240] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_241 bl[241] br[241] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_242 bl[242] br[242] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_243 bl[243] br[243] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_244 bl[244] br[244] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_245 bl[245] br[245] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_246 bl[246] br[246] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_247 bl[247] br[247] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_248 bl[248] br[248] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_249 bl[249] br[249] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_250 bl[250] br[250] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_251 bl[251] br[251] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_252 bl[252] br[252] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_253 bl[253] br[253] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_254 bl[254] br[254] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_255 bl[255] br[255] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_51_0 bl[0] br[0] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_1 bl[1] br[1] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_2 bl[2] br[2] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_3 bl[3] br[3] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_4 bl[4] br[4] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_5 bl[5] br[5] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_6 bl[6] br[6] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_7 bl[7] br[7] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_8 bl[8] br[8] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_9 bl[9] br[9] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_10 bl[10] br[10] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_11 bl[11] br[11] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_12 bl[12] br[12] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_13 bl[13] br[13] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_14 bl[14] br[14] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_15 bl[15] br[15] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_16 bl[16] br[16] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_17 bl[17] br[17] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_18 bl[18] br[18] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_19 bl[19] br[19] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_20 bl[20] br[20] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_21 bl[21] br[21] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_22 bl[22] br[22] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_23 bl[23] br[23] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_24 bl[24] br[24] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_25 bl[25] br[25] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_26 bl[26] br[26] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_27 bl[27] br[27] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_28 bl[28] br[28] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_29 bl[29] br[29] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_30 bl[30] br[30] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_31 bl[31] br[31] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_32 bl[32] br[32] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_33 bl[33] br[33] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_34 bl[34] br[34] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_35 bl[35] br[35] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_36 bl[36] br[36] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_37 bl[37] br[37] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_38 bl[38] br[38] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_39 bl[39] br[39] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_40 bl[40] br[40] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_41 bl[41] br[41] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_42 bl[42] br[42] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_43 bl[43] br[43] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_44 bl[44] br[44] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_45 bl[45] br[45] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_46 bl[46] br[46] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_47 bl[47] br[47] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_48 bl[48] br[48] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_49 bl[49] br[49] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_50 bl[50] br[50] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_51 bl[51] br[51] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_52 bl[52] br[52] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_53 bl[53] br[53] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_54 bl[54] br[54] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_55 bl[55] br[55] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_56 bl[56] br[56] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_57 bl[57] br[57] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_58 bl[58] br[58] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_59 bl[59] br[59] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_60 bl[60] br[60] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_61 bl[61] br[61] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_62 bl[62] br[62] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_63 bl[63] br[63] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_64 bl[64] br[64] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_65 bl[65] br[65] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_66 bl[66] br[66] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_67 bl[67] br[67] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_68 bl[68] br[68] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_69 bl[69] br[69] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_70 bl[70] br[70] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_71 bl[71] br[71] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_72 bl[72] br[72] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_73 bl[73] br[73] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_74 bl[74] br[74] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_75 bl[75] br[75] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_76 bl[76] br[76] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_77 bl[77] br[77] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_78 bl[78] br[78] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_79 bl[79] br[79] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_80 bl[80] br[80] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_81 bl[81] br[81] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_82 bl[82] br[82] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_83 bl[83] br[83] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_84 bl[84] br[84] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_85 bl[85] br[85] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_86 bl[86] br[86] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_87 bl[87] br[87] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_88 bl[88] br[88] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_89 bl[89] br[89] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_90 bl[90] br[90] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_91 bl[91] br[91] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_92 bl[92] br[92] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_93 bl[93] br[93] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_94 bl[94] br[94] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_95 bl[95] br[95] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_96 bl[96] br[96] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_97 bl[97] br[97] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_98 bl[98] br[98] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_99 bl[99] br[99] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_100 bl[100] br[100] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_101 bl[101] br[101] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_102 bl[102] br[102] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_103 bl[103] br[103] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_104 bl[104] br[104] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_105 bl[105] br[105] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_106 bl[106] br[106] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_107 bl[107] br[107] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_108 bl[108] br[108] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_109 bl[109] br[109] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_110 bl[110] br[110] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_111 bl[111] br[111] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_112 bl[112] br[112] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_113 bl[113] br[113] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_114 bl[114] br[114] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_115 bl[115] br[115] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_116 bl[116] br[116] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_117 bl[117] br[117] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_118 bl[118] br[118] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_119 bl[119] br[119] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_120 bl[120] br[120] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_121 bl[121] br[121] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_122 bl[122] br[122] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_123 bl[123] br[123] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_124 bl[124] br[124] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_125 bl[125] br[125] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_126 bl[126] br[126] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_127 bl[127] br[127] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_128 bl[128] br[128] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_129 bl[129] br[129] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_130 bl[130] br[130] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_131 bl[131] br[131] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_132 bl[132] br[132] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_133 bl[133] br[133] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_134 bl[134] br[134] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_135 bl[135] br[135] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_136 bl[136] br[136] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_137 bl[137] br[137] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_138 bl[138] br[138] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_139 bl[139] br[139] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_140 bl[140] br[140] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_141 bl[141] br[141] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_142 bl[142] br[142] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_143 bl[143] br[143] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_144 bl[144] br[144] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_145 bl[145] br[145] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_146 bl[146] br[146] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_147 bl[147] br[147] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_148 bl[148] br[148] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_149 bl[149] br[149] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_150 bl[150] br[150] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_151 bl[151] br[151] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_152 bl[152] br[152] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_153 bl[153] br[153] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_154 bl[154] br[154] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_155 bl[155] br[155] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_156 bl[156] br[156] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_157 bl[157] br[157] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_158 bl[158] br[158] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_159 bl[159] br[159] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_160 bl[160] br[160] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_161 bl[161] br[161] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_162 bl[162] br[162] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_163 bl[163] br[163] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_164 bl[164] br[164] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_165 bl[165] br[165] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_166 bl[166] br[166] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_167 bl[167] br[167] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_168 bl[168] br[168] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_169 bl[169] br[169] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_170 bl[170] br[170] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_171 bl[171] br[171] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_172 bl[172] br[172] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_173 bl[173] br[173] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_174 bl[174] br[174] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_175 bl[175] br[175] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_176 bl[176] br[176] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_177 bl[177] br[177] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_178 bl[178] br[178] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_179 bl[179] br[179] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_180 bl[180] br[180] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_181 bl[181] br[181] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_182 bl[182] br[182] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_183 bl[183] br[183] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_184 bl[184] br[184] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_185 bl[185] br[185] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_186 bl[186] br[186] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_187 bl[187] br[187] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_188 bl[188] br[188] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_189 bl[189] br[189] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_190 bl[190] br[190] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_191 bl[191] br[191] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_192 bl[192] br[192] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_193 bl[193] br[193] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_194 bl[194] br[194] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_195 bl[195] br[195] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_196 bl[196] br[196] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_197 bl[197] br[197] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_198 bl[198] br[198] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_199 bl[199] br[199] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_200 bl[200] br[200] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_201 bl[201] br[201] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_202 bl[202] br[202] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_203 bl[203] br[203] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_204 bl[204] br[204] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_205 bl[205] br[205] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_206 bl[206] br[206] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_207 bl[207] br[207] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_208 bl[208] br[208] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_209 bl[209] br[209] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_210 bl[210] br[210] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_211 bl[211] br[211] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_212 bl[212] br[212] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_213 bl[213] br[213] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_214 bl[214] br[214] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_215 bl[215] br[215] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_216 bl[216] br[216] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_217 bl[217] br[217] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_218 bl[218] br[218] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_219 bl[219] br[219] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_220 bl[220] br[220] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_221 bl[221] br[221] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_222 bl[222] br[222] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_223 bl[223] br[223] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_224 bl[224] br[224] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_225 bl[225] br[225] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_226 bl[226] br[226] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_227 bl[227] br[227] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_228 bl[228] br[228] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_229 bl[229] br[229] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_230 bl[230] br[230] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_231 bl[231] br[231] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_232 bl[232] br[232] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_233 bl[233] br[233] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_234 bl[234] br[234] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_235 bl[235] br[235] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_236 bl[236] br[236] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_237 bl[237] br[237] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_238 bl[238] br[238] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_239 bl[239] br[239] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_240 bl[240] br[240] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_241 bl[241] br[241] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_242 bl[242] br[242] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_243 bl[243] br[243] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_244 bl[244] br[244] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_245 bl[245] br[245] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_246 bl[246] br[246] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_247 bl[247] br[247] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_248 bl[248] br[248] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_249 bl[249] br[249] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_250 bl[250] br[250] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_251 bl[251] br[251] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_252 bl[252] br[252] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_253 bl[253] br[253] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_254 bl[254] br[254] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_255 bl[255] br[255] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_52_0 bl[0] br[0] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_1 bl[1] br[1] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_2 bl[2] br[2] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_3 bl[3] br[3] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_4 bl[4] br[4] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_5 bl[5] br[5] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_6 bl[6] br[6] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_7 bl[7] br[7] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_8 bl[8] br[8] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_9 bl[9] br[9] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_10 bl[10] br[10] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_11 bl[11] br[11] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_12 bl[12] br[12] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_13 bl[13] br[13] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_14 bl[14] br[14] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_15 bl[15] br[15] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_16 bl[16] br[16] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_17 bl[17] br[17] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_18 bl[18] br[18] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_19 bl[19] br[19] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_20 bl[20] br[20] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_21 bl[21] br[21] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_22 bl[22] br[22] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_23 bl[23] br[23] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_24 bl[24] br[24] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_25 bl[25] br[25] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_26 bl[26] br[26] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_27 bl[27] br[27] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_28 bl[28] br[28] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_29 bl[29] br[29] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_30 bl[30] br[30] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_31 bl[31] br[31] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_32 bl[32] br[32] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_33 bl[33] br[33] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_34 bl[34] br[34] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_35 bl[35] br[35] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_36 bl[36] br[36] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_37 bl[37] br[37] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_38 bl[38] br[38] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_39 bl[39] br[39] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_40 bl[40] br[40] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_41 bl[41] br[41] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_42 bl[42] br[42] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_43 bl[43] br[43] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_44 bl[44] br[44] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_45 bl[45] br[45] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_46 bl[46] br[46] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_47 bl[47] br[47] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_48 bl[48] br[48] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_49 bl[49] br[49] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_50 bl[50] br[50] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_51 bl[51] br[51] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_52 bl[52] br[52] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_53 bl[53] br[53] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_54 bl[54] br[54] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_55 bl[55] br[55] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_56 bl[56] br[56] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_57 bl[57] br[57] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_58 bl[58] br[58] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_59 bl[59] br[59] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_60 bl[60] br[60] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_61 bl[61] br[61] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_62 bl[62] br[62] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_63 bl[63] br[63] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_64 bl[64] br[64] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_65 bl[65] br[65] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_66 bl[66] br[66] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_67 bl[67] br[67] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_68 bl[68] br[68] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_69 bl[69] br[69] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_70 bl[70] br[70] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_71 bl[71] br[71] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_72 bl[72] br[72] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_73 bl[73] br[73] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_74 bl[74] br[74] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_75 bl[75] br[75] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_76 bl[76] br[76] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_77 bl[77] br[77] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_78 bl[78] br[78] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_79 bl[79] br[79] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_80 bl[80] br[80] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_81 bl[81] br[81] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_82 bl[82] br[82] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_83 bl[83] br[83] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_84 bl[84] br[84] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_85 bl[85] br[85] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_86 bl[86] br[86] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_87 bl[87] br[87] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_88 bl[88] br[88] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_89 bl[89] br[89] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_90 bl[90] br[90] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_91 bl[91] br[91] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_92 bl[92] br[92] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_93 bl[93] br[93] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_94 bl[94] br[94] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_95 bl[95] br[95] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_96 bl[96] br[96] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_97 bl[97] br[97] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_98 bl[98] br[98] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_99 bl[99] br[99] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_100 bl[100] br[100] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_101 bl[101] br[101] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_102 bl[102] br[102] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_103 bl[103] br[103] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_104 bl[104] br[104] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_105 bl[105] br[105] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_106 bl[106] br[106] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_107 bl[107] br[107] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_108 bl[108] br[108] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_109 bl[109] br[109] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_110 bl[110] br[110] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_111 bl[111] br[111] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_112 bl[112] br[112] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_113 bl[113] br[113] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_114 bl[114] br[114] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_115 bl[115] br[115] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_116 bl[116] br[116] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_117 bl[117] br[117] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_118 bl[118] br[118] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_119 bl[119] br[119] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_120 bl[120] br[120] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_121 bl[121] br[121] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_122 bl[122] br[122] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_123 bl[123] br[123] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_124 bl[124] br[124] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_125 bl[125] br[125] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_126 bl[126] br[126] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_127 bl[127] br[127] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_128 bl[128] br[128] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_129 bl[129] br[129] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_130 bl[130] br[130] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_131 bl[131] br[131] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_132 bl[132] br[132] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_133 bl[133] br[133] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_134 bl[134] br[134] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_135 bl[135] br[135] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_136 bl[136] br[136] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_137 bl[137] br[137] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_138 bl[138] br[138] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_139 bl[139] br[139] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_140 bl[140] br[140] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_141 bl[141] br[141] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_142 bl[142] br[142] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_143 bl[143] br[143] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_144 bl[144] br[144] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_145 bl[145] br[145] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_146 bl[146] br[146] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_147 bl[147] br[147] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_148 bl[148] br[148] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_149 bl[149] br[149] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_150 bl[150] br[150] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_151 bl[151] br[151] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_152 bl[152] br[152] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_153 bl[153] br[153] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_154 bl[154] br[154] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_155 bl[155] br[155] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_156 bl[156] br[156] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_157 bl[157] br[157] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_158 bl[158] br[158] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_159 bl[159] br[159] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_160 bl[160] br[160] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_161 bl[161] br[161] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_162 bl[162] br[162] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_163 bl[163] br[163] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_164 bl[164] br[164] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_165 bl[165] br[165] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_166 bl[166] br[166] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_167 bl[167] br[167] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_168 bl[168] br[168] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_169 bl[169] br[169] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_170 bl[170] br[170] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_171 bl[171] br[171] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_172 bl[172] br[172] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_173 bl[173] br[173] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_174 bl[174] br[174] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_175 bl[175] br[175] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_176 bl[176] br[176] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_177 bl[177] br[177] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_178 bl[178] br[178] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_179 bl[179] br[179] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_180 bl[180] br[180] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_181 bl[181] br[181] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_182 bl[182] br[182] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_183 bl[183] br[183] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_184 bl[184] br[184] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_185 bl[185] br[185] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_186 bl[186] br[186] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_187 bl[187] br[187] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_188 bl[188] br[188] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_189 bl[189] br[189] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_190 bl[190] br[190] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_191 bl[191] br[191] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_192 bl[192] br[192] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_193 bl[193] br[193] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_194 bl[194] br[194] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_195 bl[195] br[195] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_196 bl[196] br[196] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_197 bl[197] br[197] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_198 bl[198] br[198] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_199 bl[199] br[199] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_200 bl[200] br[200] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_201 bl[201] br[201] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_202 bl[202] br[202] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_203 bl[203] br[203] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_204 bl[204] br[204] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_205 bl[205] br[205] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_206 bl[206] br[206] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_207 bl[207] br[207] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_208 bl[208] br[208] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_209 bl[209] br[209] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_210 bl[210] br[210] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_211 bl[211] br[211] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_212 bl[212] br[212] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_213 bl[213] br[213] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_214 bl[214] br[214] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_215 bl[215] br[215] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_216 bl[216] br[216] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_217 bl[217] br[217] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_218 bl[218] br[218] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_219 bl[219] br[219] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_220 bl[220] br[220] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_221 bl[221] br[221] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_222 bl[222] br[222] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_223 bl[223] br[223] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_224 bl[224] br[224] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_225 bl[225] br[225] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_226 bl[226] br[226] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_227 bl[227] br[227] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_228 bl[228] br[228] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_229 bl[229] br[229] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_230 bl[230] br[230] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_231 bl[231] br[231] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_232 bl[232] br[232] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_233 bl[233] br[233] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_234 bl[234] br[234] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_235 bl[235] br[235] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_236 bl[236] br[236] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_237 bl[237] br[237] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_238 bl[238] br[238] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_239 bl[239] br[239] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_240 bl[240] br[240] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_241 bl[241] br[241] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_242 bl[242] br[242] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_243 bl[243] br[243] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_244 bl[244] br[244] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_245 bl[245] br[245] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_246 bl[246] br[246] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_247 bl[247] br[247] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_248 bl[248] br[248] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_249 bl[249] br[249] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_250 bl[250] br[250] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_251 bl[251] br[251] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_252 bl[252] br[252] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_253 bl[253] br[253] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_254 bl[254] br[254] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_255 bl[255] br[255] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_53_0 bl[0] br[0] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_1 bl[1] br[1] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_2 bl[2] br[2] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_3 bl[3] br[3] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_4 bl[4] br[4] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_5 bl[5] br[5] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_6 bl[6] br[6] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_7 bl[7] br[7] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_8 bl[8] br[8] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_9 bl[9] br[9] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_10 bl[10] br[10] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_11 bl[11] br[11] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_12 bl[12] br[12] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_13 bl[13] br[13] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_14 bl[14] br[14] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_15 bl[15] br[15] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_16 bl[16] br[16] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_17 bl[17] br[17] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_18 bl[18] br[18] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_19 bl[19] br[19] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_20 bl[20] br[20] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_21 bl[21] br[21] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_22 bl[22] br[22] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_23 bl[23] br[23] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_24 bl[24] br[24] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_25 bl[25] br[25] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_26 bl[26] br[26] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_27 bl[27] br[27] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_28 bl[28] br[28] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_29 bl[29] br[29] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_30 bl[30] br[30] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_31 bl[31] br[31] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_32 bl[32] br[32] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_33 bl[33] br[33] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_34 bl[34] br[34] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_35 bl[35] br[35] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_36 bl[36] br[36] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_37 bl[37] br[37] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_38 bl[38] br[38] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_39 bl[39] br[39] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_40 bl[40] br[40] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_41 bl[41] br[41] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_42 bl[42] br[42] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_43 bl[43] br[43] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_44 bl[44] br[44] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_45 bl[45] br[45] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_46 bl[46] br[46] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_47 bl[47] br[47] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_48 bl[48] br[48] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_49 bl[49] br[49] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_50 bl[50] br[50] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_51 bl[51] br[51] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_52 bl[52] br[52] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_53 bl[53] br[53] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_54 bl[54] br[54] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_55 bl[55] br[55] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_56 bl[56] br[56] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_57 bl[57] br[57] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_58 bl[58] br[58] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_59 bl[59] br[59] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_60 bl[60] br[60] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_61 bl[61] br[61] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_62 bl[62] br[62] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_63 bl[63] br[63] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_64 bl[64] br[64] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_65 bl[65] br[65] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_66 bl[66] br[66] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_67 bl[67] br[67] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_68 bl[68] br[68] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_69 bl[69] br[69] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_70 bl[70] br[70] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_71 bl[71] br[71] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_72 bl[72] br[72] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_73 bl[73] br[73] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_74 bl[74] br[74] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_75 bl[75] br[75] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_76 bl[76] br[76] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_77 bl[77] br[77] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_78 bl[78] br[78] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_79 bl[79] br[79] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_80 bl[80] br[80] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_81 bl[81] br[81] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_82 bl[82] br[82] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_83 bl[83] br[83] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_84 bl[84] br[84] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_85 bl[85] br[85] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_86 bl[86] br[86] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_87 bl[87] br[87] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_88 bl[88] br[88] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_89 bl[89] br[89] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_90 bl[90] br[90] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_91 bl[91] br[91] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_92 bl[92] br[92] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_93 bl[93] br[93] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_94 bl[94] br[94] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_95 bl[95] br[95] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_96 bl[96] br[96] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_97 bl[97] br[97] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_98 bl[98] br[98] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_99 bl[99] br[99] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_100 bl[100] br[100] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_101 bl[101] br[101] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_102 bl[102] br[102] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_103 bl[103] br[103] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_104 bl[104] br[104] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_105 bl[105] br[105] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_106 bl[106] br[106] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_107 bl[107] br[107] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_108 bl[108] br[108] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_109 bl[109] br[109] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_110 bl[110] br[110] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_111 bl[111] br[111] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_112 bl[112] br[112] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_113 bl[113] br[113] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_114 bl[114] br[114] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_115 bl[115] br[115] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_116 bl[116] br[116] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_117 bl[117] br[117] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_118 bl[118] br[118] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_119 bl[119] br[119] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_120 bl[120] br[120] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_121 bl[121] br[121] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_122 bl[122] br[122] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_123 bl[123] br[123] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_124 bl[124] br[124] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_125 bl[125] br[125] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_126 bl[126] br[126] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_127 bl[127] br[127] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_128 bl[128] br[128] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_129 bl[129] br[129] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_130 bl[130] br[130] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_131 bl[131] br[131] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_132 bl[132] br[132] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_133 bl[133] br[133] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_134 bl[134] br[134] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_135 bl[135] br[135] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_136 bl[136] br[136] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_137 bl[137] br[137] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_138 bl[138] br[138] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_139 bl[139] br[139] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_140 bl[140] br[140] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_141 bl[141] br[141] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_142 bl[142] br[142] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_143 bl[143] br[143] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_144 bl[144] br[144] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_145 bl[145] br[145] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_146 bl[146] br[146] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_147 bl[147] br[147] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_148 bl[148] br[148] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_149 bl[149] br[149] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_150 bl[150] br[150] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_151 bl[151] br[151] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_152 bl[152] br[152] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_153 bl[153] br[153] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_154 bl[154] br[154] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_155 bl[155] br[155] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_156 bl[156] br[156] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_157 bl[157] br[157] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_158 bl[158] br[158] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_159 bl[159] br[159] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_160 bl[160] br[160] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_161 bl[161] br[161] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_162 bl[162] br[162] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_163 bl[163] br[163] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_164 bl[164] br[164] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_165 bl[165] br[165] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_166 bl[166] br[166] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_167 bl[167] br[167] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_168 bl[168] br[168] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_169 bl[169] br[169] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_170 bl[170] br[170] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_171 bl[171] br[171] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_172 bl[172] br[172] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_173 bl[173] br[173] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_174 bl[174] br[174] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_175 bl[175] br[175] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_176 bl[176] br[176] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_177 bl[177] br[177] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_178 bl[178] br[178] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_179 bl[179] br[179] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_180 bl[180] br[180] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_181 bl[181] br[181] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_182 bl[182] br[182] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_183 bl[183] br[183] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_184 bl[184] br[184] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_185 bl[185] br[185] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_186 bl[186] br[186] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_187 bl[187] br[187] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_188 bl[188] br[188] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_189 bl[189] br[189] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_190 bl[190] br[190] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_191 bl[191] br[191] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_192 bl[192] br[192] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_193 bl[193] br[193] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_194 bl[194] br[194] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_195 bl[195] br[195] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_196 bl[196] br[196] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_197 bl[197] br[197] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_198 bl[198] br[198] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_199 bl[199] br[199] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_200 bl[200] br[200] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_201 bl[201] br[201] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_202 bl[202] br[202] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_203 bl[203] br[203] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_204 bl[204] br[204] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_205 bl[205] br[205] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_206 bl[206] br[206] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_207 bl[207] br[207] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_208 bl[208] br[208] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_209 bl[209] br[209] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_210 bl[210] br[210] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_211 bl[211] br[211] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_212 bl[212] br[212] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_213 bl[213] br[213] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_214 bl[214] br[214] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_215 bl[215] br[215] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_216 bl[216] br[216] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_217 bl[217] br[217] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_218 bl[218] br[218] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_219 bl[219] br[219] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_220 bl[220] br[220] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_221 bl[221] br[221] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_222 bl[222] br[222] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_223 bl[223] br[223] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_224 bl[224] br[224] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_225 bl[225] br[225] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_226 bl[226] br[226] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_227 bl[227] br[227] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_228 bl[228] br[228] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_229 bl[229] br[229] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_230 bl[230] br[230] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_231 bl[231] br[231] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_232 bl[232] br[232] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_233 bl[233] br[233] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_234 bl[234] br[234] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_235 bl[235] br[235] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_236 bl[236] br[236] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_237 bl[237] br[237] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_238 bl[238] br[238] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_239 bl[239] br[239] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_240 bl[240] br[240] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_241 bl[241] br[241] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_242 bl[242] br[242] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_243 bl[243] br[243] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_244 bl[244] br[244] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_245 bl[245] br[245] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_246 bl[246] br[246] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_247 bl[247] br[247] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_248 bl[248] br[248] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_249 bl[249] br[249] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_250 bl[250] br[250] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_251 bl[251] br[251] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_252 bl[252] br[252] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_253 bl[253] br[253] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_254 bl[254] br[254] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_255 bl[255] br[255] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_54_0 bl[0] br[0] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_1 bl[1] br[1] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_2 bl[2] br[2] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_3 bl[3] br[3] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_4 bl[4] br[4] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_5 bl[5] br[5] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_6 bl[6] br[6] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_7 bl[7] br[7] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_8 bl[8] br[8] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_9 bl[9] br[9] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_10 bl[10] br[10] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_11 bl[11] br[11] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_12 bl[12] br[12] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_13 bl[13] br[13] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_14 bl[14] br[14] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_15 bl[15] br[15] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_16 bl[16] br[16] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_17 bl[17] br[17] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_18 bl[18] br[18] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_19 bl[19] br[19] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_20 bl[20] br[20] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_21 bl[21] br[21] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_22 bl[22] br[22] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_23 bl[23] br[23] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_24 bl[24] br[24] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_25 bl[25] br[25] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_26 bl[26] br[26] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_27 bl[27] br[27] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_28 bl[28] br[28] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_29 bl[29] br[29] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_30 bl[30] br[30] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_31 bl[31] br[31] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_32 bl[32] br[32] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_33 bl[33] br[33] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_34 bl[34] br[34] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_35 bl[35] br[35] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_36 bl[36] br[36] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_37 bl[37] br[37] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_38 bl[38] br[38] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_39 bl[39] br[39] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_40 bl[40] br[40] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_41 bl[41] br[41] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_42 bl[42] br[42] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_43 bl[43] br[43] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_44 bl[44] br[44] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_45 bl[45] br[45] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_46 bl[46] br[46] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_47 bl[47] br[47] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_48 bl[48] br[48] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_49 bl[49] br[49] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_50 bl[50] br[50] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_51 bl[51] br[51] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_52 bl[52] br[52] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_53 bl[53] br[53] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_54 bl[54] br[54] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_55 bl[55] br[55] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_56 bl[56] br[56] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_57 bl[57] br[57] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_58 bl[58] br[58] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_59 bl[59] br[59] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_60 bl[60] br[60] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_61 bl[61] br[61] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_62 bl[62] br[62] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_63 bl[63] br[63] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_64 bl[64] br[64] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_65 bl[65] br[65] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_66 bl[66] br[66] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_67 bl[67] br[67] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_68 bl[68] br[68] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_69 bl[69] br[69] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_70 bl[70] br[70] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_71 bl[71] br[71] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_72 bl[72] br[72] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_73 bl[73] br[73] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_74 bl[74] br[74] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_75 bl[75] br[75] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_76 bl[76] br[76] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_77 bl[77] br[77] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_78 bl[78] br[78] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_79 bl[79] br[79] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_80 bl[80] br[80] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_81 bl[81] br[81] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_82 bl[82] br[82] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_83 bl[83] br[83] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_84 bl[84] br[84] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_85 bl[85] br[85] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_86 bl[86] br[86] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_87 bl[87] br[87] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_88 bl[88] br[88] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_89 bl[89] br[89] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_90 bl[90] br[90] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_91 bl[91] br[91] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_92 bl[92] br[92] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_93 bl[93] br[93] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_94 bl[94] br[94] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_95 bl[95] br[95] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_96 bl[96] br[96] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_97 bl[97] br[97] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_98 bl[98] br[98] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_99 bl[99] br[99] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_100 bl[100] br[100] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_101 bl[101] br[101] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_102 bl[102] br[102] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_103 bl[103] br[103] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_104 bl[104] br[104] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_105 bl[105] br[105] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_106 bl[106] br[106] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_107 bl[107] br[107] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_108 bl[108] br[108] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_109 bl[109] br[109] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_110 bl[110] br[110] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_111 bl[111] br[111] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_112 bl[112] br[112] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_113 bl[113] br[113] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_114 bl[114] br[114] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_115 bl[115] br[115] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_116 bl[116] br[116] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_117 bl[117] br[117] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_118 bl[118] br[118] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_119 bl[119] br[119] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_120 bl[120] br[120] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_121 bl[121] br[121] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_122 bl[122] br[122] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_123 bl[123] br[123] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_124 bl[124] br[124] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_125 bl[125] br[125] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_126 bl[126] br[126] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_127 bl[127] br[127] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_128 bl[128] br[128] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_129 bl[129] br[129] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_130 bl[130] br[130] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_131 bl[131] br[131] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_132 bl[132] br[132] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_133 bl[133] br[133] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_134 bl[134] br[134] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_135 bl[135] br[135] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_136 bl[136] br[136] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_137 bl[137] br[137] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_138 bl[138] br[138] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_139 bl[139] br[139] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_140 bl[140] br[140] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_141 bl[141] br[141] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_142 bl[142] br[142] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_143 bl[143] br[143] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_144 bl[144] br[144] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_145 bl[145] br[145] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_146 bl[146] br[146] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_147 bl[147] br[147] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_148 bl[148] br[148] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_149 bl[149] br[149] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_150 bl[150] br[150] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_151 bl[151] br[151] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_152 bl[152] br[152] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_153 bl[153] br[153] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_154 bl[154] br[154] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_155 bl[155] br[155] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_156 bl[156] br[156] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_157 bl[157] br[157] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_158 bl[158] br[158] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_159 bl[159] br[159] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_160 bl[160] br[160] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_161 bl[161] br[161] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_162 bl[162] br[162] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_163 bl[163] br[163] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_164 bl[164] br[164] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_165 bl[165] br[165] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_166 bl[166] br[166] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_167 bl[167] br[167] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_168 bl[168] br[168] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_169 bl[169] br[169] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_170 bl[170] br[170] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_171 bl[171] br[171] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_172 bl[172] br[172] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_173 bl[173] br[173] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_174 bl[174] br[174] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_175 bl[175] br[175] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_176 bl[176] br[176] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_177 bl[177] br[177] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_178 bl[178] br[178] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_179 bl[179] br[179] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_180 bl[180] br[180] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_181 bl[181] br[181] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_182 bl[182] br[182] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_183 bl[183] br[183] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_184 bl[184] br[184] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_185 bl[185] br[185] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_186 bl[186] br[186] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_187 bl[187] br[187] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_188 bl[188] br[188] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_189 bl[189] br[189] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_190 bl[190] br[190] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_191 bl[191] br[191] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_192 bl[192] br[192] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_193 bl[193] br[193] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_194 bl[194] br[194] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_195 bl[195] br[195] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_196 bl[196] br[196] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_197 bl[197] br[197] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_198 bl[198] br[198] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_199 bl[199] br[199] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_200 bl[200] br[200] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_201 bl[201] br[201] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_202 bl[202] br[202] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_203 bl[203] br[203] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_204 bl[204] br[204] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_205 bl[205] br[205] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_206 bl[206] br[206] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_207 bl[207] br[207] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_208 bl[208] br[208] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_209 bl[209] br[209] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_210 bl[210] br[210] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_211 bl[211] br[211] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_212 bl[212] br[212] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_213 bl[213] br[213] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_214 bl[214] br[214] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_215 bl[215] br[215] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_216 bl[216] br[216] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_217 bl[217] br[217] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_218 bl[218] br[218] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_219 bl[219] br[219] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_220 bl[220] br[220] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_221 bl[221] br[221] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_222 bl[222] br[222] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_223 bl[223] br[223] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_224 bl[224] br[224] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_225 bl[225] br[225] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_226 bl[226] br[226] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_227 bl[227] br[227] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_228 bl[228] br[228] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_229 bl[229] br[229] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_230 bl[230] br[230] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_231 bl[231] br[231] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_232 bl[232] br[232] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_233 bl[233] br[233] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_234 bl[234] br[234] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_235 bl[235] br[235] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_236 bl[236] br[236] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_237 bl[237] br[237] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_238 bl[238] br[238] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_239 bl[239] br[239] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_240 bl[240] br[240] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_241 bl[241] br[241] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_242 bl[242] br[242] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_243 bl[243] br[243] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_244 bl[244] br[244] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_245 bl[245] br[245] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_246 bl[246] br[246] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_247 bl[247] br[247] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_248 bl[248] br[248] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_249 bl[249] br[249] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_250 bl[250] br[250] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_251 bl[251] br[251] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_252 bl[252] br[252] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_253 bl[253] br[253] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_254 bl[254] br[254] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_255 bl[255] br[255] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_55_0 bl[0] br[0] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_1 bl[1] br[1] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_2 bl[2] br[2] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_3 bl[3] br[3] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_4 bl[4] br[4] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_5 bl[5] br[5] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_6 bl[6] br[6] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_7 bl[7] br[7] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_8 bl[8] br[8] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_9 bl[9] br[9] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_10 bl[10] br[10] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_11 bl[11] br[11] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_12 bl[12] br[12] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_13 bl[13] br[13] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_14 bl[14] br[14] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_15 bl[15] br[15] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_16 bl[16] br[16] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_17 bl[17] br[17] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_18 bl[18] br[18] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_19 bl[19] br[19] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_20 bl[20] br[20] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_21 bl[21] br[21] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_22 bl[22] br[22] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_23 bl[23] br[23] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_24 bl[24] br[24] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_25 bl[25] br[25] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_26 bl[26] br[26] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_27 bl[27] br[27] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_28 bl[28] br[28] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_29 bl[29] br[29] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_30 bl[30] br[30] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_31 bl[31] br[31] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_32 bl[32] br[32] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_33 bl[33] br[33] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_34 bl[34] br[34] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_35 bl[35] br[35] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_36 bl[36] br[36] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_37 bl[37] br[37] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_38 bl[38] br[38] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_39 bl[39] br[39] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_40 bl[40] br[40] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_41 bl[41] br[41] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_42 bl[42] br[42] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_43 bl[43] br[43] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_44 bl[44] br[44] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_45 bl[45] br[45] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_46 bl[46] br[46] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_47 bl[47] br[47] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_48 bl[48] br[48] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_49 bl[49] br[49] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_50 bl[50] br[50] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_51 bl[51] br[51] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_52 bl[52] br[52] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_53 bl[53] br[53] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_54 bl[54] br[54] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_55 bl[55] br[55] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_56 bl[56] br[56] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_57 bl[57] br[57] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_58 bl[58] br[58] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_59 bl[59] br[59] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_60 bl[60] br[60] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_61 bl[61] br[61] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_62 bl[62] br[62] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_63 bl[63] br[63] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_64 bl[64] br[64] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_65 bl[65] br[65] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_66 bl[66] br[66] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_67 bl[67] br[67] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_68 bl[68] br[68] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_69 bl[69] br[69] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_70 bl[70] br[70] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_71 bl[71] br[71] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_72 bl[72] br[72] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_73 bl[73] br[73] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_74 bl[74] br[74] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_75 bl[75] br[75] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_76 bl[76] br[76] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_77 bl[77] br[77] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_78 bl[78] br[78] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_79 bl[79] br[79] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_80 bl[80] br[80] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_81 bl[81] br[81] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_82 bl[82] br[82] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_83 bl[83] br[83] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_84 bl[84] br[84] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_85 bl[85] br[85] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_86 bl[86] br[86] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_87 bl[87] br[87] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_88 bl[88] br[88] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_89 bl[89] br[89] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_90 bl[90] br[90] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_91 bl[91] br[91] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_92 bl[92] br[92] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_93 bl[93] br[93] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_94 bl[94] br[94] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_95 bl[95] br[95] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_96 bl[96] br[96] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_97 bl[97] br[97] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_98 bl[98] br[98] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_99 bl[99] br[99] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_100 bl[100] br[100] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_101 bl[101] br[101] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_102 bl[102] br[102] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_103 bl[103] br[103] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_104 bl[104] br[104] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_105 bl[105] br[105] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_106 bl[106] br[106] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_107 bl[107] br[107] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_108 bl[108] br[108] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_109 bl[109] br[109] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_110 bl[110] br[110] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_111 bl[111] br[111] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_112 bl[112] br[112] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_113 bl[113] br[113] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_114 bl[114] br[114] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_115 bl[115] br[115] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_116 bl[116] br[116] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_117 bl[117] br[117] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_118 bl[118] br[118] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_119 bl[119] br[119] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_120 bl[120] br[120] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_121 bl[121] br[121] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_122 bl[122] br[122] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_123 bl[123] br[123] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_124 bl[124] br[124] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_125 bl[125] br[125] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_126 bl[126] br[126] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_127 bl[127] br[127] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_128 bl[128] br[128] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_129 bl[129] br[129] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_130 bl[130] br[130] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_131 bl[131] br[131] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_132 bl[132] br[132] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_133 bl[133] br[133] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_134 bl[134] br[134] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_135 bl[135] br[135] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_136 bl[136] br[136] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_137 bl[137] br[137] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_138 bl[138] br[138] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_139 bl[139] br[139] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_140 bl[140] br[140] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_141 bl[141] br[141] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_142 bl[142] br[142] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_143 bl[143] br[143] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_144 bl[144] br[144] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_145 bl[145] br[145] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_146 bl[146] br[146] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_147 bl[147] br[147] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_148 bl[148] br[148] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_149 bl[149] br[149] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_150 bl[150] br[150] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_151 bl[151] br[151] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_152 bl[152] br[152] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_153 bl[153] br[153] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_154 bl[154] br[154] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_155 bl[155] br[155] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_156 bl[156] br[156] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_157 bl[157] br[157] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_158 bl[158] br[158] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_159 bl[159] br[159] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_160 bl[160] br[160] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_161 bl[161] br[161] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_162 bl[162] br[162] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_163 bl[163] br[163] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_164 bl[164] br[164] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_165 bl[165] br[165] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_166 bl[166] br[166] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_167 bl[167] br[167] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_168 bl[168] br[168] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_169 bl[169] br[169] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_170 bl[170] br[170] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_171 bl[171] br[171] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_172 bl[172] br[172] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_173 bl[173] br[173] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_174 bl[174] br[174] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_175 bl[175] br[175] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_176 bl[176] br[176] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_177 bl[177] br[177] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_178 bl[178] br[178] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_179 bl[179] br[179] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_180 bl[180] br[180] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_181 bl[181] br[181] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_182 bl[182] br[182] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_183 bl[183] br[183] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_184 bl[184] br[184] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_185 bl[185] br[185] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_186 bl[186] br[186] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_187 bl[187] br[187] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_188 bl[188] br[188] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_189 bl[189] br[189] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_190 bl[190] br[190] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_191 bl[191] br[191] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_192 bl[192] br[192] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_193 bl[193] br[193] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_194 bl[194] br[194] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_195 bl[195] br[195] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_196 bl[196] br[196] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_197 bl[197] br[197] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_198 bl[198] br[198] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_199 bl[199] br[199] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_200 bl[200] br[200] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_201 bl[201] br[201] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_202 bl[202] br[202] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_203 bl[203] br[203] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_204 bl[204] br[204] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_205 bl[205] br[205] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_206 bl[206] br[206] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_207 bl[207] br[207] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_208 bl[208] br[208] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_209 bl[209] br[209] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_210 bl[210] br[210] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_211 bl[211] br[211] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_212 bl[212] br[212] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_213 bl[213] br[213] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_214 bl[214] br[214] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_215 bl[215] br[215] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_216 bl[216] br[216] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_217 bl[217] br[217] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_218 bl[218] br[218] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_219 bl[219] br[219] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_220 bl[220] br[220] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_221 bl[221] br[221] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_222 bl[222] br[222] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_223 bl[223] br[223] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_224 bl[224] br[224] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_225 bl[225] br[225] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_226 bl[226] br[226] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_227 bl[227] br[227] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_228 bl[228] br[228] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_229 bl[229] br[229] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_230 bl[230] br[230] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_231 bl[231] br[231] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_232 bl[232] br[232] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_233 bl[233] br[233] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_234 bl[234] br[234] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_235 bl[235] br[235] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_236 bl[236] br[236] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_237 bl[237] br[237] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_238 bl[238] br[238] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_239 bl[239] br[239] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_240 bl[240] br[240] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_241 bl[241] br[241] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_242 bl[242] br[242] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_243 bl[243] br[243] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_244 bl[244] br[244] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_245 bl[245] br[245] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_246 bl[246] br[246] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_247 bl[247] br[247] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_248 bl[248] br[248] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_249 bl[249] br[249] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_250 bl[250] br[250] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_251 bl[251] br[251] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_252 bl[252] br[252] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_253 bl[253] br[253] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_254 bl[254] br[254] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_255 bl[255] br[255] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_56_0 bl[0] br[0] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_1 bl[1] br[1] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_2 bl[2] br[2] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_3 bl[3] br[3] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_4 bl[4] br[4] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_5 bl[5] br[5] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_6 bl[6] br[6] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_7 bl[7] br[7] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_8 bl[8] br[8] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_9 bl[9] br[9] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_10 bl[10] br[10] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_11 bl[11] br[11] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_12 bl[12] br[12] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_13 bl[13] br[13] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_14 bl[14] br[14] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_15 bl[15] br[15] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_16 bl[16] br[16] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_17 bl[17] br[17] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_18 bl[18] br[18] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_19 bl[19] br[19] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_20 bl[20] br[20] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_21 bl[21] br[21] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_22 bl[22] br[22] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_23 bl[23] br[23] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_24 bl[24] br[24] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_25 bl[25] br[25] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_26 bl[26] br[26] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_27 bl[27] br[27] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_28 bl[28] br[28] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_29 bl[29] br[29] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_30 bl[30] br[30] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_31 bl[31] br[31] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_32 bl[32] br[32] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_33 bl[33] br[33] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_34 bl[34] br[34] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_35 bl[35] br[35] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_36 bl[36] br[36] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_37 bl[37] br[37] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_38 bl[38] br[38] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_39 bl[39] br[39] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_40 bl[40] br[40] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_41 bl[41] br[41] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_42 bl[42] br[42] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_43 bl[43] br[43] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_44 bl[44] br[44] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_45 bl[45] br[45] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_46 bl[46] br[46] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_47 bl[47] br[47] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_48 bl[48] br[48] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_49 bl[49] br[49] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_50 bl[50] br[50] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_51 bl[51] br[51] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_52 bl[52] br[52] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_53 bl[53] br[53] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_54 bl[54] br[54] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_55 bl[55] br[55] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_56 bl[56] br[56] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_57 bl[57] br[57] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_58 bl[58] br[58] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_59 bl[59] br[59] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_60 bl[60] br[60] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_61 bl[61] br[61] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_62 bl[62] br[62] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_63 bl[63] br[63] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_64 bl[64] br[64] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_65 bl[65] br[65] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_66 bl[66] br[66] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_67 bl[67] br[67] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_68 bl[68] br[68] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_69 bl[69] br[69] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_70 bl[70] br[70] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_71 bl[71] br[71] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_72 bl[72] br[72] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_73 bl[73] br[73] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_74 bl[74] br[74] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_75 bl[75] br[75] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_76 bl[76] br[76] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_77 bl[77] br[77] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_78 bl[78] br[78] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_79 bl[79] br[79] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_80 bl[80] br[80] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_81 bl[81] br[81] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_82 bl[82] br[82] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_83 bl[83] br[83] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_84 bl[84] br[84] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_85 bl[85] br[85] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_86 bl[86] br[86] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_87 bl[87] br[87] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_88 bl[88] br[88] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_89 bl[89] br[89] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_90 bl[90] br[90] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_91 bl[91] br[91] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_92 bl[92] br[92] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_93 bl[93] br[93] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_94 bl[94] br[94] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_95 bl[95] br[95] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_96 bl[96] br[96] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_97 bl[97] br[97] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_98 bl[98] br[98] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_99 bl[99] br[99] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_100 bl[100] br[100] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_101 bl[101] br[101] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_102 bl[102] br[102] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_103 bl[103] br[103] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_104 bl[104] br[104] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_105 bl[105] br[105] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_106 bl[106] br[106] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_107 bl[107] br[107] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_108 bl[108] br[108] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_109 bl[109] br[109] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_110 bl[110] br[110] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_111 bl[111] br[111] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_112 bl[112] br[112] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_113 bl[113] br[113] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_114 bl[114] br[114] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_115 bl[115] br[115] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_116 bl[116] br[116] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_117 bl[117] br[117] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_118 bl[118] br[118] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_119 bl[119] br[119] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_120 bl[120] br[120] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_121 bl[121] br[121] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_122 bl[122] br[122] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_123 bl[123] br[123] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_124 bl[124] br[124] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_125 bl[125] br[125] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_126 bl[126] br[126] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_127 bl[127] br[127] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_128 bl[128] br[128] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_129 bl[129] br[129] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_130 bl[130] br[130] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_131 bl[131] br[131] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_132 bl[132] br[132] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_133 bl[133] br[133] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_134 bl[134] br[134] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_135 bl[135] br[135] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_136 bl[136] br[136] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_137 bl[137] br[137] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_138 bl[138] br[138] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_139 bl[139] br[139] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_140 bl[140] br[140] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_141 bl[141] br[141] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_142 bl[142] br[142] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_143 bl[143] br[143] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_144 bl[144] br[144] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_145 bl[145] br[145] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_146 bl[146] br[146] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_147 bl[147] br[147] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_148 bl[148] br[148] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_149 bl[149] br[149] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_150 bl[150] br[150] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_151 bl[151] br[151] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_152 bl[152] br[152] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_153 bl[153] br[153] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_154 bl[154] br[154] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_155 bl[155] br[155] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_156 bl[156] br[156] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_157 bl[157] br[157] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_158 bl[158] br[158] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_159 bl[159] br[159] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_160 bl[160] br[160] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_161 bl[161] br[161] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_162 bl[162] br[162] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_163 bl[163] br[163] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_164 bl[164] br[164] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_165 bl[165] br[165] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_166 bl[166] br[166] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_167 bl[167] br[167] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_168 bl[168] br[168] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_169 bl[169] br[169] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_170 bl[170] br[170] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_171 bl[171] br[171] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_172 bl[172] br[172] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_173 bl[173] br[173] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_174 bl[174] br[174] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_175 bl[175] br[175] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_176 bl[176] br[176] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_177 bl[177] br[177] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_178 bl[178] br[178] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_179 bl[179] br[179] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_180 bl[180] br[180] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_181 bl[181] br[181] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_182 bl[182] br[182] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_183 bl[183] br[183] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_184 bl[184] br[184] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_185 bl[185] br[185] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_186 bl[186] br[186] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_187 bl[187] br[187] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_188 bl[188] br[188] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_189 bl[189] br[189] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_190 bl[190] br[190] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_191 bl[191] br[191] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_192 bl[192] br[192] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_193 bl[193] br[193] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_194 bl[194] br[194] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_195 bl[195] br[195] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_196 bl[196] br[196] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_197 bl[197] br[197] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_198 bl[198] br[198] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_199 bl[199] br[199] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_200 bl[200] br[200] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_201 bl[201] br[201] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_202 bl[202] br[202] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_203 bl[203] br[203] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_204 bl[204] br[204] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_205 bl[205] br[205] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_206 bl[206] br[206] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_207 bl[207] br[207] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_208 bl[208] br[208] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_209 bl[209] br[209] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_210 bl[210] br[210] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_211 bl[211] br[211] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_212 bl[212] br[212] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_213 bl[213] br[213] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_214 bl[214] br[214] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_215 bl[215] br[215] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_216 bl[216] br[216] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_217 bl[217] br[217] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_218 bl[218] br[218] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_219 bl[219] br[219] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_220 bl[220] br[220] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_221 bl[221] br[221] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_222 bl[222] br[222] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_223 bl[223] br[223] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_224 bl[224] br[224] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_225 bl[225] br[225] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_226 bl[226] br[226] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_227 bl[227] br[227] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_228 bl[228] br[228] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_229 bl[229] br[229] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_230 bl[230] br[230] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_231 bl[231] br[231] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_232 bl[232] br[232] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_233 bl[233] br[233] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_234 bl[234] br[234] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_235 bl[235] br[235] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_236 bl[236] br[236] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_237 bl[237] br[237] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_238 bl[238] br[238] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_239 bl[239] br[239] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_240 bl[240] br[240] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_241 bl[241] br[241] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_242 bl[242] br[242] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_243 bl[243] br[243] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_244 bl[244] br[244] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_245 bl[245] br[245] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_246 bl[246] br[246] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_247 bl[247] br[247] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_248 bl[248] br[248] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_249 bl[249] br[249] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_250 bl[250] br[250] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_251 bl[251] br[251] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_252 bl[252] br[252] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_253 bl[253] br[253] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_254 bl[254] br[254] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_255 bl[255] br[255] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_57_0 bl[0] br[0] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_1 bl[1] br[1] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_2 bl[2] br[2] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_3 bl[3] br[3] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_4 bl[4] br[4] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_5 bl[5] br[5] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_6 bl[6] br[6] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_7 bl[7] br[7] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_8 bl[8] br[8] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_9 bl[9] br[9] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_10 bl[10] br[10] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_11 bl[11] br[11] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_12 bl[12] br[12] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_13 bl[13] br[13] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_14 bl[14] br[14] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_15 bl[15] br[15] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_16 bl[16] br[16] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_17 bl[17] br[17] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_18 bl[18] br[18] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_19 bl[19] br[19] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_20 bl[20] br[20] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_21 bl[21] br[21] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_22 bl[22] br[22] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_23 bl[23] br[23] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_24 bl[24] br[24] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_25 bl[25] br[25] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_26 bl[26] br[26] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_27 bl[27] br[27] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_28 bl[28] br[28] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_29 bl[29] br[29] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_30 bl[30] br[30] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_31 bl[31] br[31] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_32 bl[32] br[32] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_33 bl[33] br[33] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_34 bl[34] br[34] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_35 bl[35] br[35] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_36 bl[36] br[36] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_37 bl[37] br[37] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_38 bl[38] br[38] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_39 bl[39] br[39] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_40 bl[40] br[40] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_41 bl[41] br[41] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_42 bl[42] br[42] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_43 bl[43] br[43] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_44 bl[44] br[44] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_45 bl[45] br[45] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_46 bl[46] br[46] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_47 bl[47] br[47] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_48 bl[48] br[48] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_49 bl[49] br[49] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_50 bl[50] br[50] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_51 bl[51] br[51] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_52 bl[52] br[52] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_53 bl[53] br[53] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_54 bl[54] br[54] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_55 bl[55] br[55] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_56 bl[56] br[56] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_57 bl[57] br[57] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_58 bl[58] br[58] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_59 bl[59] br[59] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_60 bl[60] br[60] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_61 bl[61] br[61] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_62 bl[62] br[62] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_63 bl[63] br[63] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_64 bl[64] br[64] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_65 bl[65] br[65] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_66 bl[66] br[66] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_67 bl[67] br[67] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_68 bl[68] br[68] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_69 bl[69] br[69] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_70 bl[70] br[70] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_71 bl[71] br[71] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_72 bl[72] br[72] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_73 bl[73] br[73] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_74 bl[74] br[74] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_75 bl[75] br[75] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_76 bl[76] br[76] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_77 bl[77] br[77] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_78 bl[78] br[78] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_79 bl[79] br[79] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_80 bl[80] br[80] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_81 bl[81] br[81] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_82 bl[82] br[82] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_83 bl[83] br[83] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_84 bl[84] br[84] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_85 bl[85] br[85] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_86 bl[86] br[86] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_87 bl[87] br[87] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_88 bl[88] br[88] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_89 bl[89] br[89] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_90 bl[90] br[90] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_91 bl[91] br[91] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_92 bl[92] br[92] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_93 bl[93] br[93] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_94 bl[94] br[94] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_95 bl[95] br[95] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_96 bl[96] br[96] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_97 bl[97] br[97] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_98 bl[98] br[98] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_99 bl[99] br[99] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_100 bl[100] br[100] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_101 bl[101] br[101] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_102 bl[102] br[102] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_103 bl[103] br[103] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_104 bl[104] br[104] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_105 bl[105] br[105] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_106 bl[106] br[106] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_107 bl[107] br[107] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_108 bl[108] br[108] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_109 bl[109] br[109] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_110 bl[110] br[110] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_111 bl[111] br[111] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_112 bl[112] br[112] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_113 bl[113] br[113] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_114 bl[114] br[114] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_115 bl[115] br[115] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_116 bl[116] br[116] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_117 bl[117] br[117] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_118 bl[118] br[118] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_119 bl[119] br[119] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_120 bl[120] br[120] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_121 bl[121] br[121] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_122 bl[122] br[122] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_123 bl[123] br[123] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_124 bl[124] br[124] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_125 bl[125] br[125] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_126 bl[126] br[126] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_127 bl[127] br[127] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_128 bl[128] br[128] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_129 bl[129] br[129] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_130 bl[130] br[130] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_131 bl[131] br[131] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_132 bl[132] br[132] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_133 bl[133] br[133] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_134 bl[134] br[134] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_135 bl[135] br[135] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_136 bl[136] br[136] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_137 bl[137] br[137] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_138 bl[138] br[138] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_139 bl[139] br[139] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_140 bl[140] br[140] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_141 bl[141] br[141] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_142 bl[142] br[142] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_143 bl[143] br[143] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_144 bl[144] br[144] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_145 bl[145] br[145] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_146 bl[146] br[146] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_147 bl[147] br[147] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_148 bl[148] br[148] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_149 bl[149] br[149] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_150 bl[150] br[150] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_151 bl[151] br[151] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_152 bl[152] br[152] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_153 bl[153] br[153] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_154 bl[154] br[154] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_155 bl[155] br[155] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_156 bl[156] br[156] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_157 bl[157] br[157] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_158 bl[158] br[158] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_159 bl[159] br[159] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_160 bl[160] br[160] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_161 bl[161] br[161] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_162 bl[162] br[162] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_163 bl[163] br[163] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_164 bl[164] br[164] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_165 bl[165] br[165] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_166 bl[166] br[166] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_167 bl[167] br[167] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_168 bl[168] br[168] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_169 bl[169] br[169] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_170 bl[170] br[170] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_171 bl[171] br[171] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_172 bl[172] br[172] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_173 bl[173] br[173] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_174 bl[174] br[174] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_175 bl[175] br[175] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_176 bl[176] br[176] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_177 bl[177] br[177] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_178 bl[178] br[178] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_179 bl[179] br[179] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_180 bl[180] br[180] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_181 bl[181] br[181] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_182 bl[182] br[182] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_183 bl[183] br[183] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_184 bl[184] br[184] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_185 bl[185] br[185] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_186 bl[186] br[186] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_187 bl[187] br[187] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_188 bl[188] br[188] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_189 bl[189] br[189] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_190 bl[190] br[190] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_191 bl[191] br[191] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_192 bl[192] br[192] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_193 bl[193] br[193] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_194 bl[194] br[194] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_195 bl[195] br[195] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_196 bl[196] br[196] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_197 bl[197] br[197] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_198 bl[198] br[198] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_199 bl[199] br[199] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_200 bl[200] br[200] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_201 bl[201] br[201] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_202 bl[202] br[202] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_203 bl[203] br[203] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_204 bl[204] br[204] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_205 bl[205] br[205] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_206 bl[206] br[206] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_207 bl[207] br[207] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_208 bl[208] br[208] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_209 bl[209] br[209] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_210 bl[210] br[210] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_211 bl[211] br[211] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_212 bl[212] br[212] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_213 bl[213] br[213] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_214 bl[214] br[214] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_215 bl[215] br[215] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_216 bl[216] br[216] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_217 bl[217] br[217] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_218 bl[218] br[218] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_219 bl[219] br[219] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_220 bl[220] br[220] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_221 bl[221] br[221] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_222 bl[222] br[222] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_223 bl[223] br[223] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_224 bl[224] br[224] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_225 bl[225] br[225] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_226 bl[226] br[226] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_227 bl[227] br[227] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_228 bl[228] br[228] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_229 bl[229] br[229] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_230 bl[230] br[230] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_231 bl[231] br[231] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_232 bl[232] br[232] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_233 bl[233] br[233] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_234 bl[234] br[234] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_235 bl[235] br[235] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_236 bl[236] br[236] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_237 bl[237] br[237] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_238 bl[238] br[238] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_239 bl[239] br[239] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_240 bl[240] br[240] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_241 bl[241] br[241] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_242 bl[242] br[242] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_243 bl[243] br[243] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_244 bl[244] br[244] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_245 bl[245] br[245] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_246 bl[246] br[246] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_247 bl[247] br[247] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_248 bl[248] br[248] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_249 bl[249] br[249] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_250 bl[250] br[250] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_251 bl[251] br[251] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_252 bl[252] br[252] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_253 bl[253] br[253] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_254 bl[254] br[254] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_255 bl[255] br[255] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_58_0 bl[0] br[0] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_1 bl[1] br[1] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_2 bl[2] br[2] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_3 bl[3] br[3] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_4 bl[4] br[4] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_5 bl[5] br[5] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_6 bl[6] br[6] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_7 bl[7] br[7] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_8 bl[8] br[8] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_9 bl[9] br[9] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_10 bl[10] br[10] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_11 bl[11] br[11] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_12 bl[12] br[12] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_13 bl[13] br[13] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_14 bl[14] br[14] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_15 bl[15] br[15] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_16 bl[16] br[16] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_17 bl[17] br[17] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_18 bl[18] br[18] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_19 bl[19] br[19] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_20 bl[20] br[20] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_21 bl[21] br[21] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_22 bl[22] br[22] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_23 bl[23] br[23] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_24 bl[24] br[24] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_25 bl[25] br[25] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_26 bl[26] br[26] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_27 bl[27] br[27] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_28 bl[28] br[28] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_29 bl[29] br[29] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_30 bl[30] br[30] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_31 bl[31] br[31] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_32 bl[32] br[32] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_33 bl[33] br[33] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_34 bl[34] br[34] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_35 bl[35] br[35] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_36 bl[36] br[36] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_37 bl[37] br[37] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_38 bl[38] br[38] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_39 bl[39] br[39] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_40 bl[40] br[40] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_41 bl[41] br[41] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_42 bl[42] br[42] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_43 bl[43] br[43] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_44 bl[44] br[44] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_45 bl[45] br[45] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_46 bl[46] br[46] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_47 bl[47] br[47] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_48 bl[48] br[48] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_49 bl[49] br[49] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_50 bl[50] br[50] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_51 bl[51] br[51] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_52 bl[52] br[52] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_53 bl[53] br[53] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_54 bl[54] br[54] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_55 bl[55] br[55] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_56 bl[56] br[56] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_57 bl[57] br[57] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_58 bl[58] br[58] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_59 bl[59] br[59] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_60 bl[60] br[60] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_61 bl[61] br[61] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_62 bl[62] br[62] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_63 bl[63] br[63] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_64 bl[64] br[64] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_65 bl[65] br[65] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_66 bl[66] br[66] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_67 bl[67] br[67] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_68 bl[68] br[68] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_69 bl[69] br[69] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_70 bl[70] br[70] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_71 bl[71] br[71] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_72 bl[72] br[72] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_73 bl[73] br[73] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_74 bl[74] br[74] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_75 bl[75] br[75] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_76 bl[76] br[76] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_77 bl[77] br[77] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_78 bl[78] br[78] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_79 bl[79] br[79] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_80 bl[80] br[80] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_81 bl[81] br[81] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_82 bl[82] br[82] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_83 bl[83] br[83] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_84 bl[84] br[84] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_85 bl[85] br[85] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_86 bl[86] br[86] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_87 bl[87] br[87] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_88 bl[88] br[88] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_89 bl[89] br[89] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_90 bl[90] br[90] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_91 bl[91] br[91] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_92 bl[92] br[92] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_93 bl[93] br[93] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_94 bl[94] br[94] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_95 bl[95] br[95] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_96 bl[96] br[96] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_97 bl[97] br[97] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_98 bl[98] br[98] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_99 bl[99] br[99] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_100 bl[100] br[100] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_101 bl[101] br[101] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_102 bl[102] br[102] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_103 bl[103] br[103] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_104 bl[104] br[104] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_105 bl[105] br[105] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_106 bl[106] br[106] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_107 bl[107] br[107] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_108 bl[108] br[108] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_109 bl[109] br[109] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_110 bl[110] br[110] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_111 bl[111] br[111] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_112 bl[112] br[112] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_113 bl[113] br[113] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_114 bl[114] br[114] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_115 bl[115] br[115] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_116 bl[116] br[116] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_117 bl[117] br[117] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_118 bl[118] br[118] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_119 bl[119] br[119] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_120 bl[120] br[120] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_121 bl[121] br[121] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_122 bl[122] br[122] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_123 bl[123] br[123] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_124 bl[124] br[124] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_125 bl[125] br[125] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_126 bl[126] br[126] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_127 bl[127] br[127] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_128 bl[128] br[128] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_129 bl[129] br[129] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_130 bl[130] br[130] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_131 bl[131] br[131] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_132 bl[132] br[132] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_133 bl[133] br[133] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_134 bl[134] br[134] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_135 bl[135] br[135] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_136 bl[136] br[136] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_137 bl[137] br[137] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_138 bl[138] br[138] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_139 bl[139] br[139] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_140 bl[140] br[140] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_141 bl[141] br[141] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_142 bl[142] br[142] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_143 bl[143] br[143] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_144 bl[144] br[144] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_145 bl[145] br[145] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_146 bl[146] br[146] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_147 bl[147] br[147] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_148 bl[148] br[148] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_149 bl[149] br[149] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_150 bl[150] br[150] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_151 bl[151] br[151] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_152 bl[152] br[152] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_153 bl[153] br[153] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_154 bl[154] br[154] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_155 bl[155] br[155] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_156 bl[156] br[156] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_157 bl[157] br[157] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_158 bl[158] br[158] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_159 bl[159] br[159] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_160 bl[160] br[160] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_161 bl[161] br[161] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_162 bl[162] br[162] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_163 bl[163] br[163] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_164 bl[164] br[164] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_165 bl[165] br[165] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_166 bl[166] br[166] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_167 bl[167] br[167] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_168 bl[168] br[168] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_169 bl[169] br[169] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_170 bl[170] br[170] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_171 bl[171] br[171] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_172 bl[172] br[172] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_173 bl[173] br[173] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_174 bl[174] br[174] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_175 bl[175] br[175] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_176 bl[176] br[176] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_177 bl[177] br[177] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_178 bl[178] br[178] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_179 bl[179] br[179] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_180 bl[180] br[180] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_181 bl[181] br[181] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_182 bl[182] br[182] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_183 bl[183] br[183] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_184 bl[184] br[184] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_185 bl[185] br[185] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_186 bl[186] br[186] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_187 bl[187] br[187] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_188 bl[188] br[188] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_189 bl[189] br[189] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_190 bl[190] br[190] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_191 bl[191] br[191] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_192 bl[192] br[192] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_193 bl[193] br[193] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_194 bl[194] br[194] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_195 bl[195] br[195] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_196 bl[196] br[196] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_197 bl[197] br[197] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_198 bl[198] br[198] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_199 bl[199] br[199] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_200 bl[200] br[200] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_201 bl[201] br[201] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_202 bl[202] br[202] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_203 bl[203] br[203] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_204 bl[204] br[204] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_205 bl[205] br[205] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_206 bl[206] br[206] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_207 bl[207] br[207] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_208 bl[208] br[208] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_209 bl[209] br[209] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_210 bl[210] br[210] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_211 bl[211] br[211] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_212 bl[212] br[212] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_213 bl[213] br[213] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_214 bl[214] br[214] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_215 bl[215] br[215] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_216 bl[216] br[216] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_217 bl[217] br[217] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_218 bl[218] br[218] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_219 bl[219] br[219] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_220 bl[220] br[220] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_221 bl[221] br[221] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_222 bl[222] br[222] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_223 bl[223] br[223] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_224 bl[224] br[224] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_225 bl[225] br[225] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_226 bl[226] br[226] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_227 bl[227] br[227] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_228 bl[228] br[228] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_229 bl[229] br[229] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_230 bl[230] br[230] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_231 bl[231] br[231] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_232 bl[232] br[232] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_233 bl[233] br[233] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_234 bl[234] br[234] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_235 bl[235] br[235] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_236 bl[236] br[236] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_237 bl[237] br[237] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_238 bl[238] br[238] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_239 bl[239] br[239] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_240 bl[240] br[240] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_241 bl[241] br[241] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_242 bl[242] br[242] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_243 bl[243] br[243] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_244 bl[244] br[244] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_245 bl[245] br[245] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_246 bl[246] br[246] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_247 bl[247] br[247] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_248 bl[248] br[248] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_249 bl[249] br[249] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_250 bl[250] br[250] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_251 bl[251] br[251] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_252 bl[252] br[252] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_253 bl[253] br[253] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_254 bl[254] br[254] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_255 bl[255] br[255] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_59_0 bl[0] br[0] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_1 bl[1] br[1] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_2 bl[2] br[2] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_3 bl[3] br[3] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_4 bl[4] br[4] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_5 bl[5] br[5] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_6 bl[6] br[6] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_7 bl[7] br[7] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_8 bl[8] br[8] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_9 bl[9] br[9] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_10 bl[10] br[10] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_11 bl[11] br[11] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_12 bl[12] br[12] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_13 bl[13] br[13] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_14 bl[14] br[14] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_15 bl[15] br[15] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_16 bl[16] br[16] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_17 bl[17] br[17] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_18 bl[18] br[18] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_19 bl[19] br[19] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_20 bl[20] br[20] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_21 bl[21] br[21] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_22 bl[22] br[22] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_23 bl[23] br[23] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_24 bl[24] br[24] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_25 bl[25] br[25] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_26 bl[26] br[26] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_27 bl[27] br[27] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_28 bl[28] br[28] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_29 bl[29] br[29] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_30 bl[30] br[30] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_31 bl[31] br[31] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_32 bl[32] br[32] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_33 bl[33] br[33] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_34 bl[34] br[34] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_35 bl[35] br[35] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_36 bl[36] br[36] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_37 bl[37] br[37] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_38 bl[38] br[38] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_39 bl[39] br[39] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_40 bl[40] br[40] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_41 bl[41] br[41] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_42 bl[42] br[42] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_43 bl[43] br[43] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_44 bl[44] br[44] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_45 bl[45] br[45] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_46 bl[46] br[46] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_47 bl[47] br[47] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_48 bl[48] br[48] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_49 bl[49] br[49] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_50 bl[50] br[50] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_51 bl[51] br[51] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_52 bl[52] br[52] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_53 bl[53] br[53] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_54 bl[54] br[54] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_55 bl[55] br[55] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_56 bl[56] br[56] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_57 bl[57] br[57] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_58 bl[58] br[58] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_59 bl[59] br[59] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_60 bl[60] br[60] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_61 bl[61] br[61] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_62 bl[62] br[62] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_63 bl[63] br[63] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_64 bl[64] br[64] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_65 bl[65] br[65] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_66 bl[66] br[66] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_67 bl[67] br[67] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_68 bl[68] br[68] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_69 bl[69] br[69] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_70 bl[70] br[70] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_71 bl[71] br[71] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_72 bl[72] br[72] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_73 bl[73] br[73] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_74 bl[74] br[74] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_75 bl[75] br[75] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_76 bl[76] br[76] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_77 bl[77] br[77] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_78 bl[78] br[78] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_79 bl[79] br[79] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_80 bl[80] br[80] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_81 bl[81] br[81] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_82 bl[82] br[82] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_83 bl[83] br[83] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_84 bl[84] br[84] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_85 bl[85] br[85] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_86 bl[86] br[86] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_87 bl[87] br[87] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_88 bl[88] br[88] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_89 bl[89] br[89] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_90 bl[90] br[90] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_91 bl[91] br[91] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_92 bl[92] br[92] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_93 bl[93] br[93] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_94 bl[94] br[94] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_95 bl[95] br[95] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_96 bl[96] br[96] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_97 bl[97] br[97] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_98 bl[98] br[98] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_99 bl[99] br[99] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_100 bl[100] br[100] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_101 bl[101] br[101] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_102 bl[102] br[102] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_103 bl[103] br[103] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_104 bl[104] br[104] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_105 bl[105] br[105] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_106 bl[106] br[106] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_107 bl[107] br[107] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_108 bl[108] br[108] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_109 bl[109] br[109] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_110 bl[110] br[110] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_111 bl[111] br[111] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_112 bl[112] br[112] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_113 bl[113] br[113] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_114 bl[114] br[114] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_115 bl[115] br[115] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_116 bl[116] br[116] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_117 bl[117] br[117] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_118 bl[118] br[118] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_119 bl[119] br[119] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_120 bl[120] br[120] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_121 bl[121] br[121] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_122 bl[122] br[122] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_123 bl[123] br[123] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_124 bl[124] br[124] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_125 bl[125] br[125] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_126 bl[126] br[126] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_127 bl[127] br[127] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_128 bl[128] br[128] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_129 bl[129] br[129] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_130 bl[130] br[130] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_131 bl[131] br[131] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_132 bl[132] br[132] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_133 bl[133] br[133] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_134 bl[134] br[134] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_135 bl[135] br[135] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_136 bl[136] br[136] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_137 bl[137] br[137] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_138 bl[138] br[138] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_139 bl[139] br[139] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_140 bl[140] br[140] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_141 bl[141] br[141] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_142 bl[142] br[142] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_143 bl[143] br[143] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_144 bl[144] br[144] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_145 bl[145] br[145] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_146 bl[146] br[146] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_147 bl[147] br[147] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_148 bl[148] br[148] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_149 bl[149] br[149] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_150 bl[150] br[150] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_151 bl[151] br[151] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_152 bl[152] br[152] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_153 bl[153] br[153] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_154 bl[154] br[154] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_155 bl[155] br[155] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_156 bl[156] br[156] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_157 bl[157] br[157] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_158 bl[158] br[158] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_159 bl[159] br[159] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_160 bl[160] br[160] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_161 bl[161] br[161] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_162 bl[162] br[162] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_163 bl[163] br[163] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_164 bl[164] br[164] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_165 bl[165] br[165] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_166 bl[166] br[166] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_167 bl[167] br[167] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_168 bl[168] br[168] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_169 bl[169] br[169] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_170 bl[170] br[170] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_171 bl[171] br[171] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_172 bl[172] br[172] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_173 bl[173] br[173] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_174 bl[174] br[174] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_175 bl[175] br[175] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_176 bl[176] br[176] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_177 bl[177] br[177] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_178 bl[178] br[178] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_179 bl[179] br[179] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_180 bl[180] br[180] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_181 bl[181] br[181] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_182 bl[182] br[182] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_183 bl[183] br[183] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_184 bl[184] br[184] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_185 bl[185] br[185] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_186 bl[186] br[186] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_187 bl[187] br[187] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_188 bl[188] br[188] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_189 bl[189] br[189] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_190 bl[190] br[190] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_191 bl[191] br[191] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_192 bl[192] br[192] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_193 bl[193] br[193] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_194 bl[194] br[194] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_195 bl[195] br[195] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_196 bl[196] br[196] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_197 bl[197] br[197] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_198 bl[198] br[198] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_199 bl[199] br[199] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_200 bl[200] br[200] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_201 bl[201] br[201] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_202 bl[202] br[202] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_203 bl[203] br[203] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_204 bl[204] br[204] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_205 bl[205] br[205] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_206 bl[206] br[206] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_207 bl[207] br[207] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_208 bl[208] br[208] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_209 bl[209] br[209] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_210 bl[210] br[210] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_211 bl[211] br[211] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_212 bl[212] br[212] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_213 bl[213] br[213] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_214 bl[214] br[214] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_215 bl[215] br[215] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_216 bl[216] br[216] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_217 bl[217] br[217] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_218 bl[218] br[218] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_219 bl[219] br[219] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_220 bl[220] br[220] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_221 bl[221] br[221] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_222 bl[222] br[222] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_223 bl[223] br[223] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_224 bl[224] br[224] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_225 bl[225] br[225] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_226 bl[226] br[226] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_227 bl[227] br[227] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_228 bl[228] br[228] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_229 bl[229] br[229] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_230 bl[230] br[230] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_231 bl[231] br[231] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_232 bl[232] br[232] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_233 bl[233] br[233] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_234 bl[234] br[234] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_235 bl[235] br[235] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_236 bl[236] br[236] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_237 bl[237] br[237] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_238 bl[238] br[238] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_239 bl[239] br[239] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_240 bl[240] br[240] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_241 bl[241] br[241] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_242 bl[242] br[242] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_243 bl[243] br[243] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_244 bl[244] br[244] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_245 bl[245] br[245] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_246 bl[246] br[246] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_247 bl[247] br[247] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_248 bl[248] br[248] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_249 bl[249] br[249] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_250 bl[250] br[250] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_251 bl[251] br[251] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_252 bl[252] br[252] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_253 bl[253] br[253] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_254 bl[254] br[254] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_255 bl[255] br[255] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_60_0 bl[0] br[0] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_1 bl[1] br[1] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_2 bl[2] br[2] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_3 bl[3] br[3] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_4 bl[4] br[4] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_5 bl[5] br[5] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_6 bl[6] br[6] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_7 bl[7] br[7] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_8 bl[8] br[8] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_9 bl[9] br[9] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_10 bl[10] br[10] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_11 bl[11] br[11] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_12 bl[12] br[12] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_13 bl[13] br[13] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_14 bl[14] br[14] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_15 bl[15] br[15] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_16 bl[16] br[16] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_17 bl[17] br[17] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_18 bl[18] br[18] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_19 bl[19] br[19] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_20 bl[20] br[20] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_21 bl[21] br[21] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_22 bl[22] br[22] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_23 bl[23] br[23] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_24 bl[24] br[24] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_25 bl[25] br[25] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_26 bl[26] br[26] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_27 bl[27] br[27] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_28 bl[28] br[28] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_29 bl[29] br[29] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_30 bl[30] br[30] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_31 bl[31] br[31] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_32 bl[32] br[32] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_33 bl[33] br[33] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_34 bl[34] br[34] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_35 bl[35] br[35] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_36 bl[36] br[36] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_37 bl[37] br[37] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_38 bl[38] br[38] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_39 bl[39] br[39] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_40 bl[40] br[40] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_41 bl[41] br[41] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_42 bl[42] br[42] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_43 bl[43] br[43] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_44 bl[44] br[44] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_45 bl[45] br[45] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_46 bl[46] br[46] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_47 bl[47] br[47] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_48 bl[48] br[48] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_49 bl[49] br[49] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_50 bl[50] br[50] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_51 bl[51] br[51] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_52 bl[52] br[52] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_53 bl[53] br[53] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_54 bl[54] br[54] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_55 bl[55] br[55] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_56 bl[56] br[56] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_57 bl[57] br[57] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_58 bl[58] br[58] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_59 bl[59] br[59] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_60 bl[60] br[60] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_61 bl[61] br[61] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_62 bl[62] br[62] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_63 bl[63] br[63] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_64 bl[64] br[64] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_65 bl[65] br[65] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_66 bl[66] br[66] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_67 bl[67] br[67] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_68 bl[68] br[68] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_69 bl[69] br[69] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_70 bl[70] br[70] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_71 bl[71] br[71] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_72 bl[72] br[72] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_73 bl[73] br[73] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_74 bl[74] br[74] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_75 bl[75] br[75] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_76 bl[76] br[76] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_77 bl[77] br[77] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_78 bl[78] br[78] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_79 bl[79] br[79] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_80 bl[80] br[80] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_81 bl[81] br[81] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_82 bl[82] br[82] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_83 bl[83] br[83] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_84 bl[84] br[84] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_85 bl[85] br[85] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_86 bl[86] br[86] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_87 bl[87] br[87] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_88 bl[88] br[88] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_89 bl[89] br[89] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_90 bl[90] br[90] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_91 bl[91] br[91] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_92 bl[92] br[92] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_93 bl[93] br[93] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_94 bl[94] br[94] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_95 bl[95] br[95] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_96 bl[96] br[96] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_97 bl[97] br[97] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_98 bl[98] br[98] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_99 bl[99] br[99] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_100 bl[100] br[100] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_101 bl[101] br[101] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_102 bl[102] br[102] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_103 bl[103] br[103] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_104 bl[104] br[104] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_105 bl[105] br[105] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_106 bl[106] br[106] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_107 bl[107] br[107] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_108 bl[108] br[108] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_109 bl[109] br[109] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_110 bl[110] br[110] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_111 bl[111] br[111] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_112 bl[112] br[112] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_113 bl[113] br[113] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_114 bl[114] br[114] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_115 bl[115] br[115] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_116 bl[116] br[116] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_117 bl[117] br[117] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_118 bl[118] br[118] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_119 bl[119] br[119] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_120 bl[120] br[120] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_121 bl[121] br[121] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_122 bl[122] br[122] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_123 bl[123] br[123] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_124 bl[124] br[124] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_125 bl[125] br[125] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_126 bl[126] br[126] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_127 bl[127] br[127] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_128 bl[128] br[128] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_129 bl[129] br[129] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_130 bl[130] br[130] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_131 bl[131] br[131] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_132 bl[132] br[132] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_133 bl[133] br[133] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_134 bl[134] br[134] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_135 bl[135] br[135] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_136 bl[136] br[136] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_137 bl[137] br[137] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_138 bl[138] br[138] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_139 bl[139] br[139] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_140 bl[140] br[140] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_141 bl[141] br[141] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_142 bl[142] br[142] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_143 bl[143] br[143] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_144 bl[144] br[144] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_145 bl[145] br[145] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_146 bl[146] br[146] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_147 bl[147] br[147] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_148 bl[148] br[148] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_149 bl[149] br[149] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_150 bl[150] br[150] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_151 bl[151] br[151] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_152 bl[152] br[152] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_153 bl[153] br[153] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_154 bl[154] br[154] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_155 bl[155] br[155] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_156 bl[156] br[156] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_157 bl[157] br[157] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_158 bl[158] br[158] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_159 bl[159] br[159] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_160 bl[160] br[160] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_161 bl[161] br[161] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_162 bl[162] br[162] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_163 bl[163] br[163] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_164 bl[164] br[164] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_165 bl[165] br[165] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_166 bl[166] br[166] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_167 bl[167] br[167] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_168 bl[168] br[168] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_169 bl[169] br[169] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_170 bl[170] br[170] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_171 bl[171] br[171] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_172 bl[172] br[172] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_173 bl[173] br[173] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_174 bl[174] br[174] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_175 bl[175] br[175] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_176 bl[176] br[176] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_177 bl[177] br[177] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_178 bl[178] br[178] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_179 bl[179] br[179] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_180 bl[180] br[180] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_181 bl[181] br[181] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_182 bl[182] br[182] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_183 bl[183] br[183] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_184 bl[184] br[184] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_185 bl[185] br[185] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_186 bl[186] br[186] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_187 bl[187] br[187] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_188 bl[188] br[188] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_189 bl[189] br[189] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_190 bl[190] br[190] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_191 bl[191] br[191] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_192 bl[192] br[192] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_193 bl[193] br[193] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_194 bl[194] br[194] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_195 bl[195] br[195] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_196 bl[196] br[196] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_197 bl[197] br[197] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_198 bl[198] br[198] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_199 bl[199] br[199] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_200 bl[200] br[200] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_201 bl[201] br[201] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_202 bl[202] br[202] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_203 bl[203] br[203] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_204 bl[204] br[204] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_205 bl[205] br[205] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_206 bl[206] br[206] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_207 bl[207] br[207] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_208 bl[208] br[208] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_209 bl[209] br[209] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_210 bl[210] br[210] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_211 bl[211] br[211] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_212 bl[212] br[212] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_213 bl[213] br[213] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_214 bl[214] br[214] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_215 bl[215] br[215] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_216 bl[216] br[216] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_217 bl[217] br[217] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_218 bl[218] br[218] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_219 bl[219] br[219] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_220 bl[220] br[220] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_221 bl[221] br[221] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_222 bl[222] br[222] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_223 bl[223] br[223] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_224 bl[224] br[224] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_225 bl[225] br[225] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_226 bl[226] br[226] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_227 bl[227] br[227] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_228 bl[228] br[228] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_229 bl[229] br[229] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_230 bl[230] br[230] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_231 bl[231] br[231] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_232 bl[232] br[232] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_233 bl[233] br[233] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_234 bl[234] br[234] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_235 bl[235] br[235] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_236 bl[236] br[236] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_237 bl[237] br[237] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_238 bl[238] br[238] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_239 bl[239] br[239] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_240 bl[240] br[240] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_241 bl[241] br[241] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_242 bl[242] br[242] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_243 bl[243] br[243] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_244 bl[244] br[244] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_245 bl[245] br[245] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_246 bl[246] br[246] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_247 bl[247] br[247] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_248 bl[248] br[248] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_249 bl[249] br[249] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_250 bl[250] br[250] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_251 bl[251] br[251] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_252 bl[252] br[252] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_253 bl[253] br[253] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_254 bl[254] br[254] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_255 bl[255] br[255] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_61_0 bl[0] br[0] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_1 bl[1] br[1] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_2 bl[2] br[2] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_3 bl[3] br[3] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_4 bl[4] br[4] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_5 bl[5] br[5] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_6 bl[6] br[6] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_7 bl[7] br[7] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_8 bl[8] br[8] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_9 bl[9] br[9] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_10 bl[10] br[10] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_11 bl[11] br[11] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_12 bl[12] br[12] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_13 bl[13] br[13] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_14 bl[14] br[14] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_15 bl[15] br[15] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_16 bl[16] br[16] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_17 bl[17] br[17] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_18 bl[18] br[18] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_19 bl[19] br[19] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_20 bl[20] br[20] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_21 bl[21] br[21] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_22 bl[22] br[22] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_23 bl[23] br[23] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_24 bl[24] br[24] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_25 bl[25] br[25] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_26 bl[26] br[26] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_27 bl[27] br[27] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_28 bl[28] br[28] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_29 bl[29] br[29] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_30 bl[30] br[30] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_31 bl[31] br[31] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_32 bl[32] br[32] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_33 bl[33] br[33] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_34 bl[34] br[34] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_35 bl[35] br[35] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_36 bl[36] br[36] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_37 bl[37] br[37] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_38 bl[38] br[38] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_39 bl[39] br[39] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_40 bl[40] br[40] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_41 bl[41] br[41] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_42 bl[42] br[42] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_43 bl[43] br[43] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_44 bl[44] br[44] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_45 bl[45] br[45] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_46 bl[46] br[46] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_47 bl[47] br[47] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_48 bl[48] br[48] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_49 bl[49] br[49] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_50 bl[50] br[50] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_51 bl[51] br[51] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_52 bl[52] br[52] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_53 bl[53] br[53] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_54 bl[54] br[54] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_55 bl[55] br[55] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_56 bl[56] br[56] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_57 bl[57] br[57] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_58 bl[58] br[58] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_59 bl[59] br[59] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_60 bl[60] br[60] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_61 bl[61] br[61] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_62 bl[62] br[62] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_63 bl[63] br[63] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_64 bl[64] br[64] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_65 bl[65] br[65] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_66 bl[66] br[66] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_67 bl[67] br[67] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_68 bl[68] br[68] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_69 bl[69] br[69] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_70 bl[70] br[70] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_71 bl[71] br[71] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_72 bl[72] br[72] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_73 bl[73] br[73] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_74 bl[74] br[74] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_75 bl[75] br[75] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_76 bl[76] br[76] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_77 bl[77] br[77] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_78 bl[78] br[78] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_79 bl[79] br[79] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_80 bl[80] br[80] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_81 bl[81] br[81] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_82 bl[82] br[82] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_83 bl[83] br[83] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_84 bl[84] br[84] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_85 bl[85] br[85] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_86 bl[86] br[86] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_87 bl[87] br[87] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_88 bl[88] br[88] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_89 bl[89] br[89] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_90 bl[90] br[90] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_91 bl[91] br[91] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_92 bl[92] br[92] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_93 bl[93] br[93] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_94 bl[94] br[94] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_95 bl[95] br[95] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_96 bl[96] br[96] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_97 bl[97] br[97] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_98 bl[98] br[98] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_99 bl[99] br[99] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_100 bl[100] br[100] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_101 bl[101] br[101] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_102 bl[102] br[102] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_103 bl[103] br[103] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_104 bl[104] br[104] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_105 bl[105] br[105] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_106 bl[106] br[106] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_107 bl[107] br[107] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_108 bl[108] br[108] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_109 bl[109] br[109] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_110 bl[110] br[110] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_111 bl[111] br[111] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_112 bl[112] br[112] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_113 bl[113] br[113] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_114 bl[114] br[114] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_115 bl[115] br[115] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_116 bl[116] br[116] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_117 bl[117] br[117] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_118 bl[118] br[118] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_119 bl[119] br[119] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_120 bl[120] br[120] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_121 bl[121] br[121] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_122 bl[122] br[122] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_123 bl[123] br[123] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_124 bl[124] br[124] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_125 bl[125] br[125] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_126 bl[126] br[126] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_127 bl[127] br[127] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_128 bl[128] br[128] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_129 bl[129] br[129] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_130 bl[130] br[130] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_131 bl[131] br[131] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_132 bl[132] br[132] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_133 bl[133] br[133] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_134 bl[134] br[134] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_135 bl[135] br[135] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_136 bl[136] br[136] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_137 bl[137] br[137] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_138 bl[138] br[138] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_139 bl[139] br[139] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_140 bl[140] br[140] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_141 bl[141] br[141] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_142 bl[142] br[142] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_143 bl[143] br[143] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_144 bl[144] br[144] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_145 bl[145] br[145] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_146 bl[146] br[146] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_147 bl[147] br[147] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_148 bl[148] br[148] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_149 bl[149] br[149] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_150 bl[150] br[150] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_151 bl[151] br[151] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_152 bl[152] br[152] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_153 bl[153] br[153] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_154 bl[154] br[154] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_155 bl[155] br[155] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_156 bl[156] br[156] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_157 bl[157] br[157] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_158 bl[158] br[158] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_159 bl[159] br[159] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_160 bl[160] br[160] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_161 bl[161] br[161] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_162 bl[162] br[162] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_163 bl[163] br[163] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_164 bl[164] br[164] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_165 bl[165] br[165] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_166 bl[166] br[166] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_167 bl[167] br[167] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_168 bl[168] br[168] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_169 bl[169] br[169] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_170 bl[170] br[170] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_171 bl[171] br[171] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_172 bl[172] br[172] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_173 bl[173] br[173] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_174 bl[174] br[174] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_175 bl[175] br[175] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_176 bl[176] br[176] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_177 bl[177] br[177] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_178 bl[178] br[178] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_179 bl[179] br[179] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_180 bl[180] br[180] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_181 bl[181] br[181] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_182 bl[182] br[182] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_183 bl[183] br[183] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_184 bl[184] br[184] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_185 bl[185] br[185] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_186 bl[186] br[186] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_187 bl[187] br[187] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_188 bl[188] br[188] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_189 bl[189] br[189] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_190 bl[190] br[190] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_191 bl[191] br[191] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_192 bl[192] br[192] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_193 bl[193] br[193] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_194 bl[194] br[194] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_195 bl[195] br[195] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_196 bl[196] br[196] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_197 bl[197] br[197] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_198 bl[198] br[198] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_199 bl[199] br[199] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_200 bl[200] br[200] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_201 bl[201] br[201] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_202 bl[202] br[202] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_203 bl[203] br[203] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_204 bl[204] br[204] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_205 bl[205] br[205] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_206 bl[206] br[206] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_207 bl[207] br[207] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_208 bl[208] br[208] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_209 bl[209] br[209] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_210 bl[210] br[210] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_211 bl[211] br[211] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_212 bl[212] br[212] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_213 bl[213] br[213] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_214 bl[214] br[214] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_215 bl[215] br[215] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_216 bl[216] br[216] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_217 bl[217] br[217] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_218 bl[218] br[218] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_219 bl[219] br[219] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_220 bl[220] br[220] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_221 bl[221] br[221] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_222 bl[222] br[222] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_223 bl[223] br[223] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_224 bl[224] br[224] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_225 bl[225] br[225] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_226 bl[226] br[226] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_227 bl[227] br[227] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_228 bl[228] br[228] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_229 bl[229] br[229] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_230 bl[230] br[230] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_231 bl[231] br[231] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_232 bl[232] br[232] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_233 bl[233] br[233] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_234 bl[234] br[234] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_235 bl[235] br[235] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_236 bl[236] br[236] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_237 bl[237] br[237] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_238 bl[238] br[238] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_239 bl[239] br[239] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_240 bl[240] br[240] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_241 bl[241] br[241] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_242 bl[242] br[242] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_243 bl[243] br[243] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_244 bl[244] br[244] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_245 bl[245] br[245] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_246 bl[246] br[246] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_247 bl[247] br[247] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_248 bl[248] br[248] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_249 bl[249] br[249] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_250 bl[250] br[250] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_251 bl[251] br[251] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_252 bl[252] br[252] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_253 bl[253] br[253] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_254 bl[254] br[254] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_255 bl[255] br[255] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_62_0 bl[0] br[0] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_1 bl[1] br[1] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_2 bl[2] br[2] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_3 bl[3] br[3] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_4 bl[4] br[4] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_5 bl[5] br[5] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_6 bl[6] br[6] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_7 bl[7] br[7] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_8 bl[8] br[8] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_9 bl[9] br[9] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_10 bl[10] br[10] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_11 bl[11] br[11] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_12 bl[12] br[12] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_13 bl[13] br[13] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_14 bl[14] br[14] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_15 bl[15] br[15] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_16 bl[16] br[16] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_17 bl[17] br[17] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_18 bl[18] br[18] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_19 bl[19] br[19] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_20 bl[20] br[20] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_21 bl[21] br[21] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_22 bl[22] br[22] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_23 bl[23] br[23] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_24 bl[24] br[24] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_25 bl[25] br[25] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_26 bl[26] br[26] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_27 bl[27] br[27] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_28 bl[28] br[28] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_29 bl[29] br[29] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_30 bl[30] br[30] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_31 bl[31] br[31] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_32 bl[32] br[32] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_33 bl[33] br[33] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_34 bl[34] br[34] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_35 bl[35] br[35] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_36 bl[36] br[36] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_37 bl[37] br[37] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_38 bl[38] br[38] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_39 bl[39] br[39] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_40 bl[40] br[40] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_41 bl[41] br[41] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_42 bl[42] br[42] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_43 bl[43] br[43] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_44 bl[44] br[44] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_45 bl[45] br[45] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_46 bl[46] br[46] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_47 bl[47] br[47] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_48 bl[48] br[48] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_49 bl[49] br[49] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_50 bl[50] br[50] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_51 bl[51] br[51] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_52 bl[52] br[52] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_53 bl[53] br[53] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_54 bl[54] br[54] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_55 bl[55] br[55] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_56 bl[56] br[56] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_57 bl[57] br[57] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_58 bl[58] br[58] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_59 bl[59] br[59] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_60 bl[60] br[60] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_61 bl[61] br[61] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_62 bl[62] br[62] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_63 bl[63] br[63] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_64 bl[64] br[64] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_65 bl[65] br[65] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_66 bl[66] br[66] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_67 bl[67] br[67] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_68 bl[68] br[68] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_69 bl[69] br[69] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_70 bl[70] br[70] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_71 bl[71] br[71] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_72 bl[72] br[72] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_73 bl[73] br[73] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_74 bl[74] br[74] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_75 bl[75] br[75] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_76 bl[76] br[76] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_77 bl[77] br[77] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_78 bl[78] br[78] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_79 bl[79] br[79] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_80 bl[80] br[80] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_81 bl[81] br[81] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_82 bl[82] br[82] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_83 bl[83] br[83] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_84 bl[84] br[84] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_85 bl[85] br[85] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_86 bl[86] br[86] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_87 bl[87] br[87] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_88 bl[88] br[88] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_89 bl[89] br[89] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_90 bl[90] br[90] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_91 bl[91] br[91] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_92 bl[92] br[92] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_93 bl[93] br[93] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_94 bl[94] br[94] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_95 bl[95] br[95] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_96 bl[96] br[96] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_97 bl[97] br[97] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_98 bl[98] br[98] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_99 bl[99] br[99] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_100 bl[100] br[100] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_101 bl[101] br[101] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_102 bl[102] br[102] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_103 bl[103] br[103] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_104 bl[104] br[104] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_105 bl[105] br[105] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_106 bl[106] br[106] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_107 bl[107] br[107] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_108 bl[108] br[108] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_109 bl[109] br[109] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_110 bl[110] br[110] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_111 bl[111] br[111] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_112 bl[112] br[112] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_113 bl[113] br[113] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_114 bl[114] br[114] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_115 bl[115] br[115] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_116 bl[116] br[116] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_117 bl[117] br[117] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_118 bl[118] br[118] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_119 bl[119] br[119] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_120 bl[120] br[120] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_121 bl[121] br[121] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_122 bl[122] br[122] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_123 bl[123] br[123] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_124 bl[124] br[124] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_125 bl[125] br[125] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_126 bl[126] br[126] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_127 bl[127] br[127] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_128 bl[128] br[128] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_129 bl[129] br[129] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_130 bl[130] br[130] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_131 bl[131] br[131] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_132 bl[132] br[132] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_133 bl[133] br[133] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_134 bl[134] br[134] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_135 bl[135] br[135] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_136 bl[136] br[136] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_137 bl[137] br[137] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_138 bl[138] br[138] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_139 bl[139] br[139] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_140 bl[140] br[140] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_141 bl[141] br[141] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_142 bl[142] br[142] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_143 bl[143] br[143] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_144 bl[144] br[144] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_145 bl[145] br[145] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_146 bl[146] br[146] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_147 bl[147] br[147] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_148 bl[148] br[148] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_149 bl[149] br[149] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_150 bl[150] br[150] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_151 bl[151] br[151] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_152 bl[152] br[152] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_153 bl[153] br[153] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_154 bl[154] br[154] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_155 bl[155] br[155] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_156 bl[156] br[156] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_157 bl[157] br[157] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_158 bl[158] br[158] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_159 bl[159] br[159] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_160 bl[160] br[160] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_161 bl[161] br[161] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_162 bl[162] br[162] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_163 bl[163] br[163] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_164 bl[164] br[164] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_165 bl[165] br[165] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_166 bl[166] br[166] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_167 bl[167] br[167] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_168 bl[168] br[168] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_169 bl[169] br[169] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_170 bl[170] br[170] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_171 bl[171] br[171] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_172 bl[172] br[172] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_173 bl[173] br[173] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_174 bl[174] br[174] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_175 bl[175] br[175] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_176 bl[176] br[176] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_177 bl[177] br[177] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_178 bl[178] br[178] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_179 bl[179] br[179] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_180 bl[180] br[180] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_181 bl[181] br[181] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_182 bl[182] br[182] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_183 bl[183] br[183] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_184 bl[184] br[184] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_185 bl[185] br[185] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_186 bl[186] br[186] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_187 bl[187] br[187] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_188 bl[188] br[188] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_189 bl[189] br[189] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_190 bl[190] br[190] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_191 bl[191] br[191] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_192 bl[192] br[192] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_193 bl[193] br[193] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_194 bl[194] br[194] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_195 bl[195] br[195] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_196 bl[196] br[196] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_197 bl[197] br[197] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_198 bl[198] br[198] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_199 bl[199] br[199] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_200 bl[200] br[200] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_201 bl[201] br[201] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_202 bl[202] br[202] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_203 bl[203] br[203] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_204 bl[204] br[204] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_205 bl[205] br[205] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_206 bl[206] br[206] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_207 bl[207] br[207] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_208 bl[208] br[208] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_209 bl[209] br[209] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_210 bl[210] br[210] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_211 bl[211] br[211] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_212 bl[212] br[212] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_213 bl[213] br[213] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_214 bl[214] br[214] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_215 bl[215] br[215] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_216 bl[216] br[216] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_217 bl[217] br[217] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_218 bl[218] br[218] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_219 bl[219] br[219] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_220 bl[220] br[220] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_221 bl[221] br[221] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_222 bl[222] br[222] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_223 bl[223] br[223] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_224 bl[224] br[224] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_225 bl[225] br[225] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_226 bl[226] br[226] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_227 bl[227] br[227] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_228 bl[228] br[228] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_229 bl[229] br[229] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_230 bl[230] br[230] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_231 bl[231] br[231] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_232 bl[232] br[232] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_233 bl[233] br[233] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_234 bl[234] br[234] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_235 bl[235] br[235] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_236 bl[236] br[236] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_237 bl[237] br[237] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_238 bl[238] br[238] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_239 bl[239] br[239] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_240 bl[240] br[240] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_241 bl[241] br[241] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_242 bl[242] br[242] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_243 bl[243] br[243] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_244 bl[244] br[244] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_245 bl[245] br[245] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_246 bl[246] br[246] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_247 bl[247] br[247] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_248 bl[248] br[248] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_249 bl[249] br[249] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_250 bl[250] br[250] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_251 bl[251] br[251] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_252 bl[252] br[252] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_253 bl[253] br[253] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_254 bl[254] br[254] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_255 bl[255] br[255] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_63_0 bl[0] br[0] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_1 bl[1] br[1] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_2 bl[2] br[2] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_3 bl[3] br[3] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_4 bl[4] br[4] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_5 bl[5] br[5] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_6 bl[6] br[6] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_7 bl[7] br[7] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_8 bl[8] br[8] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_9 bl[9] br[9] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_10 bl[10] br[10] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_11 bl[11] br[11] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_12 bl[12] br[12] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_13 bl[13] br[13] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_14 bl[14] br[14] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_15 bl[15] br[15] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_16 bl[16] br[16] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_17 bl[17] br[17] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_18 bl[18] br[18] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_19 bl[19] br[19] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_20 bl[20] br[20] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_21 bl[21] br[21] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_22 bl[22] br[22] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_23 bl[23] br[23] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_24 bl[24] br[24] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_25 bl[25] br[25] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_26 bl[26] br[26] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_27 bl[27] br[27] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_28 bl[28] br[28] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_29 bl[29] br[29] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_30 bl[30] br[30] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_31 bl[31] br[31] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_32 bl[32] br[32] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_33 bl[33] br[33] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_34 bl[34] br[34] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_35 bl[35] br[35] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_36 bl[36] br[36] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_37 bl[37] br[37] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_38 bl[38] br[38] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_39 bl[39] br[39] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_40 bl[40] br[40] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_41 bl[41] br[41] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_42 bl[42] br[42] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_43 bl[43] br[43] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_44 bl[44] br[44] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_45 bl[45] br[45] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_46 bl[46] br[46] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_47 bl[47] br[47] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_48 bl[48] br[48] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_49 bl[49] br[49] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_50 bl[50] br[50] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_51 bl[51] br[51] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_52 bl[52] br[52] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_53 bl[53] br[53] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_54 bl[54] br[54] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_55 bl[55] br[55] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_56 bl[56] br[56] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_57 bl[57] br[57] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_58 bl[58] br[58] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_59 bl[59] br[59] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_60 bl[60] br[60] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_61 bl[61] br[61] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_62 bl[62] br[62] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_63 bl[63] br[63] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_64 bl[64] br[64] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_65 bl[65] br[65] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_66 bl[66] br[66] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_67 bl[67] br[67] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_68 bl[68] br[68] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_69 bl[69] br[69] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_70 bl[70] br[70] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_71 bl[71] br[71] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_72 bl[72] br[72] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_73 bl[73] br[73] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_74 bl[74] br[74] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_75 bl[75] br[75] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_76 bl[76] br[76] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_77 bl[77] br[77] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_78 bl[78] br[78] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_79 bl[79] br[79] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_80 bl[80] br[80] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_81 bl[81] br[81] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_82 bl[82] br[82] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_83 bl[83] br[83] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_84 bl[84] br[84] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_85 bl[85] br[85] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_86 bl[86] br[86] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_87 bl[87] br[87] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_88 bl[88] br[88] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_89 bl[89] br[89] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_90 bl[90] br[90] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_91 bl[91] br[91] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_92 bl[92] br[92] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_93 bl[93] br[93] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_94 bl[94] br[94] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_95 bl[95] br[95] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_96 bl[96] br[96] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_97 bl[97] br[97] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_98 bl[98] br[98] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_99 bl[99] br[99] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_100 bl[100] br[100] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_101 bl[101] br[101] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_102 bl[102] br[102] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_103 bl[103] br[103] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_104 bl[104] br[104] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_105 bl[105] br[105] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_106 bl[106] br[106] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_107 bl[107] br[107] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_108 bl[108] br[108] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_109 bl[109] br[109] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_110 bl[110] br[110] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_111 bl[111] br[111] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_112 bl[112] br[112] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_113 bl[113] br[113] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_114 bl[114] br[114] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_115 bl[115] br[115] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_116 bl[116] br[116] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_117 bl[117] br[117] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_118 bl[118] br[118] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_119 bl[119] br[119] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_120 bl[120] br[120] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_121 bl[121] br[121] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_122 bl[122] br[122] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_123 bl[123] br[123] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_124 bl[124] br[124] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_125 bl[125] br[125] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_126 bl[126] br[126] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_127 bl[127] br[127] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_128 bl[128] br[128] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_129 bl[129] br[129] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_130 bl[130] br[130] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_131 bl[131] br[131] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_132 bl[132] br[132] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_133 bl[133] br[133] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_134 bl[134] br[134] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_135 bl[135] br[135] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_136 bl[136] br[136] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_137 bl[137] br[137] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_138 bl[138] br[138] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_139 bl[139] br[139] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_140 bl[140] br[140] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_141 bl[141] br[141] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_142 bl[142] br[142] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_143 bl[143] br[143] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_144 bl[144] br[144] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_145 bl[145] br[145] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_146 bl[146] br[146] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_147 bl[147] br[147] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_148 bl[148] br[148] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_149 bl[149] br[149] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_150 bl[150] br[150] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_151 bl[151] br[151] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_152 bl[152] br[152] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_153 bl[153] br[153] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_154 bl[154] br[154] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_155 bl[155] br[155] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_156 bl[156] br[156] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_157 bl[157] br[157] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_158 bl[158] br[158] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_159 bl[159] br[159] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_160 bl[160] br[160] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_161 bl[161] br[161] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_162 bl[162] br[162] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_163 bl[163] br[163] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_164 bl[164] br[164] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_165 bl[165] br[165] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_166 bl[166] br[166] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_167 bl[167] br[167] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_168 bl[168] br[168] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_169 bl[169] br[169] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_170 bl[170] br[170] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_171 bl[171] br[171] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_172 bl[172] br[172] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_173 bl[173] br[173] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_174 bl[174] br[174] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_175 bl[175] br[175] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_176 bl[176] br[176] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_177 bl[177] br[177] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_178 bl[178] br[178] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_179 bl[179] br[179] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_180 bl[180] br[180] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_181 bl[181] br[181] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_182 bl[182] br[182] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_183 bl[183] br[183] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_184 bl[184] br[184] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_185 bl[185] br[185] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_186 bl[186] br[186] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_187 bl[187] br[187] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_188 bl[188] br[188] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_189 bl[189] br[189] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_190 bl[190] br[190] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_191 bl[191] br[191] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_192 bl[192] br[192] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_193 bl[193] br[193] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_194 bl[194] br[194] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_195 bl[195] br[195] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_196 bl[196] br[196] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_197 bl[197] br[197] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_198 bl[198] br[198] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_199 bl[199] br[199] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_200 bl[200] br[200] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_201 bl[201] br[201] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_202 bl[202] br[202] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_203 bl[203] br[203] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_204 bl[204] br[204] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_205 bl[205] br[205] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_206 bl[206] br[206] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_207 bl[207] br[207] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_208 bl[208] br[208] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_209 bl[209] br[209] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_210 bl[210] br[210] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_211 bl[211] br[211] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_212 bl[212] br[212] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_213 bl[213] br[213] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_214 bl[214] br[214] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_215 bl[215] br[215] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_216 bl[216] br[216] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_217 bl[217] br[217] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_218 bl[218] br[218] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_219 bl[219] br[219] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_220 bl[220] br[220] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_221 bl[221] br[221] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_222 bl[222] br[222] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_223 bl[223] br[223] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_224 bl[224] br[224] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_225 bl[225] br[225] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_226 bl[226] br[226] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_227 bl[227] br[227] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_228 bl[228] br[228] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_229 bl[229] br[229] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_230 bl[230] br[230] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_231 bl[231] br[231] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_232 bl[232] br[232] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_233 bl[233] br[233] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_234 bl[234] br[234] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_235 bl[235] br[235] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_236 bl[236] br[236] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_237 bl[237] br[237] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_238 bl[238] br[238] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_239 bl[239] br[239] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_240 bl[240] br[240] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_241 bl[241] br[241] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_242 bl[242] br[242] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_243 bl[243] br[243] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_244 bl[244] br[244] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_245 bl[245] br[245] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_246 bl[246] br[246] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_247 bl[247] br[247] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_248 bl[248] br[248] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_249 bl[249] br[249] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_250 bl[250] br[250] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_251 bl[251] br[251] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_252 bl[252] br[252] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_253 bl[253] br[253] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_254 bl[254] br[254] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_255 bl[255] br[255] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_64_0 bl[0] br[0] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_1 bl[1] br[1] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_2 bl[2] br[2] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_3 bl[3] br[3] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_4 bl[4] br[4] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_5 bl[5] br[5] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_6 bl[6] br[6] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_7 bl[7] br[7] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_8 bl[8] br[8] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_9 bl[9] br[9] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_10 bl[10] br[10] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_11 bl[11] br[11] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_12 bl[12] br[12] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_13 bl[13] br[13] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_14 bl[14] br[14] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_15 bl[15] br[15] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_16 bl[16] br[16] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_17 bl[17] br[17] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_18 bl[18] br[18] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_19 bl[19] br[19] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_20 bl[20] br[20] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_21 bl[21] br[21] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_22 bl[22] br[22] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_23 bl[23] br[23] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_24 bl[24] br[24] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_25 bl[25] br[25] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_26 bl[26] br[26] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_27 bl[27] br[27] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_28 bl[28] br[28] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_29 bl[29] br[29] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_30 bl[30] br[30] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_31 bl[31] br[31] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_32 bl[32] br[32] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_33 bl[33] br[33] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_34 bl[34] br[34] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_35 bl[35] br[35] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_36 bl[36] br[36] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_37 bl[37] br[37] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_38 bl[38] br[38] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_39 bl[39] br[39] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_40 bl[40] br[40] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_41 bl[41] br[41] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_42 bl[42] br[42] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_43 bl[43] br[43] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_44 bl[44] br[44] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_45 bl[45] br[45] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_46 bl[46] br[46] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_47 bl[47] br[47] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_48 bl[48] br[48] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_49 bl[49] br[49] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_50 bl[50] br[50] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_51 bl[51] br[51] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_52 bl[52] br[52] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_53 bl[53] br[53] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_54 bl[54] br[54] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_55 bl[55] br[55] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_56 bl[56] br[56] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_57 bl[57] br[57] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_58 bl[58] br[58] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_59 bl[59] br[59] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_60 bl[60] br[60] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_61 bl[61] br[61] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_62 bl[62] br[62] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_63 bl[63] br[63] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_64 bl[64] br[64] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_65 bl[65] br[65] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_66 bl[66] br[66] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_67 bl[67] br[67] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_68 bl[68] br[68] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_69 bl[69] br[69] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_70 bl[70] br[70] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_71 bl[71] br[71] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_72 bl[72] br[72] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_73 bl[73] br[73] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_74 bl[74] br[74] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_75 bl[75] br[75] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_76 bl[76] br[76] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_77 bl[77] br[77] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_78 bl[78] br[78] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_79 bl[79] br[79] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_80 bl[80] br[80] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_81 bl[81] br[81] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_82 bl[82] br[82] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_83 bl[83] br[83] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_84 bl[84] br[84] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_85 bl[85] br[85] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_86 bl[86] br[86] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_87 bl[87] br[87] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_88 bl[88] br[88] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_89 bl[89] br[89] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_90 bl[90] br[90] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_91 bl[91] br[91] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_92 bl[92] br[92] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_93 bl[93] br[93] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_94 bl[94] br[94] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_95 bl[95] br[95] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_96 bl[96] br[96] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_97 bl[97] br[97] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_98 bl[98] br[98] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_99 bl[99] br[99] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_100 bl[100] br[100] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_101 bl[101] br[101] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_102 bl[102] br[102] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_103 bl[103] br[103] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_104 bl[104] br[104] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_105 bl[105] br[105] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_106 bl[106] br[106] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_107 bl[107] br[107] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_108 bl[108] br[108] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_109 bl[109] br[109] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_110 bl[110] br[110] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_111 bl[111] br[111] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_112 bl[112] br[112] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_113 bl[113] br[113] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_114 bl[114] br[114] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_115 bl[115] br[115] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_116 bl[116] br[116] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_117 bl[117] br[117] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_118 bl[118] br[118] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_119 bl[119] br[119] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_120 bl[120] br[120] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_121 bl[121] br[121] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_122 bl[122] br[122] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_123 bl[123] br[123] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_124 bl[124] br[124] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_125 bl[125] br[125] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_126 bl[126] br[126] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_127 bl[127] br[127] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_128 bl[128] br[128] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_129 bl[129] br[129] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_130 bl[130] br[130] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_131 bl[131] br[131] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_132 bl[132] br[132] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_133 bl[133] br[133] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_134 bl[134] br[134] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_135 bl[135] br[135] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_136 bl[136] br[136] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_137 bl[137] br[137] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_138 bl[138] br[138] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_139 bl[139] br[139] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_140 bl[140] br[140] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_141 bl[141] br[141] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_142 bl[142] br[142] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_143 bl[143] br[143] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_144 bl[144] br[144] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_145 bl[145] br[145] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_146 bl[146] br[146] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_147 bl[147] br[147] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_148 bl[148] br[148] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_149 bl[149] br[149] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_150 bl[150] br[150] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_151 bl[151] br[151] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_152 bl[152] br[152] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_153 bl[153] br[153] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_154 bl[154] br[154] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_155 bl[155] br[155] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_156 bl[156] br[156] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_157 bl[157] br[157] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_158 bl[158] br[158] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_159 bl[159] br[159] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_160 bl[160] br[160] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_161 bl[161] br[161] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_162 bl[162] br[162] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_163 bl[163] br[163] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_164 bl[164] br[164] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_165 bl[165] br[165] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_166 bl[166] br[166] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_167 bl[167] br[167] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_168 bl[168] br[168] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_169 bl[169] br[169] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_170 bl[170] br[170] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_171 bl[171] br[171] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_172 bl[172] br[172] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_173 bl[173] br[173] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_174 bl[174] br[174] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_175 bl[175] br[175] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_176 bl[176] br[176] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_177 bl[177] br[177] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_178 bl[178] br[178] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_179 bl[179] br[179] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_180 bl[180] br[180] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_181 bl[181] br[181] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_182 bl[182] br[182] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_183 bl[183] br[183] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_184 bl[184] br[184] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_185 bl[185] br[185] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_186 bl[186] br[186] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_187 bl[187] br[187] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_188 bl[188] br[188] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_189 bl[189] br[189] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_190 bl[190] br[190] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_191 bl[191] br[191] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_192 bl[192] br[192] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_193 bl[193] br[193] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_194 bl[194] br[194] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_195 bl[195] br[195] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_196 bl[196] br[196] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_197 bl[197] br[197] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_198 bl[198] br[198] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_199 bl[199] br[199] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_200 bl[200] br[200] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_201 bl[201] br[201] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_202 bl[202] br[202] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_203 bl[203] br[203] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_204 bl[204] br[204] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_205 bl[205] br[205] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_206 bl[206] br[206] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_207 bl[207] br[207] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_208 bl[208] br[208] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_209 bl[209] br[209] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_210 bl[210] br[210] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_211 bl[211] br[211] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_212 bl[212] br[212] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_213 bl[213] br[213] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_214 bl[214] br[214] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_215 bl[215] br[215] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_216 bl[216] br[216] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_217 bl[217] br[217] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_218 bl[218] br[218] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_219 bl[219] br[219] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_220 bl[220] br[220] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_221 bl[221] br[221] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_222 bl[222] br[222] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_223 bl[223] br[223] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_224 bl[224] br[224] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_225 bl[225] br[225] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_226 bl[226] br[226] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_227 bl[227] br[227] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_228 bl[228] br[228] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_229 bl[229] br[229] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_230 bl[230] br[230] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_231 bl[231] br[231] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_232 bl[232] br[232] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_233 bl[233] br[233] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_234 bl[234] br[234] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_235 bl[235] br[235] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_236 bl[236] br[236] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_237 bl[237] br[237] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_238 bl[238] br[238] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_239 bl[239] br[239] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_240 bl[240] br[240] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_241 bl[241] br[241] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_242 bl[242] br[242] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_243 bl[243] br[243] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_244 bl[244] br[244] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_245 bl[245] br[245] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_246 bl[246] br[246] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_247 bl[247] br[247] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_248 bl[248] br[248] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_249 bl[249] br[249] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_250 bl[250] br[250] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_251 bl[251] br[251] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_252 bl[252] br[252] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_253 bl[253] br[253] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_254 bl[254] br[254] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_255 bl[255] br[255] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_65_0 bl[0] br[0] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_1 bl[1] br[1] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_2 bl[2] br[2] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_3 bl[3] br[3] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_4 bl[4] br[4] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_5 bl[5] br[5] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_6 bl[6] br[6] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_7 bl[7] br[7] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_8 bl[8] br[8] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_9 bl[9] br[9] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_10 bl[10] br[10] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_11 bl[11] br[11] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_12 bl[12] br[12] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_13 bl[13] br[13] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_14 bl[14] br[14] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_15 bl[15] br[15] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_16 bl[16] br[16] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_17 bl[17] br[17] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_18 bl[18] br[18] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_19 bl[19] br[19] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_20 bl[20] br[20] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_21 bl[21] br[21] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_22 bl[22] br[22] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_23 bl[23] br[23] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_24 bl[24] br[24] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_25 bl[25] br[25] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_26 bl[26] br[26] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_27 bl[27] br[27] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_28 bl[28] br[28] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_29 bl[29] br[29] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_30 bl[30] br[30] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_31 bl[31] br[31] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_32 bl[32] br[32] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_33 bl[33] br[33] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_34 bl[34] br[34] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_35 bl[35] br[35] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_36 bl[36] br[36] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_37 bl[37] br[37] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_38 bl[38] br[38] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_39 bl[39] br[39] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_40 bl[40] br[40] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_41 bl[41] br[41] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_42 bl[42] br[42] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_43 bl[43] br[43] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_44 bl[44] br[44] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_45 bl[45] br[45] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_46 bl[46] br[46] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_47 bl[47] br[47] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_48 bl[48] br[48] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_49 bl[49] br[49] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_50 bl[50] br[50] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_51 bl[51] br[51] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_52 bl[52] br[52] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_53 bl[53] br[53] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_54 bl[54] br[54] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_55 bl[55] br[55] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_56 bl[56] br[56] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_57 bl[57] br[57] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_58 bl[58] br[58] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_59 bl[59] br[59] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_60 bl[60] br[60] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_61 bl[61] br[61] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_62 bl[62] br[62] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_63 bl[63] br[63] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_64 bl[64] br[64] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_65 bl[65] br[65] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_66 bl[66] br[66] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_67 bl[67] br[67] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_68 bl[68] br[68] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_69 bl[69] br[69] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_70 bl[70] br[70] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_71 bl[71] br[71] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_72 bl[72] br[72] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_73 bl[73] br[73] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_74 bl[74] br[74] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_75 bl[75] br[75] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_76 bl[76] br[76] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_77 bl[77] br[77] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_78 bl[78] br[78] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_79 bl[79] br[79] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_80 bl[80] br[80] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_81 bl[81] br[81] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_82 bl[82] br[82] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_83 bl[83] br[83] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_84 bl[84] br[84] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_85 bl[85] br[85] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_86 bl[86] br[86] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_87 bl[87] br[87] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_88 bl[88] br[88] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_89 bl[89] br[89] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_90 bl[90] br[90] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_91 bl[91] br[91] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_92 bl[92] br[92] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_93 bl[93] br[93] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_94 bl[94] br[94] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_95 bl[95] br[95] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_96 bl[96] br[96] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_97 bl[97] br[97] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_98 bl[98] br[98] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_99 bl[99] br[99] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_100 bl[100] br[100] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_101 bl[101] br[101] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_102 bl[102] br[102] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_103 bl[103] br[103] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_104 bl[104] br[104] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_105 bl[105] br[105] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_106 bl[106] br[106] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_107 bl[107] br[107] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_108 bl[108] br[108] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_109 bl[109] br[109] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_110 bl[110] br[110] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_111 bl[111] br[111] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_112 bl[112] br[112] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_113 bl[113] br[113] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_114 bl[114] br[114] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_115 bl[115] br[115] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_116 bl[116] br[116] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_117 bl[117] br[117] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_118 bl[118] br[118] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_119 bl[119] br[119] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_120 bl[120] br[120] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_121 bl[121] br[121] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_122 bl[122] br[122] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_123 bl[123] br[123] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_124 bl[124] br[124] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_125 bl[125] br[125] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_126 bl[126] br[126] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_127 bl[127] br[127] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_128 bl[128] br[128] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_129 bl[129] br[129] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_130 bl[130] br[130] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_131 bl[131] br[131] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_132 bl[132] br[132] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_133 bl[133] br[133] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_134 bl[134] br[134] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_135 bl[135] br[135] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_136 bl[136] br[136] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_137 bl[137] br[137] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_138 bl[138] br[138] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_139 bl[139] br[139] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_140 bl[140] br[140] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_141 bl[141] br[141] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_142 bl[142] br[142] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_143 bl[143] br[143] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_144 bl[144] br[144] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_145 bl[145] br[145] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_146 bl[146] br[146] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_147 bl[147] br[147] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_148 bl[148] br[148] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_149 bl[149] br[149] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_150 bl[150] br[150] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_151 bl[151] br[151] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_152 bl[152] br[152] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_153 bl[153] br[153] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_154 bl[154] br[154] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_155 bl[155] br[155] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_156 bl[156] br[156] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_157 bl[157] br[157] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_158 bl[158] br[158] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_159 bl[159] br[159] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_160 bl[160] br[160] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_161 bl[161] br[161] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_162 bl[162] br[162] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_163 bl[163] br[163] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_164 bl[164] br[164] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_165 bl[165] br[165] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_166 bl[166] br[166] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_167 bl[167] br[167] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_168 bl[168] br[168] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_169 bl[169] br[169] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_170 bl[170] br[170] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_171 bl[171] br[171] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_172 bl[172] br[172] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_173 bl[173] br[173] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_174 bl[174] br[174] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_175 bl[175] br[175] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_176 bl[176] br[176] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_177 bl[177] br[177] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_178 bl[178] br[178] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_179 bl[179] br[179] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_180 bl[180] br[180] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_181 bl[181] br[181] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_182 bl[182] br[182] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_183 bl[183] br[183] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_184 bl[184] br[184] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_185 bl[185] br[185] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_186 bl[186] br[186] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_187 bl[187] br[187] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_188 bl[188] br[188] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_189 bl[189] br[189] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_190 bl[190] br[190] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_191 bl[191] br[191] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_192 bl[192] br[192] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_193 bl[193] br[193] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_194 bl[194] br[194] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_195 bl[195] br[195] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_196 bl[196] br[196] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_197 bl[197] br[197] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_198 bl[198] br[198] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_199 bl[199] br[199] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_200 bl[200] br[200] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_201 bl[201] br[201] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_202 bl[202] br[202] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_203 bl[203] br[203] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_204 bl[204] br[204] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_205 bl[205] br[205] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_206 bl[206] br[206] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_207 bl[207] br[207] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_208 bl[208] br[208] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_209 bl[209] br[209] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_210 bl[210] br[210] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_211 bl[211] br[211] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_212 bl[212] br[212] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_213 bl[213] br[213] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_214 bl[214] br[214] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_215 bl[215] br[215] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_216 bl[216] br[216] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_217 bl[217] br[217] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_218 bl[218] br[218] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_219 bl[219] br[219] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_220 bl[220] br[220] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_221 bl[221] br[221] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_222 bl[222] br[222] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_223 bl[223] br[223] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_224 bl[224] br[224] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_225 bl[225] br[225] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_226 bl[226] br[226] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_227 bl[227] br[227] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_228 bl[228] br[228] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_229 bl[229] br[229] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_230 bl[230] br[230] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_231 bl[231] br[231] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_232 bl[232] br[232] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_233 bl[233] br[233] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_234 bl[234] br[234] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_235 bl[235] br[235] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_236 bl[236] br[236] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_237 bl[237] br[237] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_238 bl[238] br[238] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_239 bl[239] br[239] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_240 bl[240] br[240] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_241 bl[241] br[241] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_242 bl[242] br[242] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_243 bl[243] br[243] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_244 bl[244] br[244] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_245 bl[245] br[245] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_246 bl[246] br[246] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_247 bl[247] br[247] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_248 bl[248] br[248] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_249 bl[249] br[249] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_250 bl[250] br[250] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_251 bl[251] br[251] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_252 bl[252] br[252] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_253 bl[253] br[253] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_254 bl[254] br[254] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_255 bl[255] br[255] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_66_0 bl[0] br[0] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_1 bl[1] br[1] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_2 bl[2] br[2] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_3 bl[3] br[3] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_4 bl[4] br[4] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_5 bl[5] br[5] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_6 bl[6] br[6] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_7 bl[7] br[7] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_8 bl[8] br[8] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_9 bl[9] br[9] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_10 bl[10] br[10] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_11 bl[11] br[11] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_12 bl[12] br[12] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_13 bl[13] br[13] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_14 bl[14] br[14] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_15 bl[15] br[15] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_16 bl[16] br[16] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_17 bl[17] br[17] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_18 bl[18] br[18] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_19 bl[19] br[19] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_20 bl[20] br[20] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_21 bl[21] br[21] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_22 bl[22] br[22] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_23 bl[23] br[23] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_24 bl[24] br[24] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_25 bl[25] br[25] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_26 bl[26] br[26] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_27 bl[27] br[27] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_28 bl[28] br[28] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_29 bl[29] br[29] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_30 bl[30] br[30] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_31 bl[31] br[31] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_32 bl[32] br[32] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_33 bl[33] br[33] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_34 bl[34] br[34] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_35 bl[35] br[35] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_36 bl[36] br[36] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_37 bl[37] br[37] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_38 bl[38] br[38] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_39 bl[39] br[39] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_40 bl[40] br[40] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_41 bl[41] br[41] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_42 bl[42] br[42] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_43 bl[43] br[43] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_44 bl[44] br[44] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_45 bl[45] br[45] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_46 bl[46] br[46] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_47 bl[47] br[47] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_48 bl[48] br[48] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_49 bl[49] br[49] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_50 bl[50] br[50] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_51 bl[51] br[51] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_52 bl[52] br[52] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_53 bl[53] br[53] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_54 bl[54] br[54] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_55 bl[55] br[55] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_56 bl[56] br[56] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_57 bl[57] br[57] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_58 bl[58] br[58] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_59 bl[59] br[59] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_60 bl[60] br[60] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_61 bl[61] br[61] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_62 bl[62] br[62] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_63 bl[63] br[63] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_64 bl[64] br[64] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_65 bl[65] br[65] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_66 bl[66] br[66] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_67 bl[67] br[67] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_68 bl[68] br[68] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_69 bl[69] br[69] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_70 bl[70] br[70] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_71 bl[71] br[71] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_72 bl[72] br[72] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_73 bl[73] br[73] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_74 bl[74] br[74] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_75 bl[75] br[75] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_76 bl[76] br[76] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_77 bl[77] br[77] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_78 bl[78] br[78] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_79 bl[79] br[79] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_80 bl[80] br[80] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_81 bl[81] br[81] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_82 bl[82] br[82] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_83 bl[83] br[83] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_84 bl[84] br[84] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_85 bl[85] br[85] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_86 bl[86] br[86] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_87 bl[87] br[87] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_88 bl[88] br[88] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_89 bl[89] br[89] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_90 bl[90] br[90] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_91 bl[91] br[91] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_92 bl[92] br[92] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_93 bl[93] br[93] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_94 bl[94] br[94] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_95 bl[95] br[95] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_96 bl[96] br[96] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_97 bl[97] br[97] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_98 bl[98] br[98] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_99 bl[99] br[99] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_100 bl[100] br[100] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_101 bl[101] br[101] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_102 bl[102] br[102] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_103 bl[103] br[103] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_104 bl[104] br[104] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_105 bl[105] br[105] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_106 bl[106] br[106] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_107 bl[107] br[107] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_108 bl[108] br[108] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_109 bl[109] br[109] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_110 bl[110] br[110] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_111 bl[111] br[111] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_112 bl[112] br[112] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_113 bl[113] br[113] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_114 bl[114] br[114] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_115 bl[115] br[115] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_116 bl[116] br[116] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_117 bl[117] br[117] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_118 bl[118] br[118] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_119 bl[119] br[119] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_120 bl[120] br[120] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_121 bl[121] br[121] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_122 bl[122] br[122] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_123 bl[123] br[123] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_124 bl[124] br[124] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_125 bl[125] br[125] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_126 bl[126] br[126] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_127 bl[127] br[127] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_128 bl[128] br[128] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_129 bl[129] br[129] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_130 bl[130] br[130] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_131 bl[131] br[131] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_132 bl[132] br[132] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_133 bl[133] br[133] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_134 bl[134] br[134] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_135 bl[135] br[135] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_136 bl[136] br[136] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_137 bl[137] br[137] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_138 bl[138] br[138] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_139 bl[139] br[139] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_140 bl[140] br[140] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_141 bl[141] br[141] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_142 bl[142] br[142] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_143 bl[143] br[143] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_144 bl[144] br[144] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_145 bl[145] br[145] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_146 bl[146] br[146] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_147 bl[147] br[147] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_148 bl[148] br[148] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_149 bl[149] br[149] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_150 bl[150] br[150] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_151 bl[151] br[151] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_152 bl[152] br[152] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_153 bl[153] br[153] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_154 bl[154] br[154] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_155 bl[155] br[155] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_156 bl[156] br[156] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_157 bl[157] br[157] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_158 bl[158] br[158] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_159 bl[159] br[159] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_160 bl[160] br[160] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_161 bl[161] br[161] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_162 bl[162] br[162] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_163 bl[163] br[163] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_164 bl[164] br[164] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_165 bl[165] br[165] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_166 bl[166] br[166] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_167 bl[167] br[167] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_168 bl[168] br[168] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_169 bl[169] br[169] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_170 bl[170] br[170] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_171 bl[171] br[171] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_172 bl[172] br[172] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_173 bl[173] br[173] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_174 bl[174] br[174] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_175 bl[175] br[175] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_176 bl[176] br[176] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_177 bl[177] br[177] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_178 bl[178] br[178] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_179 bl[179] br[179] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_180 bl[180] br[180] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_181 bl[181] br[181] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_182 bl[182] br[182] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_183 bl[183] br[183] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_184 bl[184] br[184] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_185 bl[185] br[185] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_186 bl[186] br[186] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_187 bl[187] br[187] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_188 bl[188] br[188] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_189 bl[189] br[189] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_190 bl[190] br[190] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_191 bl[191] br[191] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_192 bl[192] br[192] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_193 bl[193] br[193] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_194 bl[194] br[194] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_195 bl[195] br[195] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_196 bl[196] br[196] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_197 bl[197] br[197] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_198 bl[198] br[198] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_199 bl[199] br[199] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_200 bl[200] br[200] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_201 bl[201] br[201] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_202 bl[202] br[202] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_203 bl[203] br[203] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_204 bl[204] br[204] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_205 bl[205] br[205] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_206 bl[206] br[206] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_207 bl[207] br[207] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_208 bl[208] br[208] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_209 bl[209] br[209] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_210 bl[210] br[210] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_211 bl[211] br[211] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_212 bl[212] br[212] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_213 bl[213] br[213] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_214 bl[214] br[214] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_215 bl[215] br[215] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_216 bl[216] br[216] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_217 bl[217] br[217] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_218 bl[218] br[218] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_219 bl[219] br[219] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_220 bl[220] br[220] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_221 bl[221] br[221] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_222 bl[222] br[222] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_223 bl[223] br[223] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_224 bl[224] br[224] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_225 bl[225] br[225] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_226 bl[226] br[226] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_227 bl[227] br[227] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_228 bl[228] br[228] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_229 bl[229] br[229] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_230 bl[230] br[230] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_231 bl[231] br[231] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_232 bl[232] br[232] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_233 bl[233] br[233] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_234 bl[234] br[234] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_235 bl[235] br[235] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_236 bl[236] br[236] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_237 bl[237] br[237] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_238 bl[238] br[238] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_239 bl[239] br[239] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_240 bl[240] br[240] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_241 bl[241] br[241] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_242 bl[242] br[242] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_243 bl[243] br[243] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_244 bl[244] br[244] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_245 bl[245] br[245] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_246 bl[246] br[246] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_247 bl[247] br[247] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_248 bl[248] br[248] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_249 bl[249] br[249] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_250 bl[250] br[250] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_251 bl[251] br[251] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_252 bl[252] br[252] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_253 bl[253] br[253] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_254 bl[254] br[254] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_255 bl[255] br[255] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_67_0 bl[0] br[0] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_1 bl[1] br[1] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_2 bl[2] br[2] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_3 bl[3] br[3] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_4 bl[4] br[4] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_5 bl[5] br[5] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_6 bl[6] br[6] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_7 bl[7] br[7] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_8 bl[8] br[8] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_9 bl[9] br[9] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_10 bl[10] br[10] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_11 bl[11] br[11] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_12 bl[12] br[12] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_13 bl[13] br[13] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_14 bl[14] br[14] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_15 bl[15] br[15] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_16 bl[16] br[16] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_17 bl[17] br[17] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_18 bl[18] br[18] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_19 bl[19] br[19] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_20 bl[20] br[20] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_21 bl[21] br[21] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_22 bl[22] br[22] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_23 bl[23] br[23] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_24 bl[24] br[24] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_25 bl[25] br[25] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_26 bl[26] br[26] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_27 bl[27] br[27] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_28 bl[28] br[28] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_29 bl[29] br[29] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_30 bl[30] br[30] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_31 bl[31] br[31] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_32 bl[32] br[32] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_33 bl[33] br[33] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_34 bl[34] br[34] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_35 bl[35] br[35] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_36 bl[36] br[36] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_37 bl[37] br[37] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_38 bl[38] br[38] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_39 bl[39] br[39] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_40 bl[40] br[40] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_41 bl[41] br[41] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_42 bl[42] br[42] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_43 bl[43] br[43] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_44 bl[44] br[44] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_45 bl[45] br[45] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_46 bl[46] br[46] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_47 bl[47] br[47] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_48 bl[48] br[48] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_49 bl[49] br[49] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_50 bl[50] br[50] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_51 bl[51] br[51] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_52 bl[52] br[52] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_53 bl[53] br[53] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_54 bl[54] br[54] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_55 bl[55] br[55] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_56 bl[56] br[56] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_57 bl[57] br[57] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_58 bl[58] br[58] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_59 bl[59] br[59] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_60 bl[60] br[60] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_61 bl[61] br[61] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_62 bl[62] br[62] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_63 bl[63] br[63] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_64 bl[64] br[64] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_65 bl[65] br[65] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_66 bl[66] br[66] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_67 bl[67] br[67] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_68 bl[68] br[68] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_69 bl[69] br[69] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_70 bl[70] br[70] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_71 bl[71] br[71] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_72 bl[72] br[72] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_73 bl[73] br[73] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_74 bl[74] br[74] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_75 bl[75] br[75] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_76 bl[76] br[76] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_77 bl[77] br[77] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_78 bl[78] br[78] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_79 bl[79] br[79] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_80 bl[80] br[80] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_81 bl[81] br[81] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_82 bl[82] br[82] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_83 bl[83] br[83] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_84 bl[84] br[84] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_85 bl[85] br[85] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_86 bl[86] br[86] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_87 bl[87] br[87] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_88 bl[88] br[88] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_89 bl[89] br[89] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_90 bl[90] br[90] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_91 bl[91] br[91] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_92 bl[92] br[92] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_93 bl[93] br[93] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_94 bl[94] br[94] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_95 bl[95] br[95] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_96 bl[96] br[96] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_97 bl[97] br[97] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_98 bl[98] br[98] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_99 bl[99] br[99] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_100 bl[100] br[100] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_101 bl[101] br[101] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_102 bl[102] br[102] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_103 bl[103] br[103] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_104 bl[104] br[104] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_105 bl[105] br[105] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_106 bl[106] br[106] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_107 bl[107] br[107] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_108 bl[108] br[108] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_109 bl[109] br[109] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_110 bl[110] br[110] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_111 bl[111] br[111] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_112 bl[112] br[112] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_113 bl[113] br[113] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_114 bl[114] br[114] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_115 bl[115] br[115] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_116 bl[116] br[116] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_117 bl[117] br[117] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_118 bl[118] br[118] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_119 bl[119] br[119] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_120 bl[120] br[120] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_121 bl[121] br[121] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_122 bl[122] br[122] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_123 bl[123] br[123] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_124 bl[124] br[124] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_125 bl[125] br[125] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_126 bl[126] br[126] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_127 bl[127] br[127] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_128 bl[128] br[128] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_129 bl[129] br[129] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_130 bl[130] br[130] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_131 bl[131] br[131] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_132 bl[132] br[132] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_133 bl[133] br[133] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_134 bl[134] br[134] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_135 bl[135] br[135] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_136 bl[136] br[136] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_137 bl[137] br[137] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_138 bl[138] br[138] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_139 bl[139] br[139] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_140 bl[140] br[140] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_141 bl[141] br[141] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_142 bl[142] br[142] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_143 bl[143] br[143] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_144 bl[144] br[144] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_145 bl[145] br[145] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_146 bl[146] br[146] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_147 bl[147] br[147] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_148 bl[148] br[148] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_149 bl[149] br[149] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_150 bl[150] br[150] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_151 bl[151] br[151] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_152 bl[152] br[152] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_153 bl[153] br[153] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_154 bl[154] br[154] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_155 bl[155] br[155] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_156 bl[156] br[156] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_157 bl[157] br[157] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_158 bl[158] br[158] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_159 bl[159] br[159] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_160 bl[160] br[160] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_161 bl[161] br[161] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_162 bl[162] br[162] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_163 bl[163] br[163] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_164 bl[164] br[164] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_165 bl[165] br[165] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_166 bl[166] br[166] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_167 bl[167] br[167] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_168 bl[168] br[168] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_169 bl[169] br[169] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_170 bl[170] br[170] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_171 bl[171] br[171] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_172 bl[172] br[172] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_173 bl[173] br[173] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_174 bl[174] br[174] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_175 bl[175] br[175] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_176 bl[176] br[176] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_177 bl[177] br[177] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_178 bl[178] br[178] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_179 bl[179] br[179] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_180 bl[180] br[180] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_181 bl[181] br[181] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_182 bl[182] br[182] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_183 bl[183] br[183] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_184 bl[184] br[184] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_185 bl[185] br[185] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_186 bl[186] br[186] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_187 bl[187] br[187] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_188 bl[188] br[188] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_189 bl[189] br[189] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_190 bl[190] br[190] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_191 bl[191] br[191] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_192 bl[192] br[192] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_193 bl[193] br[193] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_194 bl[194] br[194] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_195 bl[195] br[195] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_196 bl[196] br[196] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_197 bl[197] br[197] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_198 bl[198] br[198] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_199 bl[199] br[199] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_200 bl[200] br[200] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_201 bl[201] br[201] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_202 bl[202] br[202] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_203 bl[203] br[203] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_204 bl[204] br[204] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_205 bl[205] br[205] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_206 bl[206] br[206] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_207 bl[207] br[207] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_208 bl[208] br[208] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_209 bl[209] br[209] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_210 bl[210] br[210] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_211 bl[211] br[211] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_212 bl[212] br[212] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_213 bl[213] br[213] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_214 bl[214] br[214] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_215 bl[215] br[215] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_216 bl[216] br[216] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_217 bl[217] br[217] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_218 bl[218] br[218] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_219 bl[219] br[219] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_220 bl[220] br[220] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_221 bl[221] br[221] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_222 bl[222] br[222] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_223 bl[223] br[223] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_224 bl[224] br[224] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_225 bl[225] br[225] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_226 bl[226] br[226] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_227 bl[227] br[227] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_228 bl[228] br[228] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_229 bl[229] br[229] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_230 bl[230] br[230] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_231 bl[231] br[231] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_232 bl[232] br[232] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_233 bl[233] br[233] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_234 bl[234] br[234] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_235 bl[235] br[235] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_236 bl[236] br[236] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_237 bl[237] br[237] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_238 bl[238] br[238] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_239 bl[239] br[239] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_240 bl[240] br[240] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_241 bl[241] br[241] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_242 bl[242] br[242] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_243 bl[243] br[243] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_244 bl[244] br[244] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_245 bl[245] br[245] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_246 bl[246] br[246] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_247 bl[247] br[247] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_248 bl[248] br[248] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_249 bl[249] br[249] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_250 bl[250] br[250] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_251 bl[251] br[251] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_252 bl[252] br[252] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_253 bl[253] br[253] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_254 bl[254] br[254] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_255 bl[255] br[255] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_68_0 bl[0] br[0] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_1 bl[1] br[1] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_2 bl[2] br[2] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_3 bl[3] br[3] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_4 bl[4] br[4] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_5 bl[5] br[5] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_6 bl[6] br[6] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_7 bl[7] br[7] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_8 bl[8] br[8] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_9 bl[9] br[9] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_10 bl[10] br[10] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_11 bl[11] br[11] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_12 bl[12] br[12] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_13 bl[13] br[13] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_14 bl[14] br[14] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_15 bl[15] br[15] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_16 bl[16] br[16] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_17 bl[17] br[17] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_18 bl[18] br[18] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_19 bl[19] br[19] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_20 bl[20] br[20] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_21 bl[21] br[21] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_22 bl[22] br[22] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_23 bl[23] br[23] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_24 bl[24] br[24] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_25 bl[25] br[25] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_26 bl[26] br[26] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_27 bl[27] br[27] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_28 bl[28] br[28] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_29 bl[29] br[29] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_30 bl[30] br[30] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_31 bl[31] br[31] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_32 bl[32] br[32] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_33 bl[33] br[33] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_34 bl[34] br[34] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_35 bl[35] br[35] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_36 bl[36] br[36] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_37 bl[37] br[37] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_38 bl[38] br[38] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_39 bl[39] br[39] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_40 bl[40] br[40] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_41 bl[41] br[41] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_42 bl[42] br[42] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_43 bl[43] br[43] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_44 bl[44] br[44] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_45 bl[45] br[45] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_46 bl[46] br[46] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_47 bl[47] br[47] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_48 bl[48] br[48] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_49 bl[49] br[49] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_50 bl[50] br[50] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_51 bl[51] br[51] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_52 bl[52] br[52] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_53 bl[53] br[53] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_54 bl[54] br[54] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_55 bl[55] br[55] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_56 bl[56] br[56] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_57 bl[57] br[57] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_58 bl[58] br[58] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_59 bl[59] br[59] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_60 bl[60] br[60] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_61 bl[61] br[61] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_62 bl[62] br[62] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_63 bl[63] br[63] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_64 bl[64] br[64] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_65 bl[65] br[65] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_66 bl[66] br[66] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_67 bl[67] br[67] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_68 bl[68] br[68] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_69 bl[69] br[69] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_70 bl[70] br[70] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_71 bl[71] br[71] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_72 bl[72] br[72] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_73 bl[73] br[73] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_74 bl[74] br[74] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_75 bl[75] br[75] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_76 bl[76] br[76] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_77 bl[77] br[77] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_78 bl[78] br[78] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_79 bl[79] br[79] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_80 bl[80] br[80] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_81 bl[81] br[81] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_82 bl[82] br[82] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_83 bl[83] br[83] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_84 bl[84] br[84] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_85 bl[85] br[85] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_86 bl[86] br[86] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_87 bl[87] br[87] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_88 bl[88] br[88] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_89 bl[89] br[89] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_90 bl[90] br[90] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_91 bl[91] br[91] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_92 bl[92] br[92] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_93 bl[93] br[93] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_94 bl[94] br[94] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_95 bl[95] br[95] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_96 bl[96] br[96] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_97 bl[97] br[97] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_98 bl[98] br[98] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_99 bl[99] br[99] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_100 bl[100] br[100] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_101 bl[101] br[101] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_102 bl[102] br[102] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_103 bl[103] br[103] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_104 bl[104] br[104] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_105 bl[105] br[105] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_106 bl[106] br[106] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_107 bl[107] br[107] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_108 bl[108] br[108] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_109 bl[109] br[109] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_110 bl[110] br[110] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_111 bl[111] br[111] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_112 bl[112] br[112] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_113 bl[113] br[113] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_114 bl[114] br[114] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_115 bl[115] br[115] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_116 bl[116] br[116] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_117 bl[117] br[117] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_118 bl[118] br[118] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_119 bl[119] br[119] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_120 bl[120] br[120] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_121 bl[121] br[121] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_122 bl[122] br[122] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_123 bl[123] br[123] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_124 bl[124] br[124] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_125 bl[125] br[125] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_126 bl[126] br[126] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_127 bl[127] br[127] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_128 bl[128] br[128] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_129 bl[129] br[129] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_130 bl[130] br[130] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_131 bl[131] br[131] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_132 bl[132] br[132] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_133 bl[133] br[133] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_134 bl[134] br[134] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_135 bl[135] br[135] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_136 bl[136] br[136] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_137 bl[137] br[137] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_138 bl[138] br[138] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_139 bl[139] br[139] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_140 bl[140] br[140] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_141 bl[141] br[141] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_142 bl[142] br[142] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_143 bl[143] br[143] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_144 bl[144] br[144] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_145 bl[145] br[145] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_146 bl[146] br[146] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_147 bl[147] br[147] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_148 bl[148] br[148] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_149 bl[149] br[149] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_150 bl[150] br[150] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_151 bl[151] br[151] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_152 bl[152] br[152] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_153 bl[153] br[153] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_154 bl[154] br[154] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_155 bl[155] br[155] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_156 bl[156] br[156] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_157 bl[157] br[157] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_158 bl[158] br[158] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_159 bl[159] br[159] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_160 bl[160] br[160] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_161 bl[161] br[161] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_162 bl[162] br[162] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_163 bl[163] br[163] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_164 bl[164] br[164] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_165 bl[165] br[165] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_166 bl[166] br[166] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_167 bl[167] br[167] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_168 bl[168] br[168] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_169 bl[169] br[169] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_170 bl[170] br[170] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_171 bl[171] br[171] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_172 bl[172] br[172] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_173 bl[173] br[173] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_174 bl[174] br[174] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_175 bl[175] br[175] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_176 bl[176] br[176] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_177 bl[177] br[177] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_178 bl[178] br[178] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_179 bl[179] br[179] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_180 bl[180] br[180] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_181 bl[181] br[181] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_182 bl[182] br[182] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_183 bl[183] br[183] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_184 bl[184] br[184] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_185 bl[185] br[185] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_186 bl[186] br[186] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_187 bl[187] br[187] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_188 bl[188] br[188] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_189 bl[189] br[189] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_190 bl[190] br[190] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_191 bl[191] br[191] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_192 bl[192] br[192] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_193 bl[193] br[193] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_194 bl[194] br[194] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_195 bl[195] br[195] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_196 bl[196] br[196] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_197 bl[197] br[197] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_198 bl[198] br[198] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_199 bl[199] br[199] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_200 bl[200] br[200] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_201 bl[201] br[201] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_202 bl[202] br[202] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_203 bl[203] br[203] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_204 bl[204] br[204] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_205 bl[205] br[205] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_206 bl[206] br[206] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_207 bl[207] br[207] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_208 bl[208] br[208] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_209 bl[209] br[209] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_210 bl[210] br[210] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_211 bl[211] br[211] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_212 bl[212] br[212] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_213 bl[213] br[213] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_214 bl[214] br[214] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_215 bl[215] br[215] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_216 bl[216] br[216] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_217 bl[217] br[217] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_218 bl[218] br[218] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_219 bl[219] br[219] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_220 bl[220] br[220] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_221 bl[221] br[221] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_222 bl[222] br[222] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_223 bl[223] br[223] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_224 bl[224] br[224] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_225 bl[225] br[225] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_226 bl[226] br[226] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_227 bl[227] br[227] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_228 bl[228] br[228] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_229 bl[229] br[229] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_230 bl[230] br[230] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_231 bl[231] br[231] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_232 bl[232] br[232] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_233 bl[233] br[233] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_234 bl[234] br[234] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_235 bl[235] br[235] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_236 bl[236] br[236] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_237 bl[237] br[237] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_238 bl[238] br[238] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_239 bl[239] br[239] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_240 bl[240] br[240] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_241 bl[241] br[241] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_242 bl[242] br[242] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_243 bl[243] br[243] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_244 bl[244] br[244] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_245 bl[245] br[245] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_246 bl[246] br[246] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_247 bl[247] br[247] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_248 bl[248] br[248] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_249 bl[249] br[249] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_250 bl[250] br[250] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_251 bl[251] br[251] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_252 bl[252] br[252] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_253 bl[253] br[253] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_254 bl[254] br[254] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_255 bl[255] br[255] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_69_0 bl[0] br[0] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_1 bl[1] br[1] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_2 bl[2] br[2] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_3 bl[3] br[3] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_4 bl[4] br[4] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_5 bl[5] br[5] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_6 bl[6] br[6] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_7 bl[7] br[7] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_8 bl[8] br[8] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_9 bl[9] br[9] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_10 bl[10] br[10] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_11 bl[11] br[11] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_12 bl[12] br[12] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_13 bl[13] br[13] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_14 bl[14] br[14] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_15 bl[15] br[15] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_16 bl[16] br[16] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_17 bl[17] br[17] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_18 bl[18] br[18] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_19 bl[19] br[19] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_20 bl[20] br[20] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_21 bl[21] br[21] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_22 bl[22] br[22] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_23 bl[23] br[23] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_24 bl[24] br[24] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_25 bl[25] br[25] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_26 bl[26] br[26] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_27 bl[27] br[27] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_28 bl[28] br[28] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_29 bl[29] br[29] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_30 bl[30] br[30] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_31 bl[31] br[31] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_32 bl[32] br[32] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_33 bl[33] br[33] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_34 bl[34] br[34] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_35 bl[35] br[35] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_36 bl[36] br[36] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_37 bl[37] br[37] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_38 bl[38] br[38] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_39 bl[39] br[39] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_40 bl[40] br[40] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_41 bl[41] br[41] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_42 bl[42] br[42] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_43 bl[43] br[43] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_44 bl[44] br[44] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_45 bl[45] br[45] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_46 bl[46] br[46] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_47 bl[47] br[47] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_48 bl[48] br[48] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_49 bl[49] br[49] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_50 bl[50] br[50] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_51 bl[51] br[51] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_52 bl[52] br[52] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_53 bl[53] br[53] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_54 bl[54] br[54] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_55 bl[55] br[55] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_56 bl[56] br[56] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_57 bl[57] br[57] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_58 bl[58] br[58] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_59 bl[59] br[59] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_60 bl[60] br[60] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_61 bl[61] br[61] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_62 bl[62] br[62] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_63 bl[63] br[63] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_64 bl[64] br[64] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_65 bl[65] br[65] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_66 bl[66] br[66] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_67 bl[67] br[67] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_68 bl[68] br[68] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_69 bl[69] br[69] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_70 bl[70] br[70] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_71 bl[71] br[71] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_72 bl[72] br[72] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_73 bl[73] br[73] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_74 bl[74] br[74] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_75 bl[75] br[75] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_76 bl[76] br[76] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_77 bl[77] br[77] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_78 bl[78] br[78] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_79 bl[79] br[79] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_80 bl[80] br[80] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_81 bl[81] br[81] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_82 bl[82] br[82] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_83 bl[83] br[83] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_84 bl[84] br[84] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_85 bl[85] br[85] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_86 bl[86] br[86] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_87 bl[87] br[87] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_88 bl[88] br[88] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_89 bl[89] br[89] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_90 bl[90] br[90] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_91 bl[91] br[91] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_92 bl[92] br[92] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_93 bl[93] br[93] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_94 bl[94] br[94] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_95 bl[95] br[95] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_96 bl[96] br[96] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_97 bl[97] br[97] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_98 bl[98] br[98] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_99 bl[99] br[99] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_100 bl[100] br[100] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_101 bl[101] br[101] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_102 bl[102] br[102] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_103 bl[103] br[103] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_104 bl[104] br[104] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_105 bl[105] br[105] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_106 bl[106] br[106] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_107 bl[107] br[107] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_108 bl[108] br[108] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_109 bl[109] br[109] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_110 bl[110] br[110] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_111 bl[111] br[111] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_112 bl[112] br[112] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_113 bl[113] br[113] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_114 bl[114] br[114] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_115 bl[115] br[115] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_116 bl[116] br[116] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_117 bl[117] br[117] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_118 bl[118] br[118] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_119 bl[119] br[119] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_120 bl[120] br[120] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_121 bl[121] br[121] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_122 bl[122] br[122] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_123 bl[123] br[123] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_124 bl[124] br[124] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_125 bl[125] br[125] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_126 bl[126] br[126] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_127 bl[127] br[127] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_128 bl[128] br[128] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_129 bl[129] br[129] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_130 bl[130] br[130] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_131 bl[131] br[131] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_132 bl[132] br[132] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_133 bl[133] br[133] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_134 bl[134] br[134] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_135 bl[135] br[135] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_136 bl[136] br[136] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_137 bl[137] br[137] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_138 bl[138] br[138] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_139 bl[139] br[139] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_140 bl[140] br[140] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_141 bl[141] br[141] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_142 bl[142] br[142] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_143 bl[143] br[143] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_144 bl[144] br[144] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_145 bl[145] br[145] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_146 bl[146] br[146] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_147 bl[147] br[147] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_148 bl[148] br[148] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_149 bl[149] br[149] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_150 bl[150] br[150] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_151 bl[151] br[151] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_152 bl[152] br[152] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_153 bl[153] br[153] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_154 bl[154] br[154] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_155 bl[155] br[155] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_156 bl[156] br[156] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_157 bl[157] br[157] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_158 bl[158] br[158] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_159 bl[159] br[159] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_160 bl[160] br[160] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_161 bl[161] br[161] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_162 bl[162] br[162] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_163 bl[163] br[163] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_164 bl[164] br[164] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_165 bl[165] br[165] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_166 bl[166] br[166] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_167 bl[167] br[167] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_168 bl[168] br[168] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_169 bl[169] br[169] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_170 bl[170] br[170] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_171 bl[171] br[171] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_172 bl[172] br[172] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_173 bl[173] br[173] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_174 bl[174] br[174] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_175 bl[175] br[175] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_176 bl[176] br[176] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_177 bl[177] br[177] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_178 bl[178] br[178] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_179 bl[179] br[179] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_180 bl[180] br[180] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_181 bl[181] br[181] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_182 bl[182] br[182] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_183 bl[183] br[183] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_184 bl[184] br[184] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_185 bl[185] br[185] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_186 bl[186] br[186] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_187 bl[187] br[187] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_188 bl[188] br[188] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_189 bl[189] br[189] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_190 bl[190] br[190] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_191 bl[191] br[191] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_192 bl[192] br[192] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_193 bl[193] br[193] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_194 bl[194] br[194] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_195 bl[195] br[195] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_196 bl[196] br[196] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_197 bl[197] br[197] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_198 bl[198] br[198] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_199 bl[199] br[199] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_200 bl[200] br[200] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_201 bl[201] br[201] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_202 bl[202] br[202] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_203 bl[203] br[203] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_204 bl[204] br[204] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_205 bl[205] br[205] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_206 bl[206] br[206] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_207 bl[207] br[207] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_208 bl[208] br[208] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_209 bl[209] br[209] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_210 bl[210] br[210] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_211 bl[211] br[211] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_212 bl[212] br[212] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_213 bl[213] br[213] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_214 bl[214] br[214] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_215 bl[215] br[215] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_216 bl[216] br[216] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_217 bl[217] br[217] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_218 bl[218] br[218] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_219 bl[219] br[219] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_220 bl[220] br[220] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_221 bl[221] br[221] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_222 bl[222] br[222] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_223 bl[223] br[223] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_224 bl[224] br[224] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_225 bl[225] br[225] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_226 bl[226] br[226] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_227 bl[227] br[227] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_228 bl[228] br[228] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_229 bl[229] br[229] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_230 bl[230] br[230] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_231 bl[231] br[231] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_232 bl[232] br[232] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_233 bl[233] br[233] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_234 bl[234] br[234] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_235 bl[235] br[235] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_236 bl[236] br[236] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_237 bl[237] br[237] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_238 bl[238] br[238] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_239 bl[239] br[239] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_240 bl[240] br[240] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_241 bl[241] br[241] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_242 bl[242] br[242] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_243 bl[243] br[243] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_244 bl[244] br[244] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_245 bl[245] br[245] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_246 bl[246] br[246] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_247 bl[247] br[247] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_248 bl[248] br[248] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_249 bl[249] br[249] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_250 bl[250] br[250] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_251 bl[251] br[251] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_252 bl[252] br[252] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_253 bl[253] br[253] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_254 bl[254] br[254] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_255 bl[255] br[255] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_70_0 bl[0] br[0] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_1 bl[1] br[1] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_2 bl[2] br[2] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_3 bl[3] br[3] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_4 bl[4] br[4] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_5 bl[5] br[5] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_6 bl[6] br[6] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_7 bl[7] br[7] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_8 bl[8] br[8] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_9 bl[9] br[9] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_10 bl[10] br[10] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_11 bl[11] br[11] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_12 bl[12] br[12] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_13 bl[13] br[13] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_14 bl[14] br[14] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_15 bl[15] br[15] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_16 bl[16] br[16] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_17 bl[17] br[17] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_18 bl[18] br[18] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_19 bl[19] br[19] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_20 bl[20] br[20] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_21 bl[21] br[21] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_22 bl[22] br[22] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_23 bl[23] br[23] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_24 bl[24] br[24] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_25 bl[25] br[25] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_26 bl[26] br[26] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_27 bl[27] br[27] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_28 bl[28] br[28] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_29 bl[29] br[29] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_30 bl[30] br[30] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_31 bl[31] br[31] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_32 bl[32] br[32] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_33 bl[33] br[33] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_34 bl[34] br[34] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_35 bl[35] br[35] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_36 bl[36] br[36] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_37 bl[37] br[37] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_38 bl[38] br[38] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_39 bl[39] br[39] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_40 bl[40] br[40] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_41 bl[41] br[41] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_42 bl[42] br[42] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_43 bl[43] br[43] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_44 bl[44] br[44] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_45 bl[45] br[45] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_46 bl[46] br[46] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_47 bl[47] br[47] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_48 bl[48] br[48] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_49 bl[49] br[49] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_50 bl[50] br[50] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_51 bl[51] br[51] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_52 bl[52] br[52] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_53 bl[53] br[53] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_54 bl[54] br[54] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_55 bl[55] br[55] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_56 bl[56] br[56] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_57 bl[57] br[57] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_58 bl[58] br[58] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_59 bl[59] br[59] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_60 bl[60] br[60] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_61 bl[61] br[61] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_62 bl[62] br[62] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_63 bl[63] br[63] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_64 bl[64] br[64] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_65 bl[65] br[65] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_66 bl[66] br[66] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_67 bl[67] br[67] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_68 bl[68] br[68] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_69 bl[69] br[69] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_70 bl[70] br[70] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_71 bl[71] br[71] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_72 bl[72] br[72] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_73 bl[73] br[73] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_74 bl[74] br[74] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_75 bl[75] br[75] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_76 bl[76] br[76] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_77 bl[77] br[77] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_78 bl[78] br[78] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_79 bl[79] br[79] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_80 bl[80] br[80] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_81 bl[81] br[81] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_82 bl[82] br[82] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_83 bl[83] br[83] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_84 bl[84] br[84] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_85 bl[85] br[85] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_86 bl[86] br[86] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_87 bl[87] br[87] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_88 bl[88] br[88] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_89 bl[89] br[89] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_90 bl[90] br[90] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_91 bl[91] br[91] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_92 bl[92] br[92] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_93 bl[93] br[93] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_94 bl[94] br[94] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_95 bl[95] br[95] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_96 bl[96] br[96] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_97 bl[97] br[97] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_98 bl[98] br[98] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_99 bl[99] br[99] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_100 bl[100] br[100] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_101 bl[101] br[101] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_102 bl[102] br[102] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_103 bl[103] br[103] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_104 bl[104] br[104] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_105 bl[105] br[105] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_106 bl[106] br[106] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_107 bl[107] br[107] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_108 bl[108] br[108] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_109 bl[109] br[109] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_110 bl[110] br[110] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_111 bl[111] br[111] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_112 bl[112] br[112] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_113 bl[113] br[113] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_114 bl[114] br[114] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_115 bl[115] br[115] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_116 bl[116] br[116] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_117 bl[117] br[117] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_118 bl[118] br[118] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_119 bl[119] br[119] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_120 bl[120] br[120] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_121 bl[121] br[121] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_122 bl[122] br[122] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_123 bl[123] br[123] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_124 bl[124] br[124] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_125 bl[125] br[125] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_126 bl[126] br[126] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_127 bl[127] br[127] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_128 bl[128] br[128] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_129 bl[129] br[129] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_130 bl[130] br[130] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_131 bl[131] br[131] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_132 bl[132] br[132] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_133 bl[133] br[133] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_134 bl[134] br[134] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_135 bl[135] br[135] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_136 bl[136] br[136] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_137 bl[137] br[137] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_138 bl[138] br[138] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_139 bl[139] br[139] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_140 bl[140] br[140] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_141 bl[141] br[141] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_142 bl[142] br[142] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_143 bl[143] br[143] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_144 bl[144] br[144] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_145 bl[145] br[145] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_146 bl[146] br[146] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_147 bl[147] br[147] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_148 bl[148] br[148] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_149 bl[149] br[149] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_150 bl[150] br[150] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_151 bl[151] br[151] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_152 bl[152] br[152] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_153 bl[153] br[153] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_154 bl[154] br[154] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_155 bl[155] br[155] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_156 bl[156] br[156] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_157 bl[157] br[157] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_158 bl[158] br[158] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_159 bl[159] br[159] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_160 bl[160] br[160] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_161 bl[161] br[161] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_162 bl[162] br[162] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_163 bl[163] br[163] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_164 bl[164] br[164] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_165 bl[165] br[165] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_166 bl[166] br[166] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_167 bl[167] br[167] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_168 bl[168] br[168] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_169 bl[169] br[169] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_170 bl[170] br[170] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_171 bl[171] br[171] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_172 bl[172] br[172] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_173 bl[173] br[173] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_174 bl[174] br[174] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_175 bl[175] br[175] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_176 bl[176] br[176] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_177 bl[177] br[177] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_178 bl[178] br[178] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_179 bl[179] br[179] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_180 bl[180] br[180] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_181 bl[181] br[181] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_182 bl[182] br[182] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_183 bl[183] br[183] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_184 bl[184] br[184] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_185 bl[185] br[185] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_186 bl[186] br[186] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_187 bl[187] br[187] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_188 bl[188] br[188] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_189 bl[189] br[189] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_190 bl[190] br[190] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_191 bl[191] br[191] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_192 bl[192] br[192] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_193 bl[193] br[193] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_194 bl[194] br[194] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_195 bl[195] br[195] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_196 bl[196] br[196] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_197 bl[197] br[197] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_198 bl[198] br[198] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_199 bl[199] br[199] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_200 bl[200] br[200] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_201 bl[201] br[201] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_202 bl[202] br[202] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_203 bl[203] br[203] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_204 bl[204] br[204] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_205 bl[205] br[205] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_206 bl[206] br[206] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_207 bl[207] br[207] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_208 bl[208] br[208] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_209 bl[209] br[209] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_210 bl[210] br[210] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_211 bl[211] br[211] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_212 bl[212] br[212] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_213 bl[213] br[213] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_214 bl[214] br[214] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_215 bl[215] br[215] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_216 bl[216] br[216] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_217 bl[217] br[217] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_218 bl[218] br[218] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_219 bl[219] br[219] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_220 bl[220] br[220] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_221 bl[221] br[221] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_222 bl[222] br[222] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_223 bl[223] br[223] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_224 bl[224] br[224] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_225 bl[225] br[225] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_226 bl[226] br[226] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_227 bl[227] br[227] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_228 bl[228] br[228] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_229 bl[229] br[229] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_230 bl[230] br[230] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_231 bl[231] br[231] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_232 bl[232] br[232] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_233 bl[233] br[233] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_234 bl[234] br[234] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_235 bl[235] br[235] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_236 bl[236] br[236] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_237 bl[237] br[237] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_238 bl[238] br[238] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_239 bl[239] br[239] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_240 bl[240] br[240] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_241 bl[241] br[241] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_242 bl[242] br[242] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_243 bl[243] br[243] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_244 bl[244] br[244] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_245 bl[245] br[245] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_246 bl[246] br[246] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_247 bl[247] br[247] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_248 bl[248] br[248] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_249 bl[249] br[249] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_250 bl[250] br[250] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_251 bl[251] br[251] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_252 bl[252] br[252] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_253 bl[253] br[253] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_254 bl[254] br[254] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_255 bl[255] br[255] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_71_0 bl[0] br[0] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_1 bl[1] br[1] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_2 bl[2] br[2] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_3 bl[3] br[3] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_4 bl[4] br[4] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_5 bl[5] br[5] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_6 bl[6] br[6] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_7 bl[7] br[7] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_8 bl[8] br[8] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_9 bl[9] br[9] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_10 bl[10] br[10] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_11 bl[11] br[11] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_12 bl[12] br[12] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_13 bl[13] br[13] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_14 bl[14] br[14] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_15 bl[15] br[15] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_16 bl[16] br[16] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_17 bl[17] br[17] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_18 bl[18] br[18] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_19 bl[19] br[19] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_20 bl[20] br[20] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_21 bl[21] br[21] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_22 bl[22] br[22] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_23 bl[23] br[23] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_24 bl[24] br[24] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_25 bl[25] br[25] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_26 bl[26] br[26] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_27 bl[27] br[27] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_28 bl[28] br[28] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_29 bl[29] br[29] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_30 bl[30] br[30] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_31 bl[31] br[31] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_32 bl[32] br[32] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_33 bl[33] br[33] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_34 bl[34] br[34] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_35 bl[35] br[35] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_36 bl[36] br[36] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_37 bl[37] br[37] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_38 bl[38] br[38] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_39 bl[39] br[39] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_40 bl[40] br[40] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_41 bl[41] br[41] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_42 bl[42] br[42] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_43 bl[43] br[43] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_44 bl[44] br[44] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_45 bl[45] br[45] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_46 bl[46] br[46] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_47 bl[47] br[47] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_48 bl[48] br[48] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_49 bl[49] br[49] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_50 bl[50] br[50] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_51 bl[51] br[51] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_52 bl[52] br[52] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_53 bl[53] br[53] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_54 bl[54] br[54] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_55 bl[55] br[55] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_56 bl[56] br[56] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_57 bl[57] br[57] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_58 bl[58] br[58] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_59 bl[59] br[59] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_60 bl[60] br[60] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_61 bl[61] br[61] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_62 bl[62] br[62] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_63 bl[63] br[63] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_64 bl[64] br[64] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_65 bl[65] br[65] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_66 bl[66] br[66] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_67 bl[67] br[67] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_68 bl[68] br[68] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_69 bl[69] br[69] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_70 bl[70] br[70] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_71 bl[71] br[71] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_72 bl[72] br[72] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_73 bl[73] br[73] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_74 bl[74] br[74] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_75 bl[75] br[75] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_76 bl[76] br[76] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_77 bl[77] br[77] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_78 bl[78] br[78] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_79 bl[79] br[79] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_80 bl[80] br[80] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_81 bl[81] br[81] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_82 bl[82] br[82] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_83 bl[83] br[83] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_84 bl[84] br[84] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_85 bl[85] br[85] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_86 bl[86] br[86] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_87 bl[87] br[87] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_88 bl[88] br[88] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_89 bl[89] br[89] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_90 bl[90] br[90] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_91 bl[91] br[91] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_92 bl[92] br[92] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_93 bl[93] br[93] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_94 bl[94] br[94] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_95 bl[95] br[95] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_96 bl[96] br[96] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_97 bl[97] br[97] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_98 bl[98] br[98] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_99 bl[99] br[99] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_100 bl[100] br[100] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_101 bl[101] br[101] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_102 bl[102] br[102] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_103 bl[103] br[103] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_104 bl[104] br[104] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_105 bl[105] br[105] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_106 bl[106] br[106] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_107 bl[107] br[107] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_108 bl[108] br[108] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_109 bl[109] br[109] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_110 bl[110] br[110] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_111 bl[111] br[111] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_112 bl[112] br[112] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_113 bl[113] br[113] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_114 bl[114] br[114] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_115 bl[115] br[115] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_116 bl[116] br[116] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_117 bl[117] br[117] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_118 bl[118] br[118] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_119 bl[119] br[119] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_120 bl[120] br[120] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_121 bl[121] br[121] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_122 bl[122] br[122] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_123 bl[123] br[123] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_124 bl[124] br[124] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_125 bl[125] br[125] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_126 bl[126] br[126] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_127 bl[127] br[127] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_128 bl[128] br[128] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_129 bl[129] br[129] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_130 bl[130] br[130] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_131 bl[131] br[131] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_132 bl[132] br[132] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_133 bl[133] br[133] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_134 bl[134] br[134] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_135 bl[135] br[135] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_136 bl[136] br[136] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_137 bl[137] br[137] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_138 bl[138] br[138] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_139 bl[139] br[139] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_140 bl[140] br[140] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_141 bl[141] br[141] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_142 bl[142] br[142] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_143 bl[143] br[143] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_144 bl[144] br[144] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_145 bl[145] br[145] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_146 bl[146] br[146] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_147 bl[147] br[147] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_148 bl[148] br[148] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_149 bl[149] br[149] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_150 bl[150] br[150] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_151 bl[151] br[151] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_152 bl[152] br[152] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_153 bl[153] br[153] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_154 bl[154] br[154] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_155 bl[155] br[155] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_156 bl[156] br[156] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_157 bl[157] br[157] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_158 bl[158] br[158] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_159 bl[159] br[159] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_160 bl[160] br[160] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_161 bl[161] br[161] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_162 bl[162] br[162] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_163 bl[163] br[163] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_164 bl[164] br[164] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_165 bl[165] br[165] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_166 bl[166] br[166] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_167 bl[167] br[167] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_168 bl[168] br[168] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_169 bl[169] br[169] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_170 bl[170] br[170] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_171 bl[171] br[171] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_172 bl[172] br[172] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_173 bl[173] br[173] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_174 bl[174] br[174] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_175 bl[175] br[175] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_176 bl[176] br[176] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_177 bl[177] br[177] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_178 bl[178] br[178] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_179 bl[179] br[179] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_180 bl[180] br[180] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_181 bl[181] br[181] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_182 bl[182] br[182] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_183 bl[183] br[183] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_184 bl[184] br[184] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_185 bl[185] br[185] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_186 bl[186] br[186] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_187 bl[187] br[187] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_188 bl[188] br[188] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_189 bl[189] br[189] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_190 bl[190] br[190] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_191 bl[191] br[191] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_192 bl[192] br[192] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_193 bl[193] br[193] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_194 bl[194] br[194] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_195 bl[195] br[195] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_196 bl[196] br[196] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_197 bl[197] br[197] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_198 bl[198] br[198] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_199 bl[199] br[199] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_200 bl[200] br[200] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_201 bl[201] br[201] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_202 bl[202] br[202] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_203 bl[203] br[203] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_204 bl[204] br[204] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_205 bl[205] br[205] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_206 bl[206] br[206] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_207 bl[207] br[207] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_208 bl[208] br[208] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_209 bl[209] br[209] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_210 bl[210] br[210] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_211 bl[211] br[211] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_212 bl[212] br[212] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_213 bl[213] br[213] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_214 bl[214] br[214] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_215 bl[215] br[215] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_216 bl[216] br[216] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_217 bl[217] br[217] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_218 bl[218] br[218] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_219 bl[219] br[219] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_220 bl[220] br[220] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_221 bl[221] br[221] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_222 bl[222] br[222] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_223 bl[223] br[223] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_224 bl[224] br[224] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_225 bl[225] br[225] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_226 bl[226] br[226] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_227 bl[227] br[227] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_228 bl[228] br[228] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_229 bl[229] br[229] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_230 bl[230] br[230] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_231 bl[231] br[231] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_232 bl[232] br[232] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_233 bl[233] br[233] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_234 bl[234] br[234] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_235 bl[235] br[235] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_236 bl[236] br[236] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_237 bl[237] br[237] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_238 bl[238] br[238] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_239 bl[239] br[239] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_240 bl[240] br[240] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_241 bl[241] br[241] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_242 bl[242] br[242] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_243 bl[243] br[243] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_244 bl[244] br[244] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_245 bl[245] br[245] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_246 bl[246] br[246] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_247 bl[247] br[247] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_248 bl[248] br[248] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_249 bl[249] br[249] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_250 bl[250] br[250] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_251 bl[251] br[251] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_252 bl[252] br[252] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_253 bl[253] br[253] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_254 bl[254] br[254] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_255 bl[255] br[255] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_72_0 bl[0] br[0] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_1 bl[1] br[1] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_2 bl[2] br[2] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_3 bl[3] br[3] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_4 bl[4] br[4] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_5 bl[5] br[5] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_6 bl[6] br[6] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_7 bl[7] br[7] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_8 bl[8] br[8] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_9 bl[9] br[9] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_10 bl[10] br[10] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_11 bl[11] br[11] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_12 bl[12] br[12] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_13 bl[13] br[13] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_14 bl[14] br[14] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_15 bl[15] br[15] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_16 bl[16] br[16] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_17 bl[17] br[17] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_18 bl[18] br[18] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_19 bl[19] br[19] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_20 bl[20] br[20] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_21 bl[21] br[21] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_22 bl[22] br[22] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_23 bl[23] br[23] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_24 bl[24] br[24] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_25 bl[25] br[25] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_26 bl[26] br[26] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_27 bl[27] br[27] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_28 bl[28] br[28] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_29 bl[29] br[29] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_30 bl[30] br[30] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_31 bl[31] br[31] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_32 bl[32] br[32] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_33 bl[33] br[33] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_34 bl[34] br[34] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_35 bl[35] br[35] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_36 bl[36] br[36] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_37 bl[37] br[37] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_38 bl[38] br[38] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_39 bl[39] br[39] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_40 bl[40] br[40] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_41 bl[41] br[41] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_42 bl[42] br[42] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_43 bl[43] br[43] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_44 bl[44] br[44] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_45 bl[45] br[45] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_46 bl[46] br[46] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_47 bl[47] br[47] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_48 bl[48] br[48] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_49 bl[49] br[49] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_50 bl[50] br[50] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_51 bl[51] br[51] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_52 bl[52] br[52] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_53 bl[53] br[53] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_54 bl[54] br[54] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_55 bl[55] br[55] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_56 bl[56] br[56] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_57 bl[57] br[57] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_58 bl[58] br[58] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_59 bl[59] br[59] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_60 bl[60] br[60] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_61 bl[61] br[61] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_62 bl[62] br[62] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_63 bl[63] br[63] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_64 bl[64] br[64] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_65 bl[65] br[65] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_66 bl[66] br[66] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_67 bl[67] br[67] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_68 bl[68] br[68] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_69 bl[69] br[69] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_70 bl[70] br[70] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_71 bl[71] br[71] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_72 bl[72] br[72] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_73 bl[73] br[73] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_74 bl[74] br[74] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_75 bl[75] br[75] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_76 bl[76] br[76] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_77 bl[77] br[77] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_78 bl[78] br[78] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_79 bl[79] br[79] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_80 bl[80] br[80] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_81 bl[81] br[81] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_82 bl[82] br[82] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_83 bl[83] br[83] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_84 bl[84] br[84] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_85 bl[85] br[85] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_86 bl[86] br[86] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_87 bl[87] br[87] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_88 bl[88] br[88] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_89 bl[89] br[89] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_90 bl[90] br[90] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_91 bl[91] br[91] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_92 bl[92] br[92] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_93 bl[93] br[93] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_94 bl[94] br[94] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_95 bl[95] br[95] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_96 bl[96] br[96] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_97 bl[97] br[97] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_98 bl[98] br[98] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_99 bl[99] br[99] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_100 bl[100] br[100] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_101 bl[101] br[101] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_102 bl[102] br[102] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_103 bl[103] br[103] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_104 bl[104] br[104] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_105 bl[105] br[105] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_106 bl[106] br[106] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_107 bl[107] br[107] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_108 bl[108] br[108] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_109 bl[109] br[109] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_110 bl[110] br[110] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_111 bl[111] br[111] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_112 bl[112] br[112] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_113 bl[113] br[113] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_114 bl[114] br[114] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_115 bl[115] br[115] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_116 bl[116] br[116] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_117 bl[117] br[117] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_118 bl[118] br[118] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_119 bl[119] br[119] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_120 bl[120] br[120] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_121 bl[121] br[121] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_122 bl[122] br[122] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_123 bl[123] br[123] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_124 bl[124] br[124] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_125 bl[125] br[125] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_126 bl[126] br[126] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_127 bl[127] br[127] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_128 bl[128] br[128] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_129 bl[129] br[129] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_130 bl[130] br[130] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_131 bl[131] br[131] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_132 bl[132] br[132] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_133 bl[133] br[133] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_134 bl[134] br[134] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_135 bl[135] br[135] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_136 bl[136] br[136] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_137 bl[137] br[137] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_138 bl[138] br[138] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_139 bl[139] br[139] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_140 bl[140] br[140] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_141 bl[141] br[141] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_142 bl[142] br[142] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_143 bl[143] br[143] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_144 bl[144] br[144] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_145 bl[145] br[145] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_146 bl[146] br[146] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_147 bl[147] br[147] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_148 bl[148] br[148] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_149 bl[149] br[149] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_150 bl[150] br[150] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_151 bl[151] br[151] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_152 bl[152] br[152] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_153 bl[153] br[153] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_154 bl[154] br[154] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_155 bl[155] br[155] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_156 bl[156] br[156] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_157 bl[157] br[157] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_158 bl[158] br[158] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_159 bl[159] br[159] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_160 bl[160] br[160] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_161 bl[161] br[161] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_162 bl[162] br[162] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_163 bl[163] br[163] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_164 bl[164] br[164] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_165 bl[165] br[165] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_166 bl[166] br[166] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_167 bl[167] br[167] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_168 bl[168] br[168] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_169 bl[169] br[169] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_170 bl[170] br[170] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_171 bl[171] br[171] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_172 bl[172] br[172] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_173 bl[173] br[173] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_174 bl[174] br[174] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_175 bl[175] br[175] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_176 bl[176] br[176] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_177 bl[177] br[177] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_178 bl[178] br[178] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_179 bl[179] br[179] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_180 bl[180] br[180] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_181 bl[181] br[181] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_182 bl[182] br[182] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_183 bl[183] br[183] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_184 bl[184] br[184] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_185 bl[185] br[185] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_186 bl[186] br[186] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_187 bl[187] br[187] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_188 bl[188] br[188] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_189 bl[189] br[189] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_190 bl[190] br[190] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_191 bl[191] br[191] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_192 bl[192] br[192] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_193 bl[193] br[193] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_194 bl[194] br[194] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_195 bl[195] br[195] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_196 bl[196] br[196] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_197 bl[197] br[197] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_198 bl[198] br[198] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_199 bl[199] br[199] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_200 bl[200] br[200] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_201 bl[201] br[201] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_202 bl[202] br[202] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_203 bl[203] br[203] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_204 bl[204] br[204] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_205 bl[205] br[205] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_206 bl[206] br[206] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_207 bl[207] br[207] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_208 bl[208] br[208] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_209 bl[209] br[209] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_210 bl[210] br[210] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_211 bl[211] br[211] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_212 bl[212] br[212] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_213 bl[213] br[213] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_214 bl[214] br[214] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_215 bl[215] br[215] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_216 bl[216] br[216] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_217 bl[217] br[217] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_218 bl[218] br[218] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_219 bl[219] br[219] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_220 bl[220] br[220] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_221 bl[221] br[221] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_222 bl[222] br[222] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_223 bl[223] br[223] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_224 bl[224] br[224] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_225 bl[225] br[225] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_226 bl[226] br[226] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_227 bl[227] br[227] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_228 bl[228] br[228] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_229 bl[229] br[229] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_230 bl[230] br[230] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_231 bl[231] br[231] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_232 bl[232] br[232] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_233 bl[233] br[233] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_234 bl[234] br[234] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_235 bl[235] br[235] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_236 bl[236] br[236] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_237 bl[237] br[237] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_238 bl[238] br[238] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_239 bl[239] br[239] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_240 bl[240] br[240] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_241 bl[241] br[241] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_242 bl[242] br[242] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_243 bl[243] br[243] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_244 bl[244] br[244] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_245 bl[245] br[245] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_246 bl[246] br[246] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_247 bl[247] br[247] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_248 bl[248] br[248] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_249 bl[249] br[249] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_250 bl[250] br[250] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_251 bl[251] br[251] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_252 bl[252] br[252] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_253 bl[253] br[253] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_254 bl[254] br[254] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_255 bl[255] br[255] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_73_0 bl[0] br[0] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_1 bl[1] br[1] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_2 bl[2] br[2] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_3 bl[3] br[3] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_4 bl[4] br[4] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_5 bl[5] br[5] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_6 bl[6] br[6] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_7 bl[7] br[7] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_8 bl[8] br[8] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_9 bl[9] br[9] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_10 bl[10] br[10] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_11 bl[11] br[11] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_12 bl[12] br[12] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_13 bl[13] br[13] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_14 bl[14] br[14] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_15 bl[15] br[15] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_16 bl[16] br[16] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_17 bl[17] br[17] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_18 bl[18] br[18] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_19 bl[19] br[19] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_20 bl[20] br[20] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_21 bl[21] br[21] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_22 bl[22] br[22] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_23 bl[23] br[23] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_24 bl[24] br[24] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_25 bl[25] br[25] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_26 bl[26] br[26] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_27 bl[27] br[27] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_28 bl[28] br[28] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_29 bl[29] br[29] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_30 bl[30] br[30] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_31 bl[31] br[31] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_32 bl[32] br[32] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_33 bl[33] br[33] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_34 bl[34] br[34] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_35 bl[35] br[35] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_36 bl[36] br[36] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_37 bl[37] br[37] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_38 bl[38] br[38] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_39 bl[39] br[39] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_40 bl[40] br[40] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_41 bl[41] br[41] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_42 bl[42] br[42] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_43 bl[43] br[43] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_44 bl[44] br[44] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_45 bl[45] br[45] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_46 bl[46] br[46] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_47 bl[47] br[47] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_48 bl[48] br[48] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_49 bl[49] br[49] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_50 bl[50] br[50] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_51 bl[51] br[51] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_52 bl[52] br[52] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_53 bl[53] br[53] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_54 bl[54] br[54] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_55 bl[55] br[55] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_56 bl[56] br[56] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_57 bl[57] br[57] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_58 bl[58] br[58] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_59 bl[59] br[59] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_60 bl[60] br[60] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_61 bl[61] br[61] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_62 bl[62] br[62] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_63 bl[63] br[63] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_64 bl[64] br[64] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_65 bl[65] br[65] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_66 bl[66] br[66] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_67 bl[67] br[67] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_68 bl[68] br[68] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_69 bl[69] br[69] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_70 bl[70] br[70] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_71 bl[71] br[71] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_72 bl[72] br[72] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_73 bl[73] br[73] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_74 bl[74] br[74] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_75 bl[75] br[75] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_76 bl[76] br[76] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_77 bl[77] br[77] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_78 bl[78] br[78] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_79 bl[79] br[79] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_80 bl[80] br[80] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_81 bl[81] br[81] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_82 bl[82] br[82] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_83 bl[83] br[83] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_84 bl[84] br[84] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_85 bl[85] br[85] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_86 bl[86] br[86] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_87 bl[87] br[87] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_88 bl[88] br[88] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_89 bl[89] br[89] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_90 bl[90] br[90] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_91 bl[91] br[91] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_92 bl[92] br[92] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_93 bl[93] br[93] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_94 bl[94] br[94] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_95 bl[95] br[95] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_96 bl[96] br[96] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_97 bl[97] br[97] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_98 bl[98] br[98] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_99 bl[99] br[99] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_100 bl[100] br[100] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_101 bl[101] br[101] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_102 bl[102] br[102] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_103 bl[103] br[103] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_104 bl[104] br[104] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_105 bl[105] br[105] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_106 bl[106] br[106] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_107 bl[107] br[107] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_108 bl[108] br[108] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_109 bl[109] br[109] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_110 bl[110] br[110] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_111 bl[111] br[111] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_112 bl[112] br[112] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_113 bl[113] br[113] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_114 bl[114] br[114] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_115 bl[115] br[115] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_116 bl[116] br[116] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_117 bl[117] br[117] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_118 bl[118] br[118] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_119 bl[119] br[119] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_120 bl[120] br[120] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_121 bl[121] br[121] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_122 bl[122] br[122] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_123 bl[123] br[123] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_124 bl[124] br[124] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_125 bl[125] br[125] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_126 bl[126] br[126] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_127 bl[127] br[127] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_128 bl[128] br[128] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_129 bl[129] br[129] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_130 bl[130] br[130] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_131 bl[131] br[131] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_132 bl[132] br[132] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_133 bl[133] br[133] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_134 bl[134] br[134] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_135 bl[135] br[135] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_136 bl[136] br[136] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_137 bl[137] br[137] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_138 bl[138] br[138] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_139 bl[139] br[139] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_140 bl[140] br[140] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_141 bl[141] br[141] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_142 bl[142] br[142] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_143 bl[143] br[143] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_144 bl[144] br[144] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_145 bl[145] br[145] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_146 bl[146] br[146] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_147 bl[147] br[147] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_148 bl[148] br[148] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_149 bl[149] br[149] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_150 bl[150] br[150] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_151 bl[151] br[151] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_152 bl[152] br[152] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_153 bl[153] br[153] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_154 bl[154] br[154] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_155 bl[155] br[155] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_156 bl[156] br[156] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_157 bl[157] br[157] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_158 bl[158] br[158] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_159 bl[159] br[159] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_160 bl[160] br[160] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_161 bl[161] br[161] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_162 bl[162] br[162] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_163 bl[163] br[163] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_164 bl[164] br[164] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_165 bl[165] br[165] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_166 bl[166] br[166] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_167 bl[167] br[167] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_168 bl[168] br[168] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_169 bl[169] br[169] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_170 bl[170] br[170] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_171 bl[171] br[171] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_172 bl[172] br[172] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_173 bl[173] br[173] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_174 bl[174] br[174] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_175 bl[175] br[175] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_176 bl[176] br[176] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_177 bl[177] br[177] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_178 bl[178] br[178] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_179 bl[179] br[179] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_180 bl[180] br[180] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_181 bl[181] br[181] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_182 bl[182] br[182] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_183 bl[183] br[183] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_184 bl[184] br[184] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_185 bl[185] br[185] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_186 bl[186] br[186] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_187 bl[187] br[187] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_188 bl[188] br[188] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_189 bl[189] br[189] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_190 bl[190] br[190] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_191 bl[191] br[191] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_192 bl[192] br[192] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_193 bl[193] br[193] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_194 bl[194] br[194] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_195 bl[195] br[195] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_196 bl[196] br[196] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_197 bl[197] br[197] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_198 bl[198] br[198] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_199 bl[199] br[199] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_200 bl[200] br[200] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_201 bl[201] br[201] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_202 bl[202] br[202] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_203 bl[203] br[203] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_204 bl[204] br[204] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_205 bl[205] br[205] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_206 bl[206] br[206] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_207 bl[207] br[207] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_208 bl[208] br[208] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_209 bl[209] br[209] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_210 bl[210] br[210] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_211 bl[211] br[211] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_212 bl[212] br[212] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_213 bl[213] br[213] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_214 bl[214] br[214] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_215 bl[215] br[215] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_216 bl[216] br[216] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_217 bl[217] br[217] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_218 bl[218] br[218] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_219 bl[219] br[219] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_220 bl[220] br[220] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_221 bl[221] br[221] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_222 bl[222] br[222] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_223 bl[223] br[223] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_224 bl[224] br[224] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_225 bl[225] br[225] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_226 bl[226] br[226] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_227 bl[227] br[227] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_228 bl[228] br[228] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_229 bl[229] br[229] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_230 bl[230] br[230] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_231 bl[231] br[231] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_232 bl[232] br[232] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_233 bl[233] br[233] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_234 bl[234] br[234] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_235 bl[235] br[235] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_236 bl[236] br[236] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_237 bl[237] br[237] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_238 bl[238] br[238] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_239 bl[239] br[239] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_240 bl[240] br[240] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_241 bl[241] br[241] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_242 bl[242] br[242] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_243 bl[243] br[243] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_244 bl[244] br[244] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_245 bl[245] br[245] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_246 bl[246] br[246] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_247 bl[247] br[247] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_248 bl[248] br[248] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_249 bl[249] br[249] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_250 bl[250] br[250] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_251 bl[251] br[251] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_252 bl[252] br[252] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_253 bl[253] br[253] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_254 bl[254] br[254] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_255 bl[255] br[255] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_74_0 bl[0] br[0] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_1 bl[1] br[1] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_2 bl[2] br[2] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_3 bl[3] br[3] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_4 bl[4] br[4] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_5 bl[5] br[5] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_6 bl[6] br[6] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_7 bl[7] br[7] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_8 bl[8] br[8] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_9 bl[9] br[9] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_10 bl[10] br[10] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_11 bl[11] br[11] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_12 bl[12] br[12] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_13 bl[13] br[13] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_14 bl[14] br[14] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_15 bl[15] br[15] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_16 bl[16] br[16] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_17 bl[17] br[17] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_18 bl[18] br[18] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_19 bl[19] br[19] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_20 bl[20] br[20] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_21 bl[21] br[21] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_22 bl[22] br[22] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_23 bl[23] br[23] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_24 bl[24] br[24] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_25 bl[25] br[25] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_26 bl[26] br[26] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_27 bl[27] br[27] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_28 bl[28] br[28] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_29 bl[29] br[29] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_30 bl[30] br[30] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_31 bl[31] br[31] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_32 bl[32] br[32] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_33 bl[33] br[33] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_34 bl[34] br[34] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_35 bl[35] br[35] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_36 bl[36] br[36] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_37 bl[37] br[37] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_38 bl[38] br[38] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_39 bl[39] br[39] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_40 bl[40] br[40] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_41 bl[41] br[41] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_42 bl[42] br[42] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_43 bl[43] br[43] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_44 bl[44] br[44] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_45 bl[45] br[45] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_46 bl[46] br[46] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_47 bl[47] br[47] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_48 bl[48] br[48] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_49 bl[49] br[49] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_50 bl[50] br[50] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_51 bl[51] br[51] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_52 bl[52] br[52] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_53 bl[53] br[53] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_54 bl[54] br[54] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_55 bl[55] br[55] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_56 bl[56] br[56] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_57 bl[57] br[57] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_58 bl[58] br[58] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_59 bl[59] br[59] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_60 bl[60] br[60] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_61 bl[61] br[61] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_62 bl[62] br[62] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_63 bl[63] br[63] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_64 bl[64] br[64] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_65 bl[65] br[65] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_66 bl[66] br[66] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_67 bl[67] br[67] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_68 bl[68] br[68] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_69 bl[69] br[69] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_70 bl[70] br[70] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_71 bl[71] br[71] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_72 bl[72] br[72] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_73 bl[73] br[73] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_74 bl[74] br[74] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_75 bl[75] br[75] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_76 bl[76] br[76] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_77 bl[77] br[77] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_78 bl[78] br[78] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_79 bl[79] br[79] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_80 bl[80] br[80] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_81 bl[81] br[81] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_82 bl[82] br[82] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_83 bl[83] br[83] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_84 bl[84] br[84] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_85 bl[85] br[85] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_86 bl[86] br[86] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_87 bl[87] br[87] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_88 bl[88] br[88] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_89 bl[89] br[89] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_90 bl[90] br[90] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_91 bl[91] br[91] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_92 bl[92] br[92] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_93 bl[93] br[93] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_94 bl[94] br[94] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_95 bl[95] br[95] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_96 bl[96] br[96] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_97 bl[97] br[97] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_98 bl[98] br[98] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_99 bl[99] br[99] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_100 bl[100] br[100] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_101 bl[101] br[101] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_102 bl[102] br[102] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_103 bl[103] br[103] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_104 bl[104] br[104] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_105 bl[105] br[105] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_106 bl[106] br[106] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_107 bl[107] br[107] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_108 bl[108] br[108] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_109 bl[109] br[109] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_110 bl[110] br[110] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_111 bl[111] br[111] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_112 bl[112] br[112] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_113 bl[113] br[113] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_114 bl[114] br[114] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_115 bl[115] br[115] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_116 bl[116] br[116] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_117 bl[117] br[117] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_118 bl[118] br[118] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_119 bl[119] br[119] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_120 bl[120] br[120] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_121 bl[121] br[121] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_122 bl[122] br[122] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_123 bl[123] br[123] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_124 bl[124] br[124] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_125 bl[125] br[125] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_126 bl[126] br[126] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_127 bl[127] br[127] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_128 bl[128] br[128] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_129 bl[129] br[129] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_130 bl[130] br[130] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_131 bl[131] br[131] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_132 bl[132] br[132] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_133 bl[133] br[133] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_134 bl[134] br[134] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_135 bl[135] br[135] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_136 bl[136] br[136] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_137 bl[137] br[137] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_138 bl[138] br[138] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_139 bl[139] br[139] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_140 bl[140] br[140] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_141 bl[141] br[141] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_142 bl[142] br[142] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_143 bl[143] br[143] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_144 bl[144] br[144] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_145 bl[145] br[145] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_146 bl[146] br[146] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_147 bl[147] br[147] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_148 bl[148] br[148] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_149 bl[149] br[149] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_150 bl[150] br[150] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_151 bl[151] br[151] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_152 bl[152] br[152] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_153 bl[153] br[153] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_154 bl[154] br[154] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_155 bl[155] br[155] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_156 bl[156] br[156] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_157 bl[157] br[157] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_158 bl[158] br[158] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_159 bl[159] br[159] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_160 bl[160] br[160] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_161 bl[161] br[161] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_162 bl[162] br[162] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_163 bl[163] br[163] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_164 bl[164] br[164] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_165 bl[165] br[165] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_166 bl[166] br[166] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_167 bl[167] br[167] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_168 bl[168] br[168] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_169 bl[169] br[169] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_170 bl[170] br[170] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_171 bl[171] br[171] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_172 bl[172] br[172] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_173 bl[173] br[173] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_174 bl[174] br[174] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_175 bl[175] br[175] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_176 bl[176] br[176] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_177 bl[177] br[177] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_178 bl[178] br[178] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_179 bl[179] br[179] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_180 bl[180] br[180] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_181 bl[181] br[181] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_182 bl[182] br[182] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_183 bl[183] br[183] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_184 bl[184] br[184] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_185 bl[185] br[185] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_186 bl[186] br[186] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_187 bl[187] br[187] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_188 bl[188] br[188] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_189 bl[189] br[189] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_190 bl[190] br[190] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_191 bl[191] br[191] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_192 bl[192] br[192] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_193 bl[193] br[193] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_194 bl[194] br[194] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_195 bl[195] br[195] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_196 bl[196] br[196] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_197 bl[197] br[197] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_198 bl[198] br[198] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_199 bl[199] br[199] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_200 bl[200] br[200] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_201 bl[201] br[201] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_202 bl[202] br[202] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_203 bl[203] br[203] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_204 bl[204] br[204] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_205 bl[205] br[205] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_206 bl[206] br[206] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_207 bl[207] br[207] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_208 bl[208] br[208] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_209 bl[209] br[209] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_210 bl[210] br[210] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_211 bl[211] br[211] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_212 bl[212] br[212] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_213 bl[213] br[213] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_214 bl[214] br[214] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_215 bl[215] br[215] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_216 bl[216] br[216] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_217 bl[217] br[217] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_218 bl[218] br[218] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_219 bl[219] br[219] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_220 bl[220] br[220] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_221 bl[221] br[221] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_222 bl[222] br[222] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_223 bl[223] br[223] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_224 bl[224] br[224] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_225 bl[225] br[225] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_226 bl[226] br[226] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_227 bl[227] br[227] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_228 bl[228] br[228] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_229 bl[229] br[229] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_230 bl[230] br[230] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_231 bl[231] br[231] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_232 bl[232] br[232] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_233 bl[233] br[233] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_234 bl[234] br[234] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_235 bl[235] br[235] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_236 bl[236] br[236] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_237 bl[237] br[237] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_238 bl[238] br[238] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_239 bl[239] br[239] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_240 bl[240] br[240] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_241 bl[241] br[241] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_242 bl[242] br[242] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_243 bl[243] br[243] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_244 bl[244] br[244] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_245 bl[245] br[245] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_246 bl[246] br[246] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_247 bl[247] br[247] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_248 bl[248] br[248] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_249 bl[249] br[249] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_250 bl[250] br[250] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_251 bl[251] br[251] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_252 bl[252] br[252] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_253 bl[253] br[253] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_254 bl[254] br[254] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_255 bl[255] br[255] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_75_0 bl[0] br[0] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_1 bl[1] br[1] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_2 bl[2] br[2] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_3 bl[3] br[3] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_4 bl[4] br[4] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_5 bl[5] br[5] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_6 bl[6] br[6] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_7 bl[7] br[7] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_8 bl[8] br[8] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_9 bl[9] br[9] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_10 bl[10] br[10] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_11 bl[11] br[11] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_12 bl[12] br[12] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_13 bl[13] br[13] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_14 bl[14] br[14] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_15 bl[15] br[15] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_16 bl[16] br[16] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_17 bl[17] br[17] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_18 bl[18] br[18] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_19 bl[19] br[19] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_20 bl[20] br[20] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_21 bl[21] br[21] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_22 bl[22] br[22] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_23 bl[23] br[23] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_24 bl[24] br[24] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_25 bl[25] br[25] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_26 bl[26] br[26] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_27 bl[27] br[27] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_28 bl[28] br[28] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_29 bl[29] br[29] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_30 bl[30] br[30] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_31 bl[31] br[31] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_32 bl[32] br[32] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_33 bl[33] br[33] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_34 bl[34] br[34] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_35 bl[35] br[35] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_36 bl[36] br[36] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_37 bl[37] br[37] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_38 bl[38] br[38] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_39 bl[39] br[39] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_40 bl[40] br[40] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_41 bl[41] br[41] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_42 bl[42] br[42] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_43 bl[43] br[43] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_44 bl[44] br[44] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_45 bl[45] br[45] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_46 bl[46] br[46] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_47 bl[47] br[47] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_48 bl[48] br[48] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_49 bl[49] br[49] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_50 bl[50] br[50] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_51 bl[51] br[51] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_52 bl[52] br[52] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_53 bl[53] br[53] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_54 bl[54] br[54] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_55 bl[55] br[55] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_56 bl[56] br[56] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_57 bl[57] br[57] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_58 bl[58] br[58] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_59 bl[59] br[59] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_60 bl[60] br[60] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_61 bl[61] br[61] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_62 bl[62] br[62] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_63 bl[63] br[63] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_64 bl[64] br[64] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_65 bl[65] br[65] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_66 bl[66] br[66] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_67 bl[67] br[67] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_68 bl[68] br[68] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_69 bl[69] br[69] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_70 bl[70] br[70] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_71 bl[71] br[71] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_72 bl[72] br[72] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_73 bl[73] br[73] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_74 bl[74] br[74] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_75 bl[75] br[75] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_76 bl[76] br[76] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_77 bl[77] br[77] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_78 bl[78] br[78] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_79 bl[79] br[79] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_80 bl[80] br[80] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_81 bl[81] br[81] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_82 bl[82] br[82] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_83 bl[83] br[83] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_84 bl[84] br[84] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_85 bl[85] br[85] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_86 bl[86] br[86] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_87 bl[87] br[87] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_88 bl[88] br[88] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_89 bl[89] br[89] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_90 bl[90] br[90] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_91 bl[91] br[91] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_92 bl[92] br[92] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_93 bl[93] br[93] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_94 bl[94] br[94] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_95 bl[95] br[95] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_96 bl[96] br[96] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_97 bl[97] br[97] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_98 bl[98] br[98] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_99 bl[99] br[99] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_100 bl[100] br[100] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_101 bl[101] br[101] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_102 bl[102] br[102] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_103 bl[103] br[103] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_104 bl[104] br[104] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_105 bl[105] br[105] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_106 bl[106] br[106] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_107 bl[107] br[107] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_108 bl[108] br[108] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_109 bl[109] br[109] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_110 bl[110] br[110] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_111 bl[111] br[111] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_112 bl[112] br[112] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_113 bl[113] br[113] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_114 bl[114] br[114] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_115 bl[115] br[115] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_116 bl[116] br[116] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_117 bl[117] br[117] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_118 bl[118] br[118] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_119 bl[119] br[119] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_120 bl[120] br[120] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_121 bl[121] br[121] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_122 bl[122] br[122] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_123 bl[123] br[123] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_124 bl[124] br[124] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_125 bl[125] br[125] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_126 bl[126] br[126] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_127 bl[127] br[127] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_128 bl[128] br[128] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_129 bl[129] br[129] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_130 bl[130] br[130] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_131 bl[131] br[131] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_132 bl[132] br[132] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_133 bl[133] br[133] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_134 bl[134] br[134] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_135 bl[135] br[135] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_136 bl[136] br[136] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_137 bl[137] br[137] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_138 bl[138] br[138] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_139 bl[139] br[139] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_140 bl[140] br[140] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_141 bl[141] br[141] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_142 bl[142] br[142] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_143 bl[143] br[143] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_144 bl[144] br[144] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_145 bl[145] br[145] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_146 bl[146] br[146] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_147 bl[147] br[147] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_148 bl[148] br[148] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_149 bl[149] br[149] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_150 bl[150] br[150] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_151 bl[151] br[151] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_152 bl[152] br[152] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_153 bl[153] br[153] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_154 bl[154] br[154] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_155 bl[155] br[155] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_156 bl[156] br[156] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_157 bl[157] br[157] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_158 bl[158] br[158] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_159 bl[159] br[159] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_160 bl[160] br[160] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_161 bl[161] br[161] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_162 bl[162] br[162] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_163 bl[163] br[163] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_164 bl[164] br[164] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_165 bl[165] br[165] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_166 bl[166] br[166] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_167 bl[167] br[167] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_168 bl[168] br[168] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_169 bl[169] br[169] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_170 bl[170] br[170] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_171 bl[171] br[171] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_172 bl[172] br[172] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_173 bl[173] br[173] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_174 bl[174] br[174] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_175 bl[175] br[175] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_176 bl[176] br[176] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_177 bl[177] br[177] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_178 bl[178] br[178] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_179 bl[179] br[179] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_180 bl[180] br[180] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_181 bl[181] br[181] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_182 bl[182] br[182] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_183 bl[183] br[183] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_184 bl[184] br[184] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_185 bl[185] br[185] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_186 bl[186] br[186] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_187 bl[187] br[187] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_188 bl[188] br[188] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_189 bl[189] br[189] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_190 bl[190] br[190] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_191 bl[191] br[191] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_192 bl[192] br[192] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_193 bl[193] br[193] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_194 bl[194] br[194] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_195 bl[195] br[195] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_196 bl[196] br[196] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_197 bl[197] br[197] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_198 bl[198] br[198] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_199 bl[199] br[199] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_200 bl[200] br[200] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_201 bl[201] br[201] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_202 bl[202] br[202] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_203 bl[203] br[203] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_204 bl[204] br[204] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_205 bl[205] br[205] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_206 bl[206] br[206] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_207 bl[207] br[207] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_208 bl[208] br[208] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_209 bl[209] br[209] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_210 bl[210] br[210] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_211 bl[211] br[211] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_212 bl[212] br[212] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_213 bl[213] br[213] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_214 bl[214] br[214] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_215 bl[215] br[215] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_216 bl[216] br[216] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_217 bl[217] br[217] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_218 bl[218] br[218] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_219 bl[219] br[219] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_220 bl[220] br[220] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_221 bl[221] br[221] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_222 bl[222] br[222] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_223 bl[223] br[223] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_224 bl[224] br[224] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_225 bl[225] br[225] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_226 bl[226] br[226] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_227 bl[227] br[227] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_228 bl[228] br[228] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_229 bl[229] br[229] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_230 bl[230] br[230] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_231 bl[231] br[231] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_232 bl[232] br[232] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_233 bl[233] br[233] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_234 bl[234] br[234] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_235 bl[235] br[235] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_236 bl[236] br[236] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_237 bl[237] br[237] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_238 bl[238] br[238] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_239 bl[239] br[239] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_240 bl[240] br[240] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_241 bl[241] br[241] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_242 bl[242] br[242] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_243 bl[243] br[243] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_244 bl[244] br[244] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_245 bl[245] br[245] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_246 bl[246] br[246] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_247 bl[247] br[247] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_248 bl[248] br[248] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_249 bl[249] br[249] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_250 bl[250] br[250] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_251 bl[251] br[251] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_252 bl[252] br[252] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_253 bl[253] br[253] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_254 bl[254] br[254] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_255 bl[255] br[255] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_76_0 bl[0] br[0] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_1 bl[1] br[1] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_2 bl[2] br[2] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_3 bl[3] br[3] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_4 bl[4] br[4] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_5 bl[5] br[5] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_6 bl[6] br[6] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_7 bl[7] br[7] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_8 bl[8] br[8] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_9 bl[9] br[9] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_10 bl[10] br[10] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_11 bl[11] br[11] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_12 bl[12] br[12] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_13 bl[13] br[13] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_14 bl[14] br[14] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_15 bl[15] br[15] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_16 bl[16] br[16] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_17 bl[17] br[17] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_18 bl[18] br[18] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_19 bl[19] br[19] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_20 bl[20] br[20] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_21 bl[21] br[21] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_22 bl[22] br[22] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_23 bl[23] br[23] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_24 bl[24] br[24] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_25 bl[25] br[25] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_26 bl[26] br[26] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_27 bl[27] br[27] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_28 bl[28] br[28] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_29 bl[29] br[29] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_30 bl[30] br[30] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_31 bl[31] br[31] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_32 bl[32] br[32] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_33 bl[33] br[33] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_34 bl[34] br[34] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_35 bl[35] br[35] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_36 bl[36] br[36] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_37 bl[37] br[37] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_38 bl[38] br[38] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_39 bl[39] br[39] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_40 bl[40] br[40] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_41 bl[41] br[41] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_42 bl[42] br[42] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_43 bl[43] br[43] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_44 bl[44] br[44] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_45 bl[45] br[45] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_46 bl[46] br[46] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_47 bl[47] br[47] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_48 bl[48] br[48] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_49 bl[49] br[49] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_50 bl[50] br[50] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_51 bl[51] br[51] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_52 bl[52] br[52] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_53 bl[53] br[53] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_54 bl[54] br[54] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_55 bl[55] br[55] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_56 bl[56] br[56] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_57 bl[57] br[57] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_58 bl[58] br[58] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_59 bl[59] br[59] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_60 bl[60] br[60] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_61 bl[61] br[61] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_62 bl[62] br[62] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_63 bl[63] br[63] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_64 bl[64] br[64] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_65 bl[65] br[65] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_66 bl[66] br[66] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_67 bl[67] br[67] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_68 bl[68] br[68] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_69 bl[69] br[69] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_70 bl[70] br[70] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_71 bl[71] br[71] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_72 bl[72] br[72] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_73 bl[73] br[73] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_74 bl[74] br[74] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_75 bl[75] br[75] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_76 bl[76] br[76] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_77 bl[77] br[77] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_78 bl[78] br[78] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_79 bl[79] br[79] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_80 bl[80] br[80] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_81 bl[81] br[81] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_82 bl[82] br[82] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_83 bl[83] br[83] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_84 bl[84] br[84] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_85 bl[85] br[85] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_86 bl[86] br[86] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_87 bl[87] br[87] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_88 bl[88] br[88] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_89 bl[89] br[89] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_90 bl[90] br[90] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_91 bl[91] br[91] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_92 bl[92] br[92] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_93 bl[93] br[93] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_94 bl[94] br[94] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_95 bl[95] br[95] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_96 bl[96] br[96] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_97 bl[97] br[97] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_98 bl[98] br[98] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_99 bl[99] br[99] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_100 bl[100] br[100] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_101 bl[101] br[101] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_102 bl[102] br[102] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_103 bl[103] br[103] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_104 bl[104] br[104] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_105 bl[105] br[105] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_106 bl[106] br[106] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_107 bl[107] br[107] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_108 bl[108] br[108] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_109 bl[109] br[109] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_110 bl[110] br[110] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_111 bl[111] br[111] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_112 bl[112] br[112] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_113 bl[113] br[113] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_114 bl[114] br[114] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_115 bl[115] br[115] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_116 bl[116] br[116] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_117 bl[117] br[117] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_118 bl[118] br[118] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_119 bl[119] br[119] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_120 bl[120] br[120] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_121 bl[121] br[121] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_122 bl[122] br[122] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_123 bl[123] br[123] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_124 bl[124] br[124] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_125 bl[125] br[125] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_126 bl[126] br[126] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_127 bl[127] br[127] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_128 bl[128] br[128] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_129 bl[129] br[129] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_130 bl[130] br[130] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_131 bl[131] br[131] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_132 bl[132] br[132] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_133 bl[133] br[133] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_134 bl[134] br[134] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_135 bl[135] br[135] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_136 bl[136] br[136] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_137 bl[137] br[137] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_138 bl[138] br[138] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_139 bl[139] br[139] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_140 bl[140] br[140] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_141 bl[141] br[141] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_142 bl[142] br[142] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_143 bl[143] br[143] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_144 bl[144] br[144] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_145 bl[145] br[145] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_146 bl[146] br[146] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_147 bl[147] br[147] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_148 bl[148] br[148] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_149 bl[149] br[149] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_150 bl[150] br[150] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_151 bl[151] br[151] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_152 bl[152] br[152] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_153 bl[153] br[153] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_154 bl[154] br[154] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_155 bl[155] br[155] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_156 bl[156] br[156] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_157 bl[157] br[157] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_158 bl[158] br[158] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_159 bl[159] br[159] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_160 bl[160] br[160] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_161 bl[161] br[161] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_162 bl[162] br[162] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_163 bl[163] br[163] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_164 bl[164] br[164] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_165 bl[165] br[165] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_166 bl[166] br[166] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_167 bl[167] br[167] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_168 bl[168] br[168] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_169 bl[169] br[169] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_170 bl[170] br[170] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_171 bl[171] br[171] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_172 bl[172] br[172] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_173 bl[173] br[173] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_174 bl[174] br[174] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_175 bl[175] br[175] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_176 bl[176] br[176] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_177 bl[177] br[177] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_178 bl[178] br[178] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_179 bl[179] br[179] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_180 bl[180] br[180] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_181 bl[181] br[181] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_182 bl[182] br[182] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_183 bl[183] br[183] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_184 bl[184] br[184] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_185 bl[185] br[185] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_186 bl[186] br[186] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_187 bl[187] br[187] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_188 bl[188] br[188] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_189 bl[189] br[189] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_190 bl[190] br[190] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_191 bl[191] br[191] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_192 bl[192] br[192] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_193 bl[193] br[193] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_194 bl[194] br[194] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_195 bl[195] br[195] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_196 bl[196] br[196] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_197 bl[197] br[197] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_198 bl[198] br[198] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_199 bl[199] br[199] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_200 bl[200] br[200] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_201 bl[201] br[201] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_202 bl[202] br[202] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_203 bl[203] br[203] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_204 bl[204] br[204] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_205 bl[205] br[205] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_206 bl[206] br[206] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_207 bl[207] br[207] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_208 bl[208] br[208] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_209 bl[209] br[209] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_210 bl[210] br[210] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_211 bl[211] br[211] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_212 bl[212] br[212] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_213 bl[213] br[213] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_214 bl[214] br[214] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_215 bl[215] br[215] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_216 bl[216] br[216] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_217 bl[217] br[217] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_218 bl[218] br[218] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_219 bl[219] br[219] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_220 bl[220] br[220] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_221 bl[221] br[221] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_222 bl[222] br[222] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_223 bl[223] br[223] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_224 bl[224] br[224] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_225 bl[225] br[225] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_226 bl[226] br[226] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_227 bl[227] br[227] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_228 bl[228] br[228] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_229 bl[229] br[229] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_230 bl[230] br[230] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_231 bl[231] br[231] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_232 bl[232] br[232] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_233 bl[233] br[233] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_234 bl[234] br[234] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_235 bl[235] br[235] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_236 bl[236] br[236] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_237 bl[237] br[237] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_238 bl[238] br[238] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_239 bl[239] br[239] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_240 bl[240] br[240] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_241 bl[241] br[241] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_242 bl[242] br[242] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_243 bl[243] br[243] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_244 bl[244] br[244] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_245 bl[245] br[245] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_246 bl[246] br[246] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_247 bl[247] br[247] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_248 bl[248] br[248] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_249 bl[249] br[249] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_250 bl[250] br[250] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_251 bl[251] br[251] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_252 bl[252] br[252] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_253 bl[253] br[253] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_254 bl[254] br[254] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_255 bl[255] br[255] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_77_0 bl[0] br[0] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_1 bl[1] br[1] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_2 bl[2] br[2] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_3 bl[3] br[3] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_4 bl[4] br[4] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_5 bl[5] br[5] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_6 bl[6] br[6] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_7 bl[7] br[7] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_8 bl[8] br[8] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_9 bl[9] br[9] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_10 bl[10] br[10] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_11 bl[11] br[11] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_12 bl[12] br[12] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_13 bl[13] br[13] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_14 bl[14] br[14] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_15 bl[15] br[15] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_16 bl[16] br[16] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_17 bl[17] br[17] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_18 bl[18] br[18] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_19 bl[19] br[19] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_20 bl[20] br[20] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_21 bl[21] br[21] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_22 bl[22] br[22] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_23 bl[23] br[23] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_24 bl[24] br[24] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_25 bl[25] br[25] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_26 bl[26] br[26] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_27 bl[27] br[27] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_28 bl[28] br[28] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_29 bl[29] br[29] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_30 bl[30] br[30] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_31 bl[31] br[31] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_32 bl[32] br[32] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_33 bl[33] br[33] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_34 bl[34] br[34] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_35 bl[35] br[35] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_36 bl[36] br[36] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_37 bl[37] br[37] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_38 bl[38] br[38] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_39 bl[39] br[39] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_40 bl[40] br[40] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_41 bl[41] br[41] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_42 bl[42] br[42] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_43 bl[43] br[43] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_44 bl[44] br[44] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_45 bl[45] br[45] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_46 bl[46] br[46] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_47 bl[47] br[47] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_48 bl[48] br[48] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_49 bl[49] br[49] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_50 bl[50] br[50] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_51 bl[51] br[51] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_52 bl[52] br[52] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_53 bl[53] br[53] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_54 bl[54] br[54] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_55 bl[55] br[55] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_56 bl[56] br[56] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_57 bl[57] br[57] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_58 bl[58] br[58] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_59 bl[59] br[59] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_60 bl[60] br[60] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_61 bl[61] br[61] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_62 bl[62] br[62] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_63 bl[63] br[63] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_64 bl[64] br[64] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_65 bl[65] br[65] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_66 bl[66] br[66] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_67 bl[67] br[67] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_68 bl[68] br[68] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_69 bl[69] br[69] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_70 bl[70] br[70] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_71 bl[71] br[71] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_72 bl[72] br[72] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_73 bl[73] br[73] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_74 bl[74] br[74] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_75 bl[75] br[75] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_76 bl[76] br[76] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_77 bl[77] br[77] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_78 bl[78] br[78] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_79 bl[79] br[79] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_80 bl[80] br[80] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_81 bl[81] br[81] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_82 bl[82] br[82] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_83 bl[83] br[83] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_84 bl[84] br[84] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_85 bl[85] br[85] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_86 bl[86] br[86] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_87 bl[87] br[87] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_88 bl[88] br[88] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_89 bl[89] br[89] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_90 bl[90] br[90] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_91 bl[91] br[91] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_92 bl[92] br[92] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_93 bl[93] br[93] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_94 bl[94] br[94] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_95 bl[95] br[95] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_96 bl[96] br[96] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_97 bl[97] br[97] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_98 bl[98] br[98] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_99 bl[99] br[99] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_100 bl[100] br[100] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_101 bl[101] br[101] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_102 bl[102] br[102] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_103 bl[103] br[103] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_104 bl[104] br[104] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_105 bl[105] br[105] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_106 bl[106] br[106] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_107 bl[107] br[107] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_108 bl[108] br[108] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_109 bl[109] br[109] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_110 bl[110] br[110] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_111 bl[111] br[111] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_112 bl[112] br[112] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_113 bl[113] br[113] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_114 bl[114] br[114] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_115 bl[115] br[115] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_116 bl[116] br[116] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_117 bl[117] br[117] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_118 bl[118] br[118] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_119 bl[119] br[119] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_120 bl[120] br[120] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_121 bl[121] br[121] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_122 bl[122] br[122] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_123 bl[123] br[123] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_124 bl[124] br[124] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_125 bl[125] br[125] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_126 bl[126] br[126] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_127 bl[127] br[127] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_128 bl[128] br[128] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_129 bl[129] br[129] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_130 bl[130] br[130] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_131 bl[131] br[131] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_132 bl[132] br[132] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_133 bl[133] br[133] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_134 bl[134] br[134] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_135 bl[135] br[135] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_136 bl[136] br[136] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_137 bl[137] br[137] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_138 bl[138] br[138] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_139 bl[139] br[139] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_140 bl[140] br[140] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_141 bl[141] br[141] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_142 bl[142] br[142] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_143 bl[143] br[143] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_144 bl[144] br[144] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_145 bl[145] br[145] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_146 bl[146] br[146] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_147 bl[147] br[147] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_148 bl[148] br[148] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_149 bl[149] br[149] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_150 bl[150] br[150] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_151 bl[151] br[151] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_152 bl[152] br[152] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_153 bl[153] br[153] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_154 bl[154] br[154] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_155 bl[155] br[155] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_156 bl[156] br[156] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_157 bl[157] br[157] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_158 bl[158] br[158] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_159 bl[159] br[159] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_160 bl[160] br[160] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_161 bl[161] br[161] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_162 bl[162] br[162] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_163 bl[163] br[163] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_164 bl[164] br[164] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_165 bl[165] br[165] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_166 bl[166] br[166] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_167 bl[167] br[167] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_168 bl[168] br[168] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_169 bl[169] br[169] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_170 bl[170] br[170] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_171 bl[171] br[171] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_172 bl[172] br[172] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_173 bl[173] br[173] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_174 bl[174] br[174] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_175 bl[175] br[175] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_176 bl[176] br[176] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_177 bl[177] br[177] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_178 bl[178] br[178] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_179 bl[179] br[179] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_180 bl[180] br[180] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_181 bl[181] br[181] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_182 bl[182] br[182] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_183 bl[183] br[183] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_184 bl[184] br[184] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_185 bl[185] br[185] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_186 bl[186] br[186] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_187 bl[187] br[187] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_188 bl[188] br[188] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_189 bl[189] br[189] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_190 bl[190] br[190] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_191 bl[191] br[191] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_192 bl[192] br[192] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_193 bl[193] br[193] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_194 bl[194] br[194] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_195 bl[195] br[195] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_196 bl[196] br[196] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_197 bl[197] br[197] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_198 bl[198] br[198] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_199 bl[199] br[199] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_200 bl[200] br[200] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_201 bl[201] br[201] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_202 bl[202] br[202] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_203 bl[203] br[203] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_204 bl[204] br[204] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_205 bl[205] br[205] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_206 bl[206] br[206] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_207 bl[207] br[207] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_208 bl[208] br[208] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_209 bl[209] br[209] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_210 bl[210] br[210] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_211 bl[211] br[211] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_212 bl[212] br[212] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_213 bl[213] br[213] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_214 bl[214] br[214] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_215 bl[215] br[215] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_216 bl[216] br[216] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_217 bl[217] br[217] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_218 bl[218] br[218] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_219 bl[219] br[219] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_220 bl[220] br[220] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_221 bl[221] br[221] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_222 bl[222] br[222] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_223 bl[223] br[223] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_224 bl[224] br[224] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_225 bl[225] br[225] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_226 bl[226] br[226] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_227 bl[227] br[227] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_228 bl[228] br[228] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_229 bl[229] br[229] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_230 bl[230] br[230] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_231 bl[231] br[231] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_232 bl[232] br[232] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_233 bl[233] br[233] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_234 bl[234] br[234] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_235 bl[235] br[235] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_236 bl[236] br[236] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_237 bl[237] br[237] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_238 bl[238] br[238] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_239 bl[239] br[239] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_240 bl[240] br[240] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_241 bl[241] br[241] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_242 bl[242] br[242] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_243 bl[243] br[243] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_244 bl[244] br[244] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_245 bl[245] br[245] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_246 bl[246] br[246] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_247 bl[247] br[247] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_248 bl[248] br[248] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_249 bl[249] br[249] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_250 bl[250] br[250] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_251 bl[251] br[251] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_252 bl[252] br[252] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_253 bl[253] br[253] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_254 bl[254] br[254] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_255 bl[255] br[255] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_78_0 bl[0] br[0] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_1 bl[1] br[1] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_2 bl[2] br[2] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_3 bl[3] br[3] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_4 bl[4] br[4] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_5 bl[5] br[5] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_6 bl[6] br[6] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_7 bl[7] br[7] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_8 bl[8] br[8] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_9 bl[9] br[9] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_10 bl[10] br[10] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_11 bl[11] br[11] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_12 bl[12] br[12] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_13 bl[13] br[13] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_14 bl[14] br[14] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_15 bl[15] br[15] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_16 bl[16] br[16] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_17 bl[17] br[17] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_18 bl[18] br[18] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_19 bl[19] br[19] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_20 bl[20] br[20] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_21 bl[21] br[21] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_22 bl[22] br[22] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_23 bl[23] br[23] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_24 bl[24] br[24] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_25 bl[25] br[25] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_26 bl[26] br[26] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_27 bl[27] br[27] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_28 bl[28] br[28] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_29 bl[29] br[29] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_30 bl[30] br[30] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_31 bl[31] br[31] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_32 bl[32] br[32] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_33 bl[33] br[33] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_34 bl[34] br[34] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_35 bl[35] br[35] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_36 bl[36] br[36] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_37 bl[37] br[37] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_38 bl[38] br[38] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_39 bl[39] br[39] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_40 bl[40] br[40] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_41 bl[41] br[41] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_42 bl[42] br[42] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_43 bl[43] br[43] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_44 bl[44] br[44] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_45 bl[45] br[45] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_46 bl[46] br[46] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_47 bl[47] br[47] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_48 bl[48] br[48] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_49 bl[49] br[49] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_50 bl[50] br[50] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_51 bl[51] br[51] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_52 bl[52] br[52] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_53 bl[53] br[53] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_54 bl[54] br[54] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_55 bl[55] br[55] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_56 bl[56] br[56] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_57 bl[57] br[57] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_58 bl[58] br[58] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_59 bl[59] br[59] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_60 bl[60] br[60] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_61 bl[61] br[61] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_62 bl[62] br[62] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_63 bl[63] br[63] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_64 bl[64] br[64] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_65 bl[65] br[65] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_66 bl[66] br[66] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_67 bl[67] br[67] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_68 bl[68] br[68] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_69 bl[69] br[69] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_70 bl[70] br[70] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_71 bl[71] br[71] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_72 bl[72] br[72] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_73 bl[73] br[73] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_74 bl[74] br[74] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_75 bl[75] br[75] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_76 bl[76] br[76] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_77 bl[77] br[77] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_78 bl[78] br[78] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_79 bl[79] br[79] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_80 bl[80] br[80] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_81 bl[81] br[81] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_82 bl[82] br[82] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_83 bl[83] br[83] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_84 bl[84] br[84] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_85 bl[85] br[85] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_86 bl[86] br[86] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_87 bl[87] br[87] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_88 bl[88] br[88] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_89 bl[89] br[89] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_90 bl[90] br[90] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_91 bl[91] br[91] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_92 bl[92] br[92] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_93 bl[93] br[93] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_94 bl[94] br[94] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_95 bl[95] br[95] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_96 bl[96] br[96] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_97 bl[97] br[97] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_98 bl[98] br[98] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_99 bl[99] br[99] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_100 bl[100] br[100] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_101 bl[101] br[101] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_102 bl[102] br[102] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_103 bl[103] br[103] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_104 bl[104] br[104] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_105 bl[105] br[105] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_106 bl[106] br[106] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_107 bl[107] br[107] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_108 bl[108] br[108] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_109 bl[109] br[109] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_110 bl[110] br[110] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_111 bl[111] br[111] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_112 bl[112] br[112] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_113 bl[113] br[113] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_114 bl[114] br[114] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_115 bl[115] br[115] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_116 bl[116] br[116] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_117 bl[117] br[117] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_118 bl[118] br[118] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_119 bl[119] br[119] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_120 bl[120] br[120] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_121 bl[121] br[121] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_122 bl[122] br[122] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_123 bl[123] br[123] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_124 bl[124] br[124] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_125 bl[125] br[125] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_126 bl[126] br[126] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_127 bl[127] br[127] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_128 bl[128] br[128] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_129 bl[129] br[129] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_130 bl[130] br[130] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_131 bl[131] br[131] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_132 bl[132] br[132] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_133 bl[133] br[133] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_134 bl[134] br[134] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_135 bl[135] br[135] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_136 bl[136] br[136] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_137 bl[137] br[137] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_138 bl[138] br[138] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_139 bl[139] br[139] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_140 bl[140] br[140] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_141 bl[141] br[141] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_142 bl[142] br[142] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_143 bl[143] br[143] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_144 bl[144] br[144] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_145 bl[145] br[145] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_146 bl[146] br[146] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_147 bl[147] br[147] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_148 bl[148] br[148] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_149 bl[149] br[149] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_150 bl[150] br[150] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_151 bl[151] br[151] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_152 bl[152] br[152] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_153 bl[153] br[153] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_154 bl[154] br[154] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_155 bl[155] br[155] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_156 bl[156] br[156] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_157 bl[157] br[157] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_158 bl[158] br[158] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_159 bl[159] br[159] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_160 bl[160] br[160] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_161 bl[161] br[161] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_162 bl[162] br[162] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_163 bl[163] br[163] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_164 bl[164] br[164] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_165 bl[165] br[165] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_166 bl[166] br[166] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_167 bl[167] br[167] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_168 bl[168] br[168] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_169 bl[169] br[169] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_170 bl[170] br[170] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_171 bl[171] br[171] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_172 bl[172] br[172] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_173 bl[173] br[173] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_174 bl[174] br[174] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_175 bl[175] br[175] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_176 bl[176] br[176] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_177 bl[177] br[177] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_178 bl[178] br[178] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_179 bl[179] br[179] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_180 bl[180] br[180] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_181 bl[181] br[181] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_182 bl[182] br[182] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_183 bl[183] br[183] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_184 bl[184] br[184] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_185 bl[185] br[185] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_186 bl[186] br[186] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_187 bl[187] br[187] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_188 bl[188] br[188] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_189 bl[189] br[189] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_190 bl[190] br[190] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_191 bl[191] br[191] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_192 bl[192] br[192] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_193 bl[193] br[193] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_194 bl[194] br[194] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_195 bl[195] br[195] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_196 bl[196] br[196] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_197 bl[197] br[197] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_198 bl[198] br[198] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_199 bl[199] br[199] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_200 bl[200] br[200] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_201 bl[201] br[201] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_202 bl[202] br[202] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_203 bl[203] br[203] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_204 bl[204] br[204] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_205 bl[205] br[205] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_206 bl[206] br[206] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_207 bl[207] br[207] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_208 bl[208] br[208] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_209 bl[209] br[209] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_210 bl[210] br[210] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_211 bl[211] br[211] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_212 bl[212] br[212] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_213 bl[213] br[213] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_214 bl[214] br[214] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_215 bl[215] br[215] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_216 bl[216] br[216] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_217 bl[217] br[217] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_218 bl[218] br[218] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_219 bl[219] br[219] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_220 bl[220] br[220] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_221 bl[221] br[221] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_222 bl[222] br[222] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_223 bl[223] br[223] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_224 bl[224] br[224] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_225 bl[225] br[225] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_226 bl[226] br[226] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_227 bl[227] br[227] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_228 bl[228] br[228] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_229 bl[229] br[229] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_230 bl[230] br[230] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_231 bl[231] br[231] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_232 bl[232] br[232] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_233 bl[233] br[233] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_234 bl[234] br[234] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_235 bl[235] br[235] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_236 bl[236] br[236] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_237 bl[237] br[237] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_238 bl[238] br[238] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_239 bl[239] br[239] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_240 bl[240] br[240] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_241 bl[241] br[241] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_242 bl[242] br[242] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_243 bl[243] br[243] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_244 bl[244] br[244] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_245 bl[245] br[245] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_246 bl[246] br[246] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_247 bl[247] br[247] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_248 bl[248] br[248] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_249 bl[249] br[249] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_250 bl[250] br[250] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_251 bl[251] br[251] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_252 bl[252] br[252] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_253 bl[253] br[253] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_254 bl[254] br[254] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_255 bl[255] br[255] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_79_0 bl[0] br[0] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_1 bl[1] br[1] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_2 bl[2] br[2] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_3 bl[3] br[3] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_4 bl[4] br[4] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_5 bl[5] br[5] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_6 bl[6] br[6] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_7 bl[7] br[7] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_8 bl[8] br[8] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_9 bl[9] br[9] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_10 bl[10] br[10] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_11 bl[11] br[11] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_12 bl[12] br[12] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_13 bl[13] br[13] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_14 bl[14] br[14] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_15 bl[15] br[15] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_16 bl[16] br[16] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_17 bl[17] br[17] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_18 bl[18] br[18] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_19 bl[19] br[19] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_20 bl[20] br[20] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_21 bl[21] br[21] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_22 bl[22] br[22] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_23 bl[23] br[23] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_24 bl[24] br[24] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_25 bl[25] br[25] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_26 bl[26] br[26] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_27 bl[27] br[27] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_28 bl[28] br[28] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_29 bl[29] br[29] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_30 bl[30] br[30] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_31 bl[31] br[31] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_32 bl[32] br[32] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_33 bl[33] br[33] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_34 bl[34] br[34] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_35 bl[35] br[35] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_36 bl[36] br[36] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_37 bl[37] br[37] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_38 bl[38] br[38] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_39 bl[39] br[39] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_40 bl[40] br[40] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_41 bl[41] br[41] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_42 bl[42] br[42] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_43 bl[43] br[43] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_44 bl[44] br[44] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_45 bl[45] br[45] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_46 bl[46] br[46] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_47 bl[47] br[47] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_48 bl[48] br[48] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_49 bl[49] br[49] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_50 bl[50] br[50] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_51 bl[51] br[51] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_52 bl[52] br[52] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_53 bl[53] br[53] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_54 bl[54] br[54] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_55 bl[55] br[55] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_56 bl[56] br[56] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_57 bl[57] br[57] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_58 bl[58] br[58] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_59 bl[59] br[59] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_60 bl[60] br[60] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_61 bl[61] br[61] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_62 bl[62] br[62] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_63 bl[63] br[63] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_64 bl[64] br[64] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_65 bl[65] br[65] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_66 bl[66] br[66] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_67 bl[67] br[67] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_68 bl[68] br[68] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_69 bl[69] br[69] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_70 bl[70] br[70] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_71 bl[71] br[71] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_72 bl[72] br[72] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_73 bl[73] br[73] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_74 bl[74] br[74] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_75 bl[75] br[75] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_76 bl[76] br[76] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_77 bl[77] br[77] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_78 bl[78] br[78] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_79 bl[79] br[79] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_80 bl[80] br[80] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_81 bl[81] br[81] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_82 bl[82] br[82] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_83 bl[83] br[83] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_84 bl[84] br[84] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_85 bl[85] br[85] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_86 bl[86] br[86] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_87 bl[87] br[87] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_88 bl[88] br[88] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_89 bl[89] br[89] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_90 bl[90] br[90] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_91 bl[91] br[91] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_92 bl[92] br[92] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_93 bl[93] br[93] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_94 bl[94] br[94] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_95 bl[95] br[95] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_96 bl[96] br[96] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_97 bl[97] br[97] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_98 bl[98] br[98] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_99 bl[99] br[99] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_100 bl[100] br[100] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_101 bl[101] br[101] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_102 bl[102] br[102] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_103 bl[103] br[103] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_104 bl[104] br[104] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_105 bl[105] br[105] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_106 bl[106] br[106] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_107 bl[107] br[107] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_108 bl[108] br[108] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_109 bl[109] br[109] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_110 bl[110] br[110] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_111 bl[111] br[111] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_112 bl[112] br[112] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_113 bl[113] br[113] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_114 bl[114] br[114] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_115 bl[115] br[115] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_116 bl[116] br[116] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_117 bl[117] br[117] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_118 bl[118] br[118] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_119 bl[119] br[119] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_120 bl[120] br[120] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_121 bl[121] br[121] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_122 bl[122] br[122] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_123 bl[123] br[123] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_124 bl[124] br[124] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_125 bl[125] br[125] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_126 bl[126] br[126] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_127 bl[127] br[127] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_128 bl[128] br[128] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_129 bl[129] br[129] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_130 bl[130] br[130] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_131 bl[131] br[131] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_132 bl[132] br[132] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_133 bl[133] br[133] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_134 bl[134] br[134] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_135 bl[135] br[135] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_136 bl[136] br[136] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_137 bl[137] br[137] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_138 bl[138] br[138] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_139 bl[139] br[139] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_140 bl[140] br[140] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_141 bl[141] br[141] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_142 bl[142] br[142] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_143 bl[143] br[143] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_144 bl[144] br[144] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_145 bl[145] br[145] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_146 bl[146] br[146] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_147 bl[147] br[147] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_148 bl[148] br[148] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_149 bl[149] br[149] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_150 bl[150] br[150] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_151 bl[151] br[151] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_152 bl[152] br[152] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_153 bl[153] br[153] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_154 bl[154] br[154] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_155 bl[155] br[155] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_156 bl[156] br[156] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_157 bl[157] br[157] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_158 bl[158] br[158] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_159 bl[159] br[159] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_160 bl[160] br[160] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_161 bl[161] br[161] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_162 bl[162] br[162] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_163 bl[163] br[163] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_164 bl[164] br[164] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_165 bl[165] br[165] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_166 bl[166] br[166] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_167 bl[167] br[167] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_168 bl[168] br[168] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_169 bl[169] br[169] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_170 bl[170] br[170] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_171 bl[171] br[171] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_172 bl[172] br[172] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_173 bl[173] br[173] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_174 bl[174] br[174] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_175 bl[175] br[175] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_176 bl[176] br[176] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_177 bl[177] br[177] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_178 bl[178] br[178] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_179 bl[179] br[179] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_180 bl[180] br[180] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_181 bl[181] br[181] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_182 bl[182] br[182] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_183 bl[183] br[183] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_184 bl[184] br[184] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_185 bl[185] br[185] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_186 bl[186] br[186] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_187 bl[187] br[187] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_188 bl[188] br[188] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_189 bl[189] br[189] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_190 bl[190] br[190] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_191 bl[191] br[191] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_192 bl[192] br[192] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_193 bl[193] br[193] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_194 bl[194] br[194] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_195 bl[195] br[195] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_196 bl[196] br[196] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_197 bl[197] br[197] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_198 bl[198] br[198] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_199 bl[199] br[199] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_200 bl[200] br[200] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_201 bl[201] br[201] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_202 bl[202] br[202] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_203 bl[203] br[203] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_204 bl[204] br[204] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_205 bl[205] br[205] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_206 bl[206] br[206] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_207 bl[207] br[207] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_208 bl[208] br[208] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_209 bl[209] br[209] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_210 bl[210] br[210] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_211 bl[211] br[211] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_212 bl[212] br[212] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_213 bl[213] br[213] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_214 bl[214] br[214] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_215 bl[215] br[215] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_216 bl[216] br[216] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_217 bl[217] br[217] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_218 bl[218] br[218] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_219 bl[219] br[219] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_220 bl[220] br[220] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_221 bl[221] br[221] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_222 bl[222] br[222] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_223 bl[223] br[223] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_224 bl[224] br[224] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_225 bl[225] br[225] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_226 bl[226] br[226] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_227 bl[227] br[227] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_228 bl[228] br[228] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_229 bl[229] br[229] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_230 bl[230] br[230] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_231 bl[231] br[231] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_232 bl[232] br[232] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_233 bl[233] br[233] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_234 bl[234] br[234] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_235 bl[235] br[235] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_236 bl[236] br[236] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_237 bl[237] br[237] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_238 bl[238] br[238] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_239 bl[239] br[239] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_240 bl[240] br[240] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_241 bl[241] br[241] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_242 bl[242] br[242] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_243 bl[243] br[243] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_244 bl[244] br[244] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_245 bl[245] br[245] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_246 bl[246] br[246] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_247 bl[247] br[247] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_248 bl[248] br[248] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_249 bl[249] br[249] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_250 bl[250] br[250] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_251 bl[251] br[251] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_252 bl[252] br[252] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_253 bl[253] br[253] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_254 bl[254] br[254] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_255 bl[255] br[255] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_80_0 bl[0] br[0] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_1 bl[1] br[1] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_2 bl[2] br[2] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_3 bl[3] br[3] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_4 bl[4] br[4] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_5 bl[5] br[5] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_6 bl[6] br[6] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_7 bl[7] br[7] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_8 bl[8] br[8] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_9 bl[9] br[9] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_10 bl[10] br[10] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_11 bl[11] br[11] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_12 bl[12] br[12] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_13 bl[13] br[13] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_14 bl[14] br[14] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_15 bl[15] br[15] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_16 bl[16] br[16] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_17 bl[17] br[17] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_18 bl[18] br[18] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_19 bl[19] br[19] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_20 bl[20] br[20] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_21 bl[21] br[21] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_22 bl[22] br[22] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_23 bl[23] br[23] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_24 bl[24] br[24] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_25 bl[25] br[25] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_26 bl[26] br[26] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_27 bl[27] br[27] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_28 bl[28] br[28] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_29 bl[29] br[29] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_30 bl[30] br[30] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_31 bl[31] br[31] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_32 bl[32] br[32] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_33 bl[33] br[33] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_34 bl[34] br[34] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_35 bl[35] br[35] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_36 bl[36] br[36] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_37 bl[37] br[37] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_38 bl[38] br[38] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_39 bl[39] br[39] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_40 bl[40] br[40] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_41 bl[41] br[41] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_42 bl[42] br[42] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_43 bl[43] br[43] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_44 bl[44] br[44] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_45 bl[45] br[45] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_46 bl[46] br[46] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_47 bl[47] br[47] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_48 bl[48] br[48] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_49 bl[49] br[49] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_50 bl[50] br[50] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_51 bl[51] br[51] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_52 bl[52] br[52] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_53 bl[53] br[53] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_54 bl[54] br[54] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_55 bl[55] br[55] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_56 bl[56] br[56] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_57 bl[57] br[57] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_58 bl[58] br[58] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_59 bl[59] br[59] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_60 bl[60] br[60] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_61 bl[61] br[61] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_62 bl[62] br[62] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_63 bl[63] br[63] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_64 bl[64] br[64] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_65 bl[65] br[65] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_66 bl[66] br[66] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_67 bl[67] br[67] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_68 bl[68] br[68] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_69 bl[69] br[69] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_70 bl[70] br[70] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_71 bl[71] br[71] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_72 bl[72] br[72] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_73 bl[73] br[73] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_74 bl[74] br[74] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_75 bl[75] br[75] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_76 bl[76] br[76] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_77 bl[77] br[77] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_78 bl[78] br[78] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_79 bl[79] br[79] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_80 bl[80] br[80] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_81 bl[81] br[81] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_82 bl[82] br[82] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_83 bl[83] br[83] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_84 bl[84] br[84] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_85 bl[85] br[85] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_86 bl[86] br[86] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_87 bl[87] br[87] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_88 bl[88] br[88] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_89 bl[89] br[89] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_90 bl[90] br[90] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_91 bl[91] br[91] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_92 bl[92] br[92] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_93 bl[93] br[93] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_94 bl[94] br[94] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_95 bl[95] br[95] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_96 bl[96] br[96] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_97 bl[97] br[97] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_98 bl[98] br[98] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_99 bl[99] br[99] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_100 bl[100] br[100] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_101 bl[101] br[101] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_102 bl[102] br[102] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_103 bl[103] br[103] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_104 bl[104] br[104] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_105 bl[105] br[105] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_106 bl[106] br[106] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_107 bl[107] br[107] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_108 bl[108] br[108] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_109 bl[109] br[109] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_110 bl[110] br[110] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_111 bl[111] br[111] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_112 bl[112] br[112] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_113 bl[113] br[113] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_114 bl[114] br[114] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_115 bl[115] br[115] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_116 bl[116] br[116] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_117 bl[117] br[117] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_118 bl[118] br[118] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_119 bl[119] br[119] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_120 bl[120] br[120] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_121 bl[121] br[121] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_122 bl[122] br[122] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_123 bl[123] br[123] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_124 bl[124] br[124] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_125 bl[125] br[125] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_126 bl[126] br[126] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_127 bl[127] br[127] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_128 bl[128] br[128] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_129 bl[129] br[129] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_130 bl[130] br[130] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_131 bl[131] br[131] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_132 bl[132] br[132] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_133 bl[133] br[133] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_134 bl[134] br[134] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_135 bl[135] br[135] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_136 bl[136] br[136] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_137 bl[137] br[137] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_138 bl[138] br[138] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_139 bl[139] br[139] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_140 bl[140] br[140] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_141 bl[141] br[141] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_142 bl[142] br[142] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_143 bl[143] br[143] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_144 bl[144] br[144] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_145 bl[145] br[145] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_146 bl[146] br[146] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_147 bl[147] br[147] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_148 bl[148] br[148] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_149 bl[149] br[149] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_150 bl[150] br[150] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_151 bl[151] br[151] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_152 bl[152] br[152] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_153 bl[153] br[153] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_154 bl[154] br[154] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_155 bl[155] br[155] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_156 bl[156] br[156] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_157 bl[157] br[157] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_158 bl[158] br[158] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_159 bl[159] br[159] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_160 bl[160] br[160] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_161 bl[161] br[161] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_162 bl[162] br[162] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_163 bl[163] br[163] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_164 bl[164] br[164] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_165 bl[165] br[165] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_166 bl[166] br[166] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_167 bl[167] br[167] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_168 bl[168] br[168] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_169 bl[169] br[169] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_170 bl[170] br[170] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_171 bl[171] br[171] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_172 bl[172] br[172] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_173 bl[173] br[173] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_174 bl[174] br[174] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_175 bl[175] br[175] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_176 bl[176] br[176] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_177 bl[177] br[177] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_178 bl[178] br[178] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_179 bl[179] br[179] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_180 bl[180] br[180] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_181 bl[181] br[181] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_182 bl[182] br[182] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_183 bl[183] br[183] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_184 bl[184] br[184] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_185 bl[185] br[185] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_186 bl[186] br[186] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_187 bl[187] br[187] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_188 bl[188] br[188] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_189 bl[189] br[189] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_190 bl[190] br[190] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_191 bl[191] br[191] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_192 bl[192] br[192] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_193 bl[193] br[193] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_194 bl[194] br[194] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_195 bl[195] br[195] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_196 bl[196] br[196] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_197 bl[197] br[197] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_198 bl[198] br[198] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_199 bl[199] br[199] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_200 bl[200] br[200] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_201 bl[201] br[201] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_202 bl[202] br[202] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_203 bl[203] br[203] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_204 bl[204] br[204] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_205 bl[205] br[205] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_206 bl[206] br[206] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_207 bl[207] br[207] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_208 bl[208] br[208] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_209 bl[209] br[209] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_210 bl[210] br[210] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_211 bl[211] br[211] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_212 bl[212] br[212] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_213 bl[213] br[213] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_214 bl[214] br[214] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_215 bl[215] br[215] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_216 bl[216] br[216] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_217 bl[217] br[217] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_218 bl[218] br[218] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_219 bl[219] br[219] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_220 bl[220] br[220] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_221 bl[221] br[221] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_222 bl[222] br[222] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_223 bl[223] br[223] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_224 bl[224] br[224] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_225 bl[225] br[225] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_226 bl[226] br[226] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_227 bl[227] br[227] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_228 bl[228] br[228] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_229 bl[229] br[229] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_230 bl[230] br[230] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_231 bl[231] br[231] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_232 bl[232] br[232] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_233 bl[233] br[233] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_234 bl[234] br[234] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_235 bl[235] br[235] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_236 bl[236] br[236] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_237 bl[237] br[237] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_238 bl[238] br[238] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_239 bl[239] br[239] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_240 bl[240] br[240] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_241 bl[241] br[241] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_242 bl[242] br[242] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_243 bl[243] br[243] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_244 bl[244] br[244] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_245 bl[245] br[245] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_246 bl[246] br[246] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_247 bl[247] br[247] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_248 bl[248] br[248] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_249 bl[249] br[249] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_250 bl[250] br[250] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_251 bl[251] br[251] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_252 bl[252] br[252] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_253 bl[253] br[253] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_254 bl[254] br[254] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_255 bl[255] br[255] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_81_0 bl[0] br[0] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_1 bl[1] br[1] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_2 bl[2] br[2] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_3 bl[3] br[3] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_4 bl[4] br[4] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_5 bl[5] br[5] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_6 bl[6] br[6] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_7 bl[7] br[7] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_8 bl[8] br[8] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_9 bl[9] br[9] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_10 bl[10] br[10] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_11 bl[11] br[11] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_12 bl[12] br[12] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_13 bl[13] br[13] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_14 bl[14] br[14] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_15 bl[15] br[15] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_16 bl[16] br[16] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_17 bl[17] br[17] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_18 bl[18] br[18] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_19 bl[19] br[19] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_20 bl[20] br[20] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_21 bl[21] br[21] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_22 bl[22] br[22] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_23 bl[23] br[23] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_24 bl[24] br[24] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_25 bl[25] br[25] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_26 bl[26] br[26] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_27 bl[27] br[27] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_28 bl[28] br[28] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_29 bl[29] br[29] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_30 bl[30] br[30] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_31 bl[31] br[31] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_32 bl[32] br[32] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_33 bl[33] br[33] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_34 bl[34] br[34] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_35 bl[35] br[35] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_36 bl[36] br[36] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_37 bl[37] br[37] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_38 bl[38] br[38] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_39 bl[39] br[39] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_40 bl[40] br[40] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_41 bl[41] br[41] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_42 bl[42] br[42] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_43 bl[43] br[43] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_44 bl[44] br[44] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_45 bl[45] br[45] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_46 bl[46] br[46] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_47 bl[47] br[47] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_48 bl[48] br[48] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_49 bl[49] br[49] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_50 bl[50] br[50] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_51 bl[51] br[51] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_52 bl[52] br[52] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_53 bl[53] br[53] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_54 bl[54] br[54] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_55 bl[55] br[55] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_56 bl[56] br[56] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_57 bl[57] br[57] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_58 bl[58] br[58] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_59 bl[59] br[59] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_60 bl[60] br[60] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_61 bl[61] br[61] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_62 bl[62] br[62] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_63 bl[63] br[63] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_64 bl[64] br[64] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_65 bl[65] br[65] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_66 bl[66] br[66] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_67 bl[67] br[67] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_68 bl[68] br[68] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_69 bl[69] br[69] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_70 bl[70] br[70] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_71 bl[71] br[71] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_72 bl[72] br[72] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_73 bl[73] br[73] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_74 bl[74] br[74] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_75 bl[75] br[75] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_76 bl[76] br[76] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_77 bl[77] br[77] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_78 bl[78] br[78] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_79 bl[79] br[79] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_80 bl[80] br[80] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_81 bl[81] br[81] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_82 bl[82] br[82] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_83 bl[83] br[83] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_84 bl[84] br[84] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_85 bl[85] br[85] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_86 bl[86] br[86] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_87 bl[87] br[87] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_88 bl[88] br[88] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_89 bl[89] br[89] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_90 bl[90] br[90] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_91 bl[91] br[91] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_92 bl[92] br[92] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_93 bl[93] br[93] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_94 bl[94] br[94] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_95 bl[95] br[95] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_96 bl[96] br[96] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_97 bl[97] br[97] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_98 bl[98] br[98] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_99 bl[99] br[99] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_100 bl[100] br[100] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_101 bl[101] br[101] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_102 bl[102] br[102] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_103 bl[103] br[103] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_104 bl[104] br[104] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_105 bl[105] br[105] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_106 bl[106] br[106] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_107 bl[107] br[107] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_108 bl[108] br[108] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_109 bl[109] br[109] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_110 bl[110] br[110] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_111 bl[111] br[111] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_112 bl[112] br[112] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_113 bl[113] br[113] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_114 bl[114] br[114] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_115 bl[115] br[115] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_116 bl[116] br[116] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_117 bl[117] br[117] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_118 bl[118] br[118] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_119 bl[119] br[119] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_120 bl[120] br[120] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_121 bl[121] br[121] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_122 bl[122] br[122] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_123 bl[123] br[123] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_124 bl[124] br[124] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_125 bl[125] br[125] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_126 bl[126] br[126] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_127 bl[127] br[127] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_128 bl[128] br[128] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_129 bl[129] br[129] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_130 bl[130] br[130] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_131 bl[131] br[131] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_132 bl[132] br[132] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_133 bl[133] br[133] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_134 bl[134] br[134] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_135 bl[135] br[135] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_136 bl[136] br[136] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_137 bl[137] br[137] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_138 bl[138] br[138] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_139 bl[139] br[139] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_140 bl[140] br[140] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_141 bl[141] br[141] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_142 bl[142] br[142] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_143 bl[143] br[143] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_144 bl[144] br[144] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_145 bl[145] br[145] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_146 bl[146] br[146] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_147 bl[147] br[147] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_148 bl[148] br[148] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_149 bl[149] br[149] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_150 bl[150] br[150] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_151 bl[151] br[151] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_152 bl[152] br[152] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_153 bl[153] br[153] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_154 bl[154] br[154] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_155 bl[155] br[155] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_156 bl[156] br[156] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_157 bl[157] br[157] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_158 bl[158] br[158] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_159 bl[159] br[159] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_160 bl[160] br[160] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_161 bl[161] br[161] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_162 bl[162] br[162] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_163 bl[163] br[163] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_164 bl[164] br[164] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_165 bl[165] br[165] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_166 bl[166] br[166] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_167 bl[167] br[167] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_168 bl[168] br[168] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_169 bl[169] br[169] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_170 bl[170] br[170] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_171 bl[171] br[171] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_172 bl[172] br[172] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_173 bl[173] br[173] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_174 bl[174] br[174] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_175 bl[175] br[175] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_176 bl[176] br[176] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_177 bl[177] br[177] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_178 bl[178] br[178] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_179 bl[179] br[179] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_180 bl[180] br[180] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_181 bl[181] br[181] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_182 bl[182] br[182] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_183 bl[183] br[183] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_184 bl[184] br[184] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_185 bl[185] br[185] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_186 bl[186] br[186] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_187 bl[187] br[187] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_188 bl[188] br[188] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_189 bl[189] br[189] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_190 bl[190] br[190] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_191 bl[191] br[191] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_192 bl[192] br[192] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_193 bl[193] br[193] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_194 bl[194] br[194] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_195 bl[195] br[195] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_196 bl[196] br[196] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_197 bl[197] br[197] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_198 bl[198] br[198] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_199 bl[199] br[199] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_200 bl[200] br[200] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_201 bl[201] br[201] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_202 bl[202] br[202] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_203 bl[203] br[203] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_204 bl[204] br[204] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_205 bl[205] br[205] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_206 bl[206] br[206] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_207 bl[207] br[207] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_208 bl[208] br[208] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_209 bl[209] br[209] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_210 bl[210] br[210] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_211 bl[211] br[211] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_212 bl[212] br[212] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_213 bl[213] br[213] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_214 bl[214] br[214] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_215 bl[215] br[215] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_216 bl[216] br[216] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_217 bl[217] br[217] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_218 bl[218] br[218] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_219 bl[219] br[219] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_220 bl[220] br[220] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_221 bl[221] br[221] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_222 bl[222] br[222] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_223 bl[223] br[223] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_224 bl[224] br[224] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_225 bl[225] br[225] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_226 bl[226] br[226] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_227 bl[227] br[227] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_228 bl[228] br[228] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_229 bl[229] br[229] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_230 bl[230] br[230] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_231 bl[231] br[231] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_232 bl[232] br[232] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_233 bl[233] br[233] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_234 bl[234] br[234] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_235 bl[235] br[235] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_236 bl[236] br[236] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_237 bl[237] br[237] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_238 bl[238] br[238] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_239 bl[239] br[239] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_240 bl[240] br[240] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_241 bl[241] br[241] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_242 bl[242] br[242] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_243 bl[243] br[243] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_244 bl[244] br[244] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_245 bl[245] br[245] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_246 bl[246] br[246] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_247 bl[247] br[247] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_248 bl[248] br[248] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_249 bl[249] br[249] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_250 bl[250] br[250] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_251 bl[251] br[251] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_252 bl[252] br[252] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_253 bl[253] br[253] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_254 bl[254] br[254] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_255 bl[255] br[255] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_82_0 bl[0] br[0] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_1 bl[1] br[1] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_2 bl[2] br[2] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_3 bl[3] br[3] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_4 bl[4] br[4] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_5 bl[5] br[5] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_6 bl[6] br[6] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_7 bl[7] br[7] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_8 bl[8] br[8] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_9 bl[9] br[9] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_10 bl[10] br[10] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_11 bl[11] br[11] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_12 bl[12] br[12] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_13 bl[13] br[13] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_14 bl[14] br[14] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_15 bl[15] br[15] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_16 bl[16] br[16] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_17 bl[17] br[17] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_18 bl[18] br[18] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_19 bl[19] br[19] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_20 bl[20] br[20] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_21 bl[21] br[21] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_22 bl[22] br[22] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_23 bl[23] br[23] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_24 bl[24] br[24] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_25 bl[25] br[25] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_26 bl[26] br[26] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_27 bl[27] br[27] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_28 bl[28] br[28] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_29 bl[29] br[29] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_30 bl[30] br[30] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_31 bl[31] br[31] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_32 bl[32] br[32] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_33 bl[33] br[33] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_34 bl[34] br[34] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_35 bl[35] br[35] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_36 bl[36] br[36] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_37 bl[37] br[37] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_38 bl[38] br[38] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_39 bl[39] br[39] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_40 bl[40] br[40] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_41 bl[41] br[41] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_42 bl[42] br[42] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_43 bl[43] br[43] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_44 bl[44] br[44] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_45 bl[45] br[45] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_46 bl[46] br[46] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_47 bl[47] br[47] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_48 bl[48] br[48] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_49 bl[49] br[49] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_50 bl[50] br[50] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_51 bl[51] br[51] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_52 bl[52] br[52] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_53 bl[53] br[53] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_54 bl[54] br[54] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_55 bl[55] br[55] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_56 bl[56] br[56] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_57 bl[57] br[57] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_58 bl[58] br[58] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_59 bl[59] br[59] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_60 bl[60] br[60] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_61 bl[61] br[61] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_62 bl[62] br[62] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_63 bl[63] br[63] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_64 bl[64] br[64] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_65 bl[65] br[65] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_66 bl[66] br[66] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_67 bl[67] br[67] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_68 bl[68] br[68] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_69 bl[69] br[69] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_70 bl[70] br[70] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_71 bl[71] br[71] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_72 bl[72] br[72] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_73 bl[73] br[73] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_74 bl[74] br[74] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_75 bl[75] br[75] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_76 bl[76] br[76] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_77 bl[77] br[77] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_78 bl[78] br[78] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_79 bl[79] br[79] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_80 bl[80] br[80] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_81 bl[81] br[81] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_82 bl[82] br[82] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_83 bl[83] br[83] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_84 bl[84] br[84] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_85 bl[85] br[85] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_86 bl[86] br[86] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_87 bl[87] br[87] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_88 bl[88] br[88] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_89 bl[89] br[89] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_90 bl[90] br[90] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_91 bl[91] br[91] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_92 bl[92] br[92] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_93 bl[93] br[93] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_94 bl[94] br[94] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_95 bl[95] br[95] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_96 bl[96] br[96] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_97 bl[97] br[97] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_98 bl[98] br[98] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_99 bl[99] br[99] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_100 bl[100] br[100] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_101 bl[101] br[101] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_102 bl[102] br[102] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_103 bl[103] br[103] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_104 bl[104] br[104] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_105 bl[105] br[105] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_106 bl[106] br[106] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_107 bl[107] br[107] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_108 bl[108] br[108] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_109 bl[109] br[109] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_110 bl[110] br[110] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_111 bl[111] br[111] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_112 bl[112] br[112] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_113 bl[113] br[113] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_114 bl[114] br[114] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_115 bl[115] br[115] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_116 bl[116] br[116] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_117 bl[117] br[117] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_118 bl[118] br[118] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_119 bl[119] br[119] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_120 bl[120] br[120] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_121 bl[121] br[121] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_122 bl[122] br[122] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_123 bl[123] br[123] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_124 bl[124] br[124] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_125 bl[125] br[125] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_126 bl[126] br[126] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_127 bl[127] br[127] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_128 bl[128] br[128] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_129 bl[129] br[129] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_130 bl[130] br[130] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_131 bl[131] br[131] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_132 bl[132] br[132] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_133 bl[133] br[133] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_134 bl[134] br[134] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_135 bl[135] br[135] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_136 bl[136] br[136] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_137 bl[137] br[137] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_138 bl[138] br[138] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_139 bl[139] br[139] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_140 bl[140] br[140] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_141 bl[141] br[141] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_142 bl[142] br[142] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_143 bl[143] br[143] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_144 bl[144] br[144] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_145 bl[145] br[145] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_146 bl[146] br[146] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_147 bl[147] br[147] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_148 bl[148] br[148] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_149 bl[149] br[149] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_150 bl[150] br[150] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_151 bl[151] br[151] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_152 bl[152] br[152] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_153 bl[153] br[153] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_154 bl[154] br[154] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_155 bl[155] br[155] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_156 bl[156] br[156] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_157 bl[157] br[157] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_158 bl[158] br[158] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_159 bl[159] br[159] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_160 bl[160] br[160] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_161 bl[161] br[161] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_162 bl[162] br[162] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_163 bl[163] br[163] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_164 bl[164] br[164] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_165 bl[165] br[165] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_166 bl[166] br[166] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_167 bl[167] br[167] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_168 bl[168] br[168] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_169 bl[169] br[169] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_170 bl[170] br[170] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_171 bl[171] br[171] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_172 bl[172] br[172] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_173 bl[173] br[173] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_174 bl[174] br[174] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_175 bl[175] br[175] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_176 bl[176] br[176] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_177 bl[177] br[177] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_178 bl[178] br[178] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_179 bl[179] br[179] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_180 bl[180] br[180] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_181 bl[181] br[181] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_182 bl[182] br[182] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_183 bl[183] br[183] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_184 bl[184] br[184] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_185 bl[185] br[185] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_186 bl[186] br[186] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_187 bl[187] br[187] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_188 bl[188] br[188] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_189 bl[189] br[189] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_190 bl[190] br[190] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_191 bl[191] br[191] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_192 bl[192] br[192] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_193 bl[193] br[193] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_194 bl[194] br[194] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_195 bl[195] br[195] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_196 bl[196] br[196] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_197 bl[197] br[197] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_198 bl[198] br[198] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_199 bl[199] br[199] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_200 bl[200] br[200] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_201 bl[201] br[201] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_202 bl[202] br[202] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_203 bl[203] br[203] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_204 bl[204] br[204] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_205 bl[205] br[205] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_206 bl[206] br[206] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_207 bl[207] br[207] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_208 bl[208] br[208] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_209 bl[209] br[209] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_210 bl[210] br[210] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_211 bl[211] br[211] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_212 bl[212] br[212] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_213 bl[213] br[213] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_214 bl[214] br[214] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_215 bl[215] br[215] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_216 bl[216] br[216] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_217 bl[217] br[217] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_218 bl[218] br[218] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_219 bl[219] br[219] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_220 bl[220] br[220] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_221 bl[221] br[221] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_222 bl[222] br[222] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_223 bl[223] br[223] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_224 bl[224] br[224] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_225 bl[225] br[225] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_226 bl[226] br[226] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_227 bl[227] br[227] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_228 bl[228] br[228] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_229 bl[229] br[229] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_230 bl[230] br[230] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_231 bl[231] br[231] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_232 bl[232] br[232] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_233 bl[233] br[233] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_234 bl[234] br[234] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_235 bl[235] br[235] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_236 bl[236] br[236] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_237 bl[237] br[237] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_238 bl[238] br[238] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_239 bl[239] br[239] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_240 bl[240] br[240] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_241 bl[241] br[241] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_242 bl[242] br[242] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_243 bl[243] br[243] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_244 bl[244] br[244] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_245 bl[245] br[245] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_246 bl[246] br[246] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_247 bl[247] br[247] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_248 bl[248] br[248] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_249 bl[249] br[249] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_250 bl[250] br[250] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_251 bl[251] br[251] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_252 bl[252] br[252] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_253 bl[253] br[253] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_254 bl[254] br[254] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_255 bl[255] br[255] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_83_0 bl[0] br[0] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_1 bl[1] br[1] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_2 bl[2] br[2] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_3 bl[3] br[3] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_4 bl[4] br[4] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_5 bl[5] br[5] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_6 bl[6] br[6] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_7 bl[7] br[7] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_8 bl[8] br[8] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_9 bl[9] br[9] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_10 bl[10] br[10] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_11 bl[11] br[11] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_12 bl[12] br[12] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_13 bl[13] br[13] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_14 bl[14] br[14] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_15 bl[15] br[15] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_16 bl[16] br[16] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_17 bl[17] br[17] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_18 bl[18] br[18] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_19 bl[19] br[19] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_20 bl[20] br[20] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_21 bl[21] br[21] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_22 bl[22] br[22] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_23 bl[23] br[23] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_24 bl[24] br[24] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_25 bl[25] br[25] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_26 bl[26] br[26] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_27 bl[27] br[27] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_28 bl[28] br[28] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_29 bl[29] br[29] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_30 bl[30] br[30] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_31 bl[31] br[31] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_32 bl[32] br[32] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_33 bl[33] br[33] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_34 bl[34] br[34] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_35 bl[35] br[35] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_36 bl[36] br[36] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_37 bl[37] br[37] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_38 bl[38] br[38] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_39 bl[39] br[39] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_40 bl[40] br[40] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_41 bl[41] br[41] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_42 bl[42] br[42] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_43 bl[43] br[43] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_44 bl[44] br[44] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_45 bl[45] br[45] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_46 bl[46] br[46] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_47 bl[47] br[47] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_48 bl[48] br[48] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_49 bl[49] br[49] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_50 bl[50] br[50] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_51 bl[51] br[51] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_52 bl[52] br[52] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_53 bl[53] br[53] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_54 bl[54] br[54] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_55 bl[55] br[55] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_56 bl[56] br[56] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_57 bl[57] br[57] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_58 bl[58] br[58] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_59 bl[59] br[59] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_60 bl[60] br[60] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_61 bl[61] br[61] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_62 bl[62] br[62] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_63 bl[63] br[63] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_64 bl[64] br[64] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_65 bl[65] br[65] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_66 bl[66] br[66] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_67 bl[67] br[67] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_68 bl[68] br[68] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_69 bl[69] br[69] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_70 bl[70] br[70] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_71 bl[71] br[71] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_72 bl[72] br[72] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_73 bl[73] br[73] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_74 bl[74] br[74] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_75 bl[75] br[75] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_76 bl[76] br[76] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_77 bl[77] br[77] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_78 bl[78] br[78] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_79 bl[79] br[79] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_80 bl[80] br[80] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_81 bl[81] br[81] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_82 bl[82] br[82] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_83 bl[83] br[83] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_84 bl[84] br[84] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_85 bl[85] br[85] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_86 bl[86] br[86] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_87 bl[87] br[87] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_88 bl[88] br[88] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_89 bl[89] br[89] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_90 bl[90] br[90] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_91 bl[91] br[91] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_92 bl[92] br[92] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_93 bl[93] br[93] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_94 bl[94] br[94] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_95 bl[95] br[95] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_96 bl[96] br[96] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_97 bl[97] br[97] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_98 bl[98] br[98] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_99 bl[99] br[99] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_100 bl[100] br[100] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_101 bl[101] br[101] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_102 bl[102] br[102] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_103 bl[103] br[103] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_104 bl[104] br[104] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_105 bl[105] br[105] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_106 bl[106] br[106] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_107 bl[107] br[107] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_108 bl[108] br[108] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_109 bl[109] br[109] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_110 bl[110] br[110] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_111 bl[111] br[111] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_112 bl[112] br[112] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_113 bl[113] br[113] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_114 bl[114] br[114] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_115 bl[115] br[115] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_116 bl[116] br[116] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_117 bl[117] br[117] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_118 bl[118] br[118] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_119 bl[119] br[119] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_120 bl[120] br[120] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_121 bl[121] br[121] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_122 bl[122] br[122] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_123 bl[123] br[123] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_124 bl[124] br[124] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_125 bl[125] br[125] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_126 bl[126] br[126] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_127 bl[127] br[127] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_128 bl[128] br[128] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_129 bl[129] br[129] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_130 bl[130] br[130] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_131 bl[131] br[131] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_132 bl[132] br[132] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_133 bl[133] br[133] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_134 bl[134] br[134] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_135 bl[135] br[135] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_136 bl[136] br[136] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_137 bl[137] br[137] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_138 bl[138] br[138] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_139 bl[139] br[139] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_140 bl[140] br[140] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_141 bl[141] br[141] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_142 bl[142] br[142] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_143 bl[143] br[143] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_144 bl[144] br[144] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_145 bl[145] br[145] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_146 bl[146] br[146] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_147 bl[147] br[147] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_148 bl[148] br[148] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_149 bl[149] br[149] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_150 bl[150] br[150] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_151 bl[151] br[151] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_152 bl[152] br[152] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_153 bl[153] br[153] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_154 bl[154] br[154] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_155 bl[155] br[155] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_156 bl[156] br[156] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_157 bl[157] br[157] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_158 bl[158] br[158] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_159 bl[159] br[159] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_160 bl[160] br[160] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_161 bl[161] br[161] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_162 bl[162] br[162] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_163 bl[163] br[163] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_164 bl[164] br[164] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_165 bl[165] br[165] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_166 bl[166] br[166] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_167 bl[167] br[167] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_168 bl[168] br[168] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_169 bl[169] br[169] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_170 bl[170] br[170] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_171 bl[171] br[171] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_172 bl[172] br[172] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_173 bl[173] br[173] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_174 bl[174] br[174] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_175 bl[175] br[175] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_176 bl[176] br[176] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_177 bl[177] br[177] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_178 bl[178] br[178] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_179 bl[179] br[179] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_180 bl[180] br[180] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_181 bl[181] br[181] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_182 bl[182] br[182] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_183 bl[183] br[183] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_184 bl[184] br[184] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_185 bl[185] br[185] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_186 bl[186] br[186] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_187 bl[187] br[187] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_188 bl[188] br[188] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_189 bl[189] br[189] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_190 bl[190] br[190] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_191 bl[191] br[191] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_192 bl[192] br[192] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_193 bl[193] br[193] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_194 bl[194] br[194] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_195 bl[195] br[195] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_196 bl[196] br[196] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_197 bl[197] br[197] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_198 bl[198] br[198] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_199 bl[199] br[199] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_200 bl[200] br[200] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_201 bl[201] br[201] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_202 bl[202] br[202] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_203 bl[203] br[203] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_204 bl[204] br[204] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_205 bl[205] br[205] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_206 bl[206] br[206] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_207 bl[207] br[207] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_208 bl[208] br[208] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_209 bl[209] br[209] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_210 bl[210] br[210] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_211 bl[211] br[211] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_212 bl[212] br[212] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_213 bl[213] br[213] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_214 bl[214] br[214] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_215 bl[215] br[215] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_216 bl[216] br[216] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_217 bl[217] br[217] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_218 bl[218] br[218] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_219 bl[219] br[219] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_220 bl[220] br[220] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_221 bl[221] br[221] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_222 bl[222] br[222] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_223 bl[223] br[223] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_224 bl[224] br[224] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_225 bl[225] br[225] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_226 bl[226] br[226] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_227 bl[227] br[227] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_228 bl[228] br[228] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_229 bl[229] br[229] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_230 bl[230] br[230] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_231 bl[231] br[231] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_232 bl[232] br[232] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_233 bl[233] br[233] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_234 bl[234] br[234] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_235 bl[235] br[235] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_236 bl[236] br[236] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_237 bl[237] br[237] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_238 bl[238] br[238] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_239 bl[239] br[239] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_240 bl[240] br[240] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_241 bl[241] br[241] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_242 bl[242] br[242] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_243 bl[243] br[243] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_244 bl[244] br[244] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_245 bl[245] br[245] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_246 bl[246] br[246] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_247 bl[247] br[247] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_248 bl[248] br[248] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_249 bl[249] br[249] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_250 bl[250] br[250] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_251 bl[251] br[251] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_252 bl[252] br[252] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_253 bl[253] br[253] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_254 bl[254] br[254] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_255 bl[255] br[255] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_84_0 bl[0] br[0] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_1 bl[1] br[1] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_2 bl[2] br[2] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_3 bl[3] br[3] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_4 bl[4] br[4] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_5 bl[5] br[5] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_6 bl[6] br[6] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_7 bl[7] br[7] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_8 bl[8] br[8] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_9 bl[9] br[9] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_10 bl[10] br[10] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_11 bl[11] br[11] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_12 bl[12] br[12] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_13 bl[13] br[13] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_14 bl[14] br[14] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_15 bl[15] br[15] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_16 bl[16] br[16] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_17 bl[17] br[17] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_18 bl[18] br[18] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_19 bl[19] br[19] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_20 bl[20] br[20] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_21 bl[21] br[21] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_22 bl[22] br[22] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_23 bl[23] br[23] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_24 bl[24] br[24] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_25 bl[25] br[25] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_26 bl[26] br[26] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_27 bl[27] br[27] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_28 bl[28] br[28] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_29 bl[29] br[29] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_30 bl[30] br[30] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_31 bl[31] br[31] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_32 bl[32] br[32] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_33 bl[33] br[33] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_34 bl[34] br[34] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_35 bl[35] br[35] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_36 bl[36] br[36] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_37 bl[37] br[37] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_38 bl[38] br[38] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_39 bl[39] br[39] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_40 bl[40] br[40] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_41 bl[41] br[41] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_42 bl[42] br[42] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_43 bl[43] br[43] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_44 bl[44] br[44] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_45 bl[45] br[45] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_46 bl[46] br[46] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_47 bl[47] br[47] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_48 bl[48] br[48] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_49 bl[49] br[49] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_50 bl[50] br[50] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_51 bl[51] br[51] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_52 bl[52] br[52] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_53 bl[53] br[53] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_54 bl[54] br[54] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_55 bl[55] br[55] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_56 bl[56] br[56] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_57 bl[57] br[57] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_58 bl[58] br[58] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_59 bl[59] br[59] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_60 bl[60] br[60] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_61 bl[61] br[61] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_62 bl[62] br[62] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_63 bl[63] br[63] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_64 bl[64] br[64] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_65 bl[65] br[65] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_66 bl[66] br[66] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_67 bl[67] br[67] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_68 bl[68] br[68] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_69 bl[69] br[69] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_70 bl[70] br[70] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_71 bl[71] br[71] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_72 bl[72] br[72] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_73 bl[73] br[73] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_74 bl[74] br[74] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_75 bl[75] br[75] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_76 bl[76] br[76] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_77 bl[77] br[77] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_78 bl[78] br[78] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_79 bl[79] br[79] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_80 bl[80] br[80] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_81 bl[81] br[81] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_82 bl[82] br[82] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_83 bl[83] br[83] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_84 bl[84] br[84] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_85 bl[85] br[85] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_86 bl[86] br[86] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_87 bl[87] br[87] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_88 bl[88] br[88] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_89 bl[89] br[89] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_90 bl[90] br[90] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_91 bl[91] br[91] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_92 bl[92] br[92] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_93 bl[93] br[93] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_94 bl[94] br[94] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_95 bl[95] br[95] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_96 bl[96] br[96] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_97 bl[97] br[97] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_98 bl[98] br[98] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_99 bl[99] br[99] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_100 bl[100] br[100] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_101 bl[101] br[101] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_102 bl[102] br[102] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_103 bl[103] br[103] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_104 bl[104] br[104] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_105 bl[105] br[105] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_106 bl[106] br[106] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_107 bl[107] br[107] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_108 bl[108] br[108] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_109 bl[109] br[109] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_110 bl[110] br[110] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_111 bl[111] br[111] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_112 bl[112] br[112] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_113 bl[113] br[113] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_114 bl[114] br[114] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_115 bl[115] br[115] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_116 bl[116] br[116] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_117 bl[117] br[117] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_118 bl[118] br[118] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_119 bl[119] br[119] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_120 bl[120] br[120] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_121 bl[121] br[121] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_122 bl[122] br[122] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_123 bl[123] br[123] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_124 bl[124] br[124] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_125 bl[125] br[125] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_126 bl[126] br[126] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_127 bl[127] br[127] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_128 bl[128] br[128] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_129 bl[129] br[129] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_130 bl[130] br[130] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_131 bl[131] br[131] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_132 bl[132] br[132] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_133 bl[133] br[133] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_134 bl[134] br[134] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_135 bl[135] br[135] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_136 bl[136] br[136] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_137 bl[137] br[137] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_138 bl[138] br[138] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_139 bl[139] br[139] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_140 bl[140] br[140] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_141 bl[141] br[141] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_142 bl[142] br[142] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_143 bl[143] br[143] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_144 bl[144] br[144] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_145 bl[145] br[145] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_146 bl[146] br[146] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_147 bl[147] br[147] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_148 bl[148] br[148] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_149 bl[149] br[149] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_150 bl[150] br[150] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_151 bl[151] br[151] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_152 bl[152] br[152] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_153 bl[153] br[153] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_154 bl[154] br[154] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_155 bl[155] br[155] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_156 bl[156] br[156] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_157 bl[157] br[157] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_158 bl[158] br[158] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_159 bl[159] br[159] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_160 bl[160] br[160] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_161 bl[161] br[161] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_162 bl[162] br[162] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_163 bl[163] br[163] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_164 bl[164] br[164] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_165 bl[165] br[165] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_166 bl[166] br[166] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_167 bl[167] br[167] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_168 bl[168] br[168] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_169 bl[169] br[169] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_170 bl[170] br[170] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_171 bl[171] br[171] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_172 bl[172] br[172] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_173 bl[173] br[173] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_174 bl[174] br[174] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_175 bl[175] br[175] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_176 bl[176] br[176] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_177 bl[177] br[177] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_178 bl[178] br[178] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_179 bl[179] br[179] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_180 bl[180] br[180] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_181 bl[181] br[181] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_182 bl[182] br[182] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_183 bl[183] br[183] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_184 bl[184] br[184] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_185 bl[185] br[185] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_186 bl[186] br[186] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_187 bl[187] br[187] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_188 bl[188] br[188] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_189 bl[189] br[189] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_190 bl[190] br[190] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_191 bl[191] br[191] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_192 bl[192] br[192] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_193 bl[193] br[193] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_194 bl[194] br[194] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_195 bl[195] br[195] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_196 bl[196] br[196] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_197 bl[197] br[197] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_198 bl[198] br[198] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_199 bl[199] br[199] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_200 bl[200] br[200] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_201 bl[201] br[201] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_202 bl[202] br[202] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_203 bl[203] br[203] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_204 bl[204] br[204] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_205 bl[205] br[205] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_206 bl[206] br[206] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_207 bl[207] br[207] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_208 bl[208] br[208] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_209 bl[209] br[209] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_210 bl[210] br[210] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_211 bl[211] br[211] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_212 bl[212] br[212] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_213 bl[213] br[213] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_214 bl[214] br[214] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_215 bl[215] br[215] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_216 bl[216] br[216] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_217 bl[217] br[217] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_218 bl[218] br[218] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_219 bl[219] br[219] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_220 bl[220] br[220] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_221 bl[221] br[221] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_222 bl[222] br[222] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_223 bl[223] br[223] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_224 bl[224] br[224] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_225 bl[225] br[225] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_226 bl[226] br[226] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_227 bl[227] br[227] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_228 bl[228] br[228] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_229 bl[229] br[229] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_230 bl[230] br[230] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_231 bl[231] br[231] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_232 bl[232] br[232] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_233 bl[233] br[233] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_234 bl[234] br[234] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_235 bl[235] br[235] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_236 bl[236] br[236] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_237 bl[237] br[237] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_238 bl[238] br[238] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_239 bl[239] br[239] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_240 bl[240] br[240] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_241 bl[241] br[241] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_242 bl[242] br[242] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_243 bl[243] br[243] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_244 bl[244] br[244] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_245 bl[245] br[245] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_246 bl[246] br[246] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_247 bl[247] br[247] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_248 bl[248] br[248] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_249 bl[249] br[249] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_250 bl[250] br[250] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_251 bl[251] br[251] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_252 bl[252] br[252] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_253 bl[253] br[253] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_254 bl[254] br[254] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_255 bl[255] br[255] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_85_0 bl[0] br[0] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_1 bl[1] br[1] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_2 bl[2] br[2] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_3 bl[3] br[3] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_4 bl[4] br[4] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_5 bl[5] br[5] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_6 bl[6] br[6] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_7 bl[7] br[7] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_8 bl[8] br[8] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_9 bl[9] br[9] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_10 bl[10] br[10] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_11 bl[11] br[11] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_12 bl[12] br[12] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_13 bl[13] br[13] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_14 bl[14] br[14] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_15 bl[15] br[15] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_16 bl[16] br[16] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_17 bl[17] br[17] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_18 bl[18] br[18] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_19 bl[19] br[19] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_20 bl[20] br[20] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_21 bl[21] br[21] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_22 bl[22] br[22] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_23 bl[23] br[23] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_24 bl[24] br[24] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_25 bl[25] br[25] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_26 bl[26] br[26] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_27 bl[27] br[27] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_28 bl[28] br[28] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_29 bl[29] br[29] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_30 bl[30] br[30] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_31 bl[31] br[31] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_32 bl[32] br[32] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_33 bl[33] br[33] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_34 bl[34] br[34] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_35 bl[35] br[35] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_36 bl[36] br[36] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_37 bl[37] br[37] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_38 bl[38] br[38] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_39 bl[39] br[39] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_40 bl[40] br[40] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_41 bl[41] br[41] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_42 bl[42] br[42] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_43 bl[43] br[43] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_44 bl[44] br[44] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_45 bl[45] br[45] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_46 bl[46] br[46] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_47 bl[47] br[47] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_48 bl[48] br[48] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_49 bl[49] br[49] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_50 bl[50] br[50] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_51 bl[51] br[51] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_52 bl[52] br[52] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_53 bl[53] br[53] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_54 bl[54] br[54] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_55 bl[55] br[55] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_56 bl[56] br[56] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_57 bl[57] br[57] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_58 bl[58] br[58] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_59 bl[59] br[59] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_60 bl[60] br[60] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_61 bl[61] br[61] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_62 bl[62] br[62] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_63 bl[63] br[63] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_64 bl[64] br[64] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_65 bl[65] br[65] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_66 bl[66] br[66] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_67 bl[67] br[67] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_68 bl[68] br[68] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_69 bl[69] br[69] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_70 bl[70] br[70] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_71 bl[71] br[71] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_72 bl[72] br[72] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_73 bl[73] br[73] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_74 bl[74] br[74] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_75 bl[75] br[75] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_76 bl[76] br[76] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_77 bl[77] br[77] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_78 bl[78] br[78] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_79 bl[79] br[79] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_80 bl[80] br[80] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_81 bl[81] br[81] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_82 bl[82] br[82] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_83 bl[83] br[83] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_84 bl[84] br[84] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_85 bl[85] br[85] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_86 bl[86] br[86] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_87 bl[87] br[87] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_88 bl[88] br[88] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_89 bl[89] br[89] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_90 bl[90] br[90] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_91 bl[91] br[91] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_92 bl[92] br[92] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_93 bl[93] br[93] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_94 bl[94] br[94] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_95 bl[95] br[95] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_96 bl[96] br[96] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_97 bl[97] br[97] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_98 bl[98] br[98] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_99 bl[99] br[99] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_100 bl[100] br[100] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_101 bl[101] br[101] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_102 bl[102] br[102] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_103 bl[103] br[103] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_104 bl[104] br[104] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_105 bl[105] br[105] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_106 bl[106] br[106] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_107 bl[107] br[107] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_108 bl[108] br[108] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_109 bl[109] br[109] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_110 bl[110] br[110] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_111 bl[111] br[111] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_112 bl[112] br[112] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_113 bl[113] br[113] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_114 bl[114] br[114] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_115 bl[115] br[115] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_116 bl[116] br[116] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_117 bl[117] br[117] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_118 bl[118] br[118] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_119 bl[119] br[119] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_120 bl[120] br[120] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_121 bl[121] br[121] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_122 bl[122] br[122] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_123 bl[123] br[123] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_124 bl[124] br[124] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_125 bl[125] br[125] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_126 bl[126] br[126] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_127 bl[127] br[127] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_128 bl[128] br[128] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_129 bl[129] br[129] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_130 bl[130] br[130] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_131 bl[131] br[131] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_132 bl[132] br[132] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_133 bl[133] br[133] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_134 bl[134] br[134] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_135 bl[135] br[135] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_136 bl[136] br[136] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_137 bl[137] br[137] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_138 bl[138] br[138] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_139 bl[139] br[139] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_140 bl[140] br[140] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_141 bl[141] br[141] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_142 bl[142] br[142] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_143 bl[143] br[143] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_144 bl[144] br[144] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_145 bl[145] br[145] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_146 bl[146] br[146] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_147 bl[147] br[147] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_148 bl[148] br[148] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_149 bl[149] br[149] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_150 bl[150] br[150] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_151 bl[151] br[151] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_152 bl[152] br[152] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_153 bl[153] br[153] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_154 bl[154] br[154] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_155 bl[155] br[155] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_156 bl[156] br[156] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_157 bl[157] br[157] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_158 bl[158] br[158] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_159 bl[159] br[159] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_160 bl[160] br[160] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_161 bl[161] br[161] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_162 bl[162] br[162] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_163 bl[163] br[163] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_164 bl[164] br[164] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_165 bl[165] br[165] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_166 bl[166] br[166] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_167 bl[167] br[167] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_168 bl[168] br[168] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_169 bl[169] br[169] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_170 bl[170] br[170] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_171 bl[171] br[171] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_172 bl[172] br[172] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_173 bl[173] br[173] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_174 bl[174] br[174] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_175 bl[175] br[175] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_176 bl[176] br[176] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_177 bl[177] br[177] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_178 bl[178] br[178] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_179 bl[179] br[179] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_180 bl[180] br[180] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_181 bl[181] br[181] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_182 bl[182] br[182] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_183 bl[183] br[183] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_184 bl[184] br[184] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_185 bl[185] br[185] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_186 bl[186] br[186] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_187 bl[187] br[187] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_188 bl[188] br[188] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_189 bl[189] br[189] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_190 bl[190] br[190] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_191 bl[191] br[191] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_192 bl[192] br[192] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_193 bl[193] br[193] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_194 bl[194] br[194] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_195 bl[195] br[195] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_196 bl[196] br[196] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_197 bl[197] br[197] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_198 bl[198] br[198] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_199 bl[199] br[199] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_200 bl[200] br[200] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_201 bl[201] br[201] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_202 bl[202] br[202] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_203 bl[203] br[203] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_204 bl[204] br[204] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_205 bl[205] br[205] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_206 bl[206] br[206] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_207 bl[207] br[207] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_208 bl[208] br[208] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_209 bl[209] br[209] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_210 bl[210] br[210] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_211 bl[211] br[211] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_212 bl[212] br[212] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_213 bl[213] br[213] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_214 bl[214] br[214] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_215 bl[215] br[215] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_216 bl[216] br[216] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_217 bl[217] br[217] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_218 bl[218] br[218] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_219 bl[219] br[219] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_220 bl[220] br[220] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_221 bl[221] br[221] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_222 bl[222] br[222] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_223 bl[223] br[223] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_224 bl[224] br[224] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_225 bl[225] br[225] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_226 bl[226] br[226] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_227 bl[227] br[227] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_228 bl[228] br[228] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_229 bl[229] br[229] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_230 bl[230] br[230] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_231 bl[231] br[231] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_232 bl[232] br[232] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_233 bl[233] br[233] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_234 bl[234] br[234] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_235 bl[235] br[235] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_236 bl[236] br[236] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_237 bl[237] br[237] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_238 bl[238] br[238] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_239 bl[239] br[239] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_240 bl[240] br[240] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_241 bl[241] br[241] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_242 bl[242] br[242] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_243 bl[243] br[243] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_244 bl[244] br[244] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_245 bl[245] br[245] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_246 bl[246] br[246] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_247 bl[247] br[247] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_248 bl[248] br[248] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_249 bl[249] br[249] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_250 bl[250] br[250] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_251 bl[251] br[251] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_252 bl[252] br[252] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_253 bl[253] br[253] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_254 bl[254] br[254] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_255 bl[255] br[255] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_86_0 bl[0] br[0] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_1 bl[1] br[1] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_2 bl[2] br[2] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_3 bl[3] br[3] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_4 bl[4] br[4] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_5 bl[5] br[5] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_6 bl[6] br[6] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_7 bl[7] br[7] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_8 bl[8] br[8] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_9 bl[9] br[9] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_10 bl[10] br[10] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_11 bl[11] br[11] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_12 bl[12] br[12] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_13 bl[13] br[13] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_14 bl[14] br[14] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_15 bl[15] br[15] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_16 bl[16] br[16] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_17 bl[17] br[17] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_18 bl[18] br[18] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_19 bl[19] br[19] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_20 bl[20] br[20] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_21 bl[21] br[21] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_22 bl[22] br[22] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_23 bl[23] br[23] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_24 bl[24] br[24] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_25 bl[25] br[25] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_26 bl[26] br[26] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_27 bl[27] br[27] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_28 bl[28] br[28] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_29 bl[29] br[29] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_30 bl[30] br[30] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_31 bl[31] br[31] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_32 bl[32] br[32] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_33 bl[33] br[33] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_34 bl[34] br[34] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_35 bl[35] br[35] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_36 bl[36] br[36] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_37 bl[37] br[37] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_38 bl[38] br[38] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_39 bl[39] br[39] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_40 bl[40] br[40] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_41 bl[41] br[41] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_42 bl[42] br[42] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_43 bl[43] br[43] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_44 bl[44] br[44] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_45 bl[45] br[45] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_46 bl[46] br[46] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_47 bl[47] br[47] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_48 bl[48] br[48] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_49 bl[49] br[49] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_50 bl[50] br[50] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_51 bl[51] br[51] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_52 bl[52] br[52] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_53 bl[53] br[53] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_54 bl[54] br[54] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_55 bl[55] br[55] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_56 bl[56] br[56] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_57 bl[57] br[57] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_58 bl[58] br[58] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_59 bl[59] br[59] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_60 bl[60] br[60] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_61 bl[61] br[61] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_62 bl[62] br[62] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_63 bl[63] br[63] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_64 bl[64] br[64] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_65 bl[65] br[65] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_66 bl[66] br[66] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_67 bl[67] br[67] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_68 bl[68] br[68] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_69 bl[69] br[69] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_70 bl[70] br[70] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_71 bl[71] br[71] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_72 bl[72] br[72] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_73 bl[73] br[73] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_74 bl[74] br[74] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_75 bl[75] br[75] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_76 bl[76] br[76] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_77 bl[77] br[77] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_78 bl[78] br[78] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_79 bl[79] br[79] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_80 bl[80] br[80] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_81 bl[81] br[81] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_82 bl[82] br[82] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_83 bl[83] br[83] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_84 bl[84] br[84] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_85 bl[85] br[85] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_86 bl[86] br[86] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_87 bl[87] br[87] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_88 bl[88] br[88] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_89 bl[89] br[89] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_90 bl[90] br[90] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_91 bl[91] br[91] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_92 bl[92] br[92] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_93 bl[93] br[93] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_94 bl[94] br[94] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_95 bl[95] br[95] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_96 bl[96] br[96] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_97 bl[97] br[97] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_98 bl[98] br[98] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_99 bl[99] br[99] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_100 bl[100] br[100] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_101 bl[101] br[101] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_102 bl[102] br[102] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_103 bl[103] br[103] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_104 bl[104] br[104] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_105 bl[105] br[105] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_106 bl[106] br[106] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_107 bl[107] br[107] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_108 bl[108] br[108] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_109 bl[109] br[109] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_110 bl[110] br[110] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_111 bl[111] br[111] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_112 bl[112] br[112] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_113 bl[113] br[113] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_114 bl[114] br[114] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_115 bl[115] br[115] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_116 bl[116] br[116] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_117 bl[117] br[117] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_118 bl[118] br[118] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_119 bl[119] br[119] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_120 bl[120] br[120] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_121 bl[121] br[121] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_122 bl[122] br[122] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_123 bl[123] br[123] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_124 bl[124] br[124] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_125 bl[125] br[125] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_126 bl[126] br[126] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_127 bl[127] br[127] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_128 bl[128] br[128] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_129 bl[129] br[129] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_130 bl[130] br[130] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_131 bl[131] br[131] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_132 bl[132] br[132] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_133 bl[133] br[133] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_134 bl[134] br[134] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_135 bl[135] br[135] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_136 bl[136] br[136] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_137 bl[137] br[137] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_138 bl[138] br[138] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_139 bl[139] br[139] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_140 bl[140] br[140] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_141 bl[141] br[141] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_142 bl[142] br[142] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_143 bl[143] br[143] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_144 bl[144] br[144] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_145 bl[145] br[145] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_146 bl[146] br[146] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_147 bl[147] br[147] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_148 bl[148] br[148] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_149 bl[149] br[149] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_150 bl[150] br[150] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_151 bl[151] br[151] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_152 bl[152] br[152] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_153 bl[153] br[153] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_154 bl[154] br[154] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_155 bl[155] br[155] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_156 bl[156] br[156] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_157 bl[157] br[157] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_158 bl[158] br[158] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_159 bl[159] br[159] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_160 bl[160] br[160] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_161 bl[161] br[161] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_162 bl[162] br[162] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_163 bl[163] br[163] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_164 bl[164] br[164] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_165 bl[165] br[165] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_166 bl[166] br[166] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_167 bl[167] br[167] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_168 bl[168] br[168] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_169 bl[169] br[169] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_170 bl[170] br[170] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_171 bl[171] br[171] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_172 bl[172] br[172] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_173 bl[173] br[173] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_174 bl[174] br[174] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_175 bl[175] br[175] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_176 bl[176] br[176] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_177 bl[177] br[177] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_178 bl[178] br[178] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_179 bl[179] br[179] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_180 bl[180] br[180] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_181 bl[181] br[181] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_182 bl[182] br[182] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_183 bl[183] br[183] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_184 bl[184] br[184] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_185 bl[185] br[185] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_186 bl[186] br[186] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_187 bl[187] br[187] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_188 bl[188] br[188] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_189 bl[189] br[189] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_190 bl[190] br[190] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_191 bl[191] br[191] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_192 bl[192] br[192] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_193 bl[193] br[193] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_194 bl[194] br[194] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_195 bl[195] br[195] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_196 bl[196] br[196] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_197 bl[197] br[197] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_198 bl[198] br[198] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_199 bl[199] br[199] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_200 bl[200] br[200] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_201 bl[201] br[201] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_202 bl[202] br[202] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_203 bl[203] br[203] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_204 bl[204] br[204] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_205 bl[205] br[205] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_206 bl[206] br[206] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_207 bl[207] br[207] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_208 bl[208] br[208] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_209 bl[209] br[209] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_210 bl[210] br[210] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_211 bl[211] br[211] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_212 bl[212] br[212] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_213 bl[213] br[213] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_214 bl[214] br[214] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_215 bl[215] br[215] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_216 bl[216] br[216] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_217 bl[217] br[217] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_218 bl[218] br[218] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_219 bl[219] br[219] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_220 bl[220] br[220] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_221 bl[221] br[221] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_222 bl[222] br[222] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_223 bl[223] br[223] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_224 bl[224] br[224] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_225 bl[225] br[225] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_226 bl[226] br[226] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_227 bl[227] br[227] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_228 bl[228] br[228] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_229 bl[229] br[229] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_230 bl[230] br[230] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_231 bl[231] br[231] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_232 bl[232] br[232] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_233 bl[233] br[233] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_234 bl[234] br[234] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_235 bl[235] br[235] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_236 bl[236] br[236] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_237 bl[237] br[237] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_238 bl[238] br[238] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_239 bl[239] br[239] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_240 bl[240] br[240] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_241 bl[241] br[241] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_242 bl[242] br[242] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_243 bl[243] br[243] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_244 bl[244] br[244] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_245 bl[245] br[245] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_246 bl[246] br[246] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_247 bl[247] br[247] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_248 bl[248] br[248] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_249 bl[249] br[249] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_250 bl[250] br[250] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_251 bl[251] br[251] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_252 bl[252] br[252] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_253 bl[253] br[253] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_254 bl[254] br[254] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_255 bl[255] br[255] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_87_0 bl[0] br[0] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_1 bl[1] br[1] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_2 bl[2] br[2] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_3 bl[3] br[3] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_4 bl[4] br[4] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_5 bl[5] br[5] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_6 bl[6] br[6] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_7 bl[7] br[7] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_8 bl[8] br[8] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_9 bl[9] br[9] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_10 bl[10] br[10] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_11 bl[11] br[11] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_12 bl[12] br[12] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_13 bl[13] br[13] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_14 bl[14] br[14] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_15 bl[15] br[15] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_16 bl[16] br[16] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_17 bl[17] br[17] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_18 bl[18] br[18] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_19 bl[19] br[19] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_20 bl[20] br[20] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_21 bl[21] br[21] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_22 bl[22] br[22] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_23 bl[23] br[23] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_24 bl[24] br[24] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_25 bl[25] br[25] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_26 bl[26] br[26] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_27 bl[27] br[27] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_28 bl[28] br[28] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_29 bl[29] br[29] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_30 bl[30] br[30] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_31 bl[31] br[31] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_32 bl[32] br[32] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_33 bl[33] br[33] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_34 bl[34] br[34] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_35 bl[35] br[35] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_36 bl[36] br[36] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_37 bl[37] br[37] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_38 bl[38] br[38] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_39 bl[39] br[39] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_40 bl[40] br[40] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_41 bl[41] br[41] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_42 bl[42] br[42] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_43 bl[43] br[43] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_44 bl[44] br[44] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_45 bl[45] br[45] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_46 bl[46] br[46] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_47 bl[47] br[47] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_48 bl[48] br[48] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_49 bl[49] br[49] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_50 bl[50] br[50] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_51 bl[51] br[51] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_52 bl[52] br[52] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_53 bl[53] br[53] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_54 bl[54] br[54] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_55 bl[55] br[55] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_56 bl[56] br[56] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_57 bl[57] br[57] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_58 bl[58] br[58] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_59 bl[59] br[59] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_60 bl[60] br[60] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_61 bl[61] br[61] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_62 bl[62] br[62] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_63 bl[63] br[63] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_64 bl[64] br[64] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_65 bl[65] br[65] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_66 bl[66] br[66] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_67 bl[67] br[67] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_68 bl[68] br[68] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_69 bl[69] br[69] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_70 bl[70] br[70] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_71 bl[71] br[71] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_72 bl[72] br[72] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_73 bl[73] br[73] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_74 bl[74] br[74] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_75 bl[75] br[75] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_76 bl[76] br[76] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_77 bl[77] br[77] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_78 bl[78] br[78] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_79 bl[79] br[79] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_80 bl[80] br[80] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_81 bl[81] br[81] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_82 bl[82] br[82] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_83 bl[83] br[83] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_84 bl[84] br[84] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_85 bl[85] br[85] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_86 bl[86] br[86] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_87 bl[87] br[87] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_88 bl[88] br[88] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_89 bl[89] br[89] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_90 bl[90] br[90] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_91 bl[91] br[91] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_92 bl[92] br[92] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_93 bl[93] br[93] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_94 bl[94] br[94] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_95 bl[95] br[95] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_96 bl[96] br[96] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_97 bl[97] br[97] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_98 bl[98] br[98] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_99 bl[99] br[99] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_100 bl[100] br[100] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_101 bl[101] br[101] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_102 bl[102] br[102] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_103 bl[103] br[103] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_104 bl[104] br[104] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_105 bl[105] br[105] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_106 bl[106] br[106] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_107 bl[107] br[107] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_108 bl[108] br[108] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_109 bl[109] br[109] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_110 bl[110] br[110] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_111 bl[111] br[111] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_112 bl[112] br[112] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_113 bl[113] br[113] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_114 bl[114] br[114] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_115 bl[115] br[115] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_116 bl[116] br[116] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_117 bl[117] br[117] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_118 bl[118] br[118] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_119 bl[119] br[119] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_120 bl[120] br[120] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_121 bl[121] br[121] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_122 bl[122] br[122] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_123 bl[123] br[123] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_124 bl[124] br[124] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_125 bl[125] br[125] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_126 bl[126] br[126] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_127 bl[127] br[127] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_128 bl[128] br[128] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_129 bl[129] br[129] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_130 bl[130] br[130] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_131 bl[131] br[131] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_132 bl[132] br[132] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_133 bl[133] br[133] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_134 bl[134] br[134] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_135 bl[135] br[135] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_136 bl[136] br[136] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_137 bl[137] br[137] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_138 bl[138] br[138] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_139 bl[139] br[139] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_140 bl[140] br[140] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_141 bl[141] br[141] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_142 bl[142] br[142] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_143 bl[143] br[143] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_144 bl[144] br[144] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_145 bl[145] br[145] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_146 bl[146] br[146] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_147 bl[147] br[147] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_148 bl[148] br[148] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_149 bl[149] br[149] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_150 bl[150] br[150] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_151 bl[151] br[151] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_152 bl[152] br[152] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_153 bl[153] br[153] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_154 bl[154] br[154] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_155 bl[155] br[155] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_156 bl[156] br[156] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_157 bl[157] br[157] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_158 bl[158] br[158] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_159 bl[159] br[159] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_160 bl[160] br[160] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_161 bl[161] br[161] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_162 bl[162] br[162] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_163 bl[163] br[163] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_164 bl[164] br[164] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_165 bl[165] br[165] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_166 bl[166] br[166] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_167 bl[167] br[167] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_168 bl[168] br[168] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_169 bl[169] br[169] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_170 bl[170] br[170] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_171 bl[171] br[171] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_172 bl[172] br[172] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_173 bl[173] br[173] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_174 bl[174] br[174] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_175 bl[175] br[175] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_176 bl[176] br[176] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_177 bl[177] br[177] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_178 bl[178] br[178] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_179 bl[179] br[179] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_180 bl[180] br[180] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_181 bl[181] br[181] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_182 bl[182] br[182] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_183 bl[183] br[183] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_184 bl[184] br[184] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_185 bl[185] br[185] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_186 bl[186] br[186] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_187 bl[187] br[187] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_188 bl[188] br[188] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_189 bl[189] br[189] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_190 bl[190] br[190] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_191 bl[191] br[191] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_192 bl[192] br[192] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_193 bl[193] br[193] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_194 bl[194] br[194] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_195 bl[195] br[195] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_196 bl[196] br[196] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_197 bl[197] br[197] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_198 bl[198] br[198] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_199 bl[199] br[199] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_200 bl[200] br[200] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_201 bl[201] br[201] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_202 bl[202] br[202] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_203 bl[203] br[203] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_204 bl[204] br[204] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_205 bl[205] br[205] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_206 bl[206] br[206] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_207 bl[207] br[207] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_208 bl[208] br[208] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_209 bl[209] br[209] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_210 bl[210] br[210] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_211 bl[211] br[211] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_212 bl[212] br[212] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_213 bl[213] br[213] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_214 bl[214] br[214] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_215 bl[215] br[215] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_216 bl[216] br[216] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_217 bl[217] br[217] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_218 bl[218] br[218] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_219 bl[219] br[219] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_220 bl[220] br[220] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_221 bl[221] br[221] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_222 bl[222] br[222] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_223 bl[223] br[223] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_224 bl[224] br[224] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_225 bl[225] br[225] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_226 bl[226] br[226] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_227 bl[227] br[227] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_228 bl[228] br[228] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_229 bl[229] br[229] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_230 bl[230] br[230] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_231 bl[231] br[231] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_232 bl[232] br[232] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_233 bl[233] br[233] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_234 bl[234] br[234] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_235 bl[235] br[235] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_236 bl[236] br[236] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_237 bl[237] br[237] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_238 bl[238] br[238] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_239 bl[239] br[239] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_240 bl[240] br[240] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_241 bl[241] br[241] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_242 bl[242] br[242] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_243 bl[243] br[243] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_244 bl[244] br[244] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_245 bl[245] br[245] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_246 bl[246] br[246] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_247 bl[247] br[247] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_248 bl[248] br[248] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_249 bl[249] br[249] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_250 bl[250] br[250] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_251 bl[251] br[251] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_252 bl[252] br[252] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_253 bl[253] br[253] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_254 bl[254] br[254] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_255 bl[255] br[255] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_88_0 bl[0] br[0] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_1 bl[1] br[1] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_2 bl[2] br[2] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_3 bl[3] br[3] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_4 bl[4] br[4] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_5 bl[5] br[5] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_6 bl[6] br[6] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_7 bl[7] br[7] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_8 bl[8] br[8] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_9 bl[9] br[9] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_10 bl[10] br[10] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_11 bl[11] br[11] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_12 bl[12] br[12] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_13 bl[13] br[13] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_14 bl[14] br[14] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_15 bl[15] br[15] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_16 bl[16] br[16] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_17 bl[17] br[17] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_18 bl[18] br[18] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_19 bl[19] br[19] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_20 bl[20] br[20] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_21 bl[21] br[21] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_22 bl[22] br[22] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_23 bl[23] br[23] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_24 bl[24] br[24] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_25 bl[25] br[25] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_26 bl[26] br[26] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_27 bl[27] br[27] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_28 bl[28] br[28] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_29 bl[29] br[29] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_30 bl[30] br[30] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_31 bl[31] br[31] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_32 bl[32] br[32] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_33 bl[33] br[33] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_34 bl[34] br[34] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_35 bl[35] br[35] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_36 bl[36] br[36] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_37 bl[37] br[37] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_38 bl[38] br[38] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_39 bl[39] br[39] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_40 bl[40] br[40] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_41 bl[41] br[41] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_42 bl[42] br[42] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_43 bl[43] br[43] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_44 bl[44] br[44] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_45 bl[45] br[45] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_46 bl[46] br[46] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_47 bl[47] br[47] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_48 bl[48] br[48] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_49 bl[49] br[49] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_50 bl[50] br[50] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_51 bl[51] br[51] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_52 bl[52] br[52] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_53 bl[53] br[53] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_54 bl[54] br[54] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_55 bl[55] br[55] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_56 bl[56] br[56] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_57 bl[57] br[57] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_58 bl[58] br[58] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_59 bl[59] br[59] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_60 bl[60] br[60] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_61 bl[61] br[61] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_62 bl[62] br[62] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_63 bl[63] br[63] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_64 bl[64] br[64] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_65 bl[65] br[65] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_66 bl[66] br[66] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_67 bl[67] br[67] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_68 bl[68] br[68] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_69 bl[69] br[69] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_70 bl[70] br[70] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_71 bl[71] br[71] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_72 bl[72] br[72] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_73 bl[73] br[73] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_74 bl[74] br[74] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_75 bl[75] br[75] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_76 bl[76] br[76] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_77 bl[77] br[77] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_78 bl[78] br[78] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_79 bl[79] br[79] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_80 bl[80] br[80] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_81 bl[81] br[81] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_82 bl[82] br[82] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_83 bl[83] br[83] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_84 bl[84] br[84] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_85 bl[85] br[85] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_86 bl[86] br[86] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_87 bl[87] br[87] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_88 bl[88] br[88] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_89 bl[89] br[89] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_90 bl[90] br[90] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_91 bl[91] br[91] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_92 bl[92] br[92] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_93 bl[93] br[93] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_94 bl[94] br[94] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_95 bl[95] br[95] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_96 bl[96] br[96] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_97 bl[97] br[97] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_98 bl[98] br[98] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_99 bl[99] br[99] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_100 bl[100] br[100] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_101 bl[101] br[101] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_102 bl[102] br[102] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_103 bl[103] br[103] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_104 bl[104] br[104] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_105 bl[105] br[105] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_106 bl[106] br[106] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_107 bl[107] br[107] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_108 bl[108] br[108] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_109 bl[109] br[109] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_110 bl[110] br[110] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_111 bl[111] br[111] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_112 bl[112] br[112] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_113 bl[113] br[113] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_114 bl[114] br[114] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_115 bl[115] br[115] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_116 bl[116] br[116] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_117 bl[117] br[117] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_118 bl[118] br[118] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_119 bl[119] br[119] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_120 bl[120] br[120] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_121 bl[121] br[121] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_122 bl[122] br[122] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_123 bl[123] br[123] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_124 bl[124] br[124] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_125 bl[125] br[125] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_126 bl[126] br[126] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_127 bl[127] br[127] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_128 bl[128] br[128] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_129 bl[129] br[129] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_130 bl[130] br[130] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_131 bl[131] br[131] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_132 bl[132] br[132] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_133 bl[133] br[133] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_134 bl[134] br[134] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_135 bl[135] br[135] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_136 bl[136] br[136] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_137 bl[137] br[137] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_138 bl[138] br[138] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_139 bl[139] br[139] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_140 bl[140] br[140] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_141 bl[141] br[141] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_142 bl[142] br[142] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_143 bl[143] br[143] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_144 bl[144] br[144] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_145 bl[145] br[145] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_146 bl[146] br[146] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_147 bl[147] br[147] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_148 bl[148] br[148] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_149 bl[149] br[149] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_150 bl[150] br[150] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_151 bl[151] br[151] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_152 bl[152] br[152] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_153 bl[153] br[153] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_154 bl[154] br[154] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_155 bl[155] br[155] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_156 bl[156] br[156] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_157 bl[157] br[157] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_158 bl[158] br[158] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_159 bl[159] br[159] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_160 bl[160] br[160] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_161 bl[161] br[161] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_162 bl[162] br[162] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_163 bl[163] br[163] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_164 bl[164] br[164] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_165 bl[165] br[165] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_166 bl[166] br[166] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_167 bl[167] br[167] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_168 bl[168] br[168] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_169 bl[169] br[169] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_170 bl[170] br[170] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_171 bl[171] br[171] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_172 bl[172] br[172] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_173 bl[173] br[173] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_174 bl[174] br[174] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_175 bl[175] br[175] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_176 bl[176] br[176] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_177 bl[177] br[177] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_178 bl[178] br[178] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_179 bl[179] br[179] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_180 bl[180] br[180] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_181 bl[181] br[181] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_182 bl[182] br[182] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_183 bl[183] br[183] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_184 bl[184] br[184] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_185 bl[185] br[185] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_186 bl[186] br[186] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_187 bl[187] br[187] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_188 bl[188] br[188] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_189 bl[189] br[189] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_190 bl[190] br[190] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_191 bl[191] br[191] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_192 bl[192] br[192] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_193 bl[193] br[193] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_194 bl[194] br[194] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_195 bl[195] br[195] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_196 bl[196] br[196] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_197 bl[197] br[197] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_198 bl[198] br[198] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_199 bl[199] br[199] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_200 bl[200] br[200] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_201 bl[201] br[201] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_202 bl[202] br[202] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_203 bl[203] br[203] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_204 bl[204] br[204] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_205 bl[205] br[205] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_206 bl[206] br[206] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_207 bl[207] br[207] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_208 bl[208] br[208] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_209 bl[209] br[209] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_210 bl[210] br[210] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_211 bl[211] br[211] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_212 bl[212] br[212] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_213 bl[213] br[213] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_214 bl[214] br[214] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_215 bl[215] br[215] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_216 bl[216] br[216] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_217 bl[217] br[217] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_218 bl[218] br[218] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_219 bl[219] br[219] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_220 bl[220] br[220] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_221 bl[221] br[221] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_222 bl[222] br[222] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_223 bl[223] br[223] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_224 bl[224] br[224] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_225 bl[225] br[225] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_226 bl[226] br[226] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_227 bl[227] br[227] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_228 bl[228] br[228] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_229 bl[229] br[229] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_230 bl[230] br[230] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_231 bl[231] br[231] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_232 bl[232] br[232] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_233 bl[233] br[233] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_234 bl[234] br[234] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_235 bl[235] br[235] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_236 bl[236] br[236] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_237 bl[237] br[237] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_238 bl[238] br[238] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_239 bl[239] br[239] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_240 bl[240] br[240] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_241 bl[241] br[241] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_242 bl[242] br[242] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_243 bl[243] br[243] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_244 bl[244] br[244] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_245 bl[245] br[245] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_246 bl[246] br[246] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_247 bl[247] br[247] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_248 bl[248] br[248] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_249 bl[249] br[249] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_250 bl[250] br[250] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_251 bl[251] br[251] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_252 bl[252] br[252] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_253 bl[253] br[253] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_254 bl[254] br[254] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_255 bl[255] br[255] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_89_0 bl[0] br[0] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_1 bl[1] br[1] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_2 bl[2] br[2] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_3 bl[3] br[3] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_4 bl[4] br[4] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_5 bl[5] br[5] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_6 bl[6] br[6] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_7 bl[7] br[7] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_8 bl[8] br[8] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_9 bl[9] br[9] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_10 bl[10] br[10] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_11 bl[11] br[11] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_12 bl[12] br[12] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_13 bl[13] br[13] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_14 bl[14] br[14] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_15 bl[15] br[15] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_16 bl[16] br[16] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_17 bl[17] br[17] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_18 bl[18] br[18] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_19 bl[19] br[19] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_20 bl[20] br[20] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_21 bl[21] br[21] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_22 bl[22] br[22] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_23 bl[23] br[23] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_24 bl[24] br[24] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_25 bl[25] br[25] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_26 bl[26] br[26] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_27 bl[27] br[27] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_28 bl[28] br[28] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_29 bl[29] br[29] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_30 bl[30] br[30] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_31 bl[31] br[31] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_32 bl[32] br[32] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_33 bl[33] br[33] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_34 bl[34] br[34] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_35 bl[35] br[35] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_36 bl[36] br[36] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_37 bl[37] br[37] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_38 bl[38] br[38] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_39 bl[39] br[39] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_40 bl[40] br[40] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_41 bl[41] br[41] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_42 bl[42] br[42] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_43 bl[43] br[43] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_44 bl[44] br[44] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_45 bl[45] br[45] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_46 bl[46] br[46] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_47 bl[47] br[47] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_48 bl[48] br[48] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_49 bl[49] br[49] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_50 bl[50] br[50] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_51 bl[51] br[51] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_52 bl[52] br[52] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_53 bl[53] br[53] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_54 bl[54] br[54] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_55 bl[55] br[55] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_56 bl[56] br[56] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_57 bl[57] br[57] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_58 bl[58] br[58] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_59 bl[59] br[59] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_60 bl[60] br[60] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_61 bl[61] br[61] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_62 bl[62] br[62] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_63 bl[63] br[63] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_64 bl[64] br[64] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_65 bl[65] br[65] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_66 bl[66] br[66] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_67 bl[67] br[67] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_68 bl[68] br[68] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_69 bl[69] br[69] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_70 bl[70] br[70] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_71 bl[71] br[71] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_72 bl[72] br[72] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_73 bl[73] br[73] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_74 bl[74] br[74] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_75 bl[75] br[75] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_76 bl[76] br[76] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_77 bl[77] br[77] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_78 bl[78] br[78] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_79 bl[79] br[79] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_80 bl[80] br[80] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_81 bl[81] br[81] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_82 bl[82] br[82] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_83 bl[83] br[83] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_84 bl[84] br[84] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_85 bl[85] br[85] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_86 bl[86] br[86] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_87 bl[87] br[87] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_88 bl[88] br[88] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_89 bl[89] br[89] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_90 bl[90] br[90] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_91 bl[91] br[91] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_92 bl[92] br[92] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_93 bl[93] br[93] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_94 bl[94] br[94] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_95 bl[95] br[95] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_96 bl[96] br[96] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_97 bl[97] br[97] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_98 bl[98] br[98] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_99 bl[99] br[99] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_100 bl[100] br[100] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_101 bl[101] br[101] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_102 bl[102] br[102] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_103 bl[103] br[103] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_104 bl[104] br[104] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_105 bl[105] br[105] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_106 bl[106] br[106] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_107 bl[107] br[107] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_108 bl[108] br[108] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_109 bl[109] br[109] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_110 bl[110] br[110] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_111 bl[111] br[111] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_112 bl[112] br[112] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_113 bl[113] br[113] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_114 bl[114] br[114] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_115 bl[115] br[115] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_116 bl[116] br[116] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_117 bl[117] br[117] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_118 bl[118] br[118] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_119 bl[119] br[119] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_120 bl[120] br[120] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_121 bl[121] br[121] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_122 bl[122] br[122] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_123 bl[123] br[123] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_124 bl[124] br[124] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_125 bl[125] br[125] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_126 bl[126] br[126] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_127 bl[127] br[127] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_128 bl[128] br[128] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_129 bl[129] br[129] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_130 bl[130] br[130] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_131 bl[131] br[131] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_132 bl[132] br[132] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_133 bl[133] br[133] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_134 bl[134] br[134] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_135 bl[135] br[135] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_136 bl[136] br[136] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_137 bl[137] br[137] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_138 bl[138] br[138] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_139 bl[139] br[139] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_140 bl[140] br[140] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_141 bl[141] br[141] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_142 bl[142] br[142] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_143 bl[143] br[143] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_144 bl[144] br[144] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_145 bl[145] br[145] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_146 bl[146] br[146] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_147 bl[147] br[147] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_148 bl[148] br[148] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_149 bl[149] br[149] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_150 bl[150] br[150] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_151 bl[151] br[151] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_152 bl[152] br[152] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_153 bl[153] br[153] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_154 bl[154] br[154] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_155 bl[155] br[155] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_156 bl[156] br[156] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_157 bl[157] br[157] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_158 bl[158] br[158] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_159 bl[159] br[159] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_160 bl[160] br[160] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_161 bl[161] br[161] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_162 bl[162] br[162] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_163 bl[163] br[163] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_164 bl[164] br[164] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_165 bl[165] br[165] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_166 bl[166] br[166] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_167 bl[167] br[167] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_168 bl[168] br[168] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_169 bl[169] br[169] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_170 bl[170] br[170] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_171 bl[171] br[171] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_172 bl[172] br[172] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_173 bl[173] br[173] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_174 bl[174] br[174] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_175 bl[175] br[175] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_176 bl[176] br[176] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_177 bl[177] br[177] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_178 bl[178] br[178] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_179 bl[179] br[179] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_180 bl[180] br[180] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_181 bl[181] br[181] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_182 bl[182] br[182] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_183 bl[183] br[183] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_184 bl[184] br[184] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_185 bl[185] br[185] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_186 bl[186] br[186] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_187 bl[187] br[187] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_188 bl[188] br[188] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_189 bl[189] br[189] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_190 bl[190] br[190] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_191 bl[191] br[191] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_192 bl[192] br[192] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_193 bl[193] br[193] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_194 bl[194] br[194] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_195 bl[195] br[195] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_196 bl[196] br[196] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_197 bl[197] br[197] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_198 bl[198] br[198] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_199 bl[199] br[199] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_200 bl[200] br[200] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_201 bl[201] br[201] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_202 bl[202] br[202] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_203 bl[203] br[203] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_204 bl[204] br[204] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_205 bl[205] br[205] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_206 bl[206] br[206] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_207 bl[207] br[207] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_208 bl[208] br[208] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_209 bl[209] br[209] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_210 bl[210] br[210] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_211 bl[211] br[211] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_212 bl[212] br[212] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_213 bl[213] br[213] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_214 bl[214] br[214] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_215 bl[215] br[215] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_216 bl[216] br[216] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_217 bl[217] br[217] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_218 bl[218] br[218] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_219 bl[219] br[219] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_220 bl[220] br[220] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_221 bl[221] br[221] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_222 bl[222] br[222] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_223 bl[223] br[223] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_224 bl[224] br[224] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_225 bl[225] br[225] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_226 bl[226] br[226] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_227 bl[227] br[227] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_228 bl[228] br[228] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_229 bl[229] br[229] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_230 bl[230] br[230] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_231 bl[231] br[231] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_232 bl[232] br[232] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_233 bl[233] br[233] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_234 bl[234] br[234] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_235 bl[235] br[235] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_236 bl[236] br[236] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_237 bl[237] br[237] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_238 bl[238] br[238] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_239 bl[239] br[239] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_240 bl[240] br[240] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_241 bl[241] br[241] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_242 bl[242] br[242] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_243 bl[243] br[243] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_244 bl[244] br[244] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_245 bl[245] br[245] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_246 bl[246] br[246] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_247 bl[247] br[247] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_248 bl[248] br[248] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_249 bl[249] br[249] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_250 bl[250] br[250] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_251 bl[251] br[251] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_252 bl[252] br[252] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_253 bl[253] br[253] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_254 bl[254] br[254] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_255 bl[255] br[255] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_90_0 bl[0] br[0] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_1 bl[1] br[1] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_2 bl[2] br[2] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_3 bl[3] br[3] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_4 bl[4] br[4] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_5 bl[5] br[5] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_6 bl[6] br[6] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_7 bl[7] br[7] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_8 bl[8] br[8] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_9 bl[9] br[9] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_10 bl[10] br[10] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_11 bl[11] br[11] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_12 bl[12] br[12] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_13 bl[13] br[13] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_14 bl[14] br[14] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_15 bl[15] br[15] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_16 bl[16] br[16] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_17 bl[17] br[17] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_18 bl[18] br[18] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_19 bl[19] br[19] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_20 bl[20] br[20] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_21 bl[21] br[21] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_22 bl[22] br[22] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_23 bl[23] br[23] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_24 bl[24] br[24] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_25 bl[25] br[25] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_26 bl[26] br[26] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_27 bl[27] br[27] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_28 bl[28] br[28] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_29 bl[29] br[29] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_30 bl[30] br[30] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_31 bl[31] br[31] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_32 bl[32] br[32] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_33 bl[33] br[33] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_34 bl[34] br[34] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_35 bl[35] br[35] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_36 bl[36] br[36] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_37 bl[37] br[37] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_38 bl[38] br[38] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_39 bl[39] br[39] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_40 bl[40] br[40] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_41 bl[41] br[41] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_42 bl[42] br[42] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_43 bl[43] br[43] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_44 bl[44] br[44] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_45 bl[45] br[45] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_46 bl[46] br[46] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_47 bl[47] br[47] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_48 bl[48] br[48] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_49 bl[49] br[49] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_50 bl[50] br[50] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_51 bl[51] br[51] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_52 bl[52] br[52] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_53 bl[53] br[53] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_54 bl[54] br[54] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_55 bl[55] br[55] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_56 bl[56] br[56] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_57 bl[57] br[57] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_58 bl[58] br[58] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_59 bl[59] br[59] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_60 bl[60] br[60] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_61 bl[61] br[61] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_62 bl[62] br[62] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_63 bl[63] br[63] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_64 bl[64] br[64] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_65 bl[65] br[65] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_66 bl[66] br[66] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_67 bl[67] br[67] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_68 bl[68] br[68] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_69 bl[69] br[69] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_70 bl[70] br[70] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_71 bl[71] br[71] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_72 bl[72] br[72] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_73 bl[73] br[73] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_74 bl[74] br[74] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_75 bl[75] br[75] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_76 bl[76] br[76] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_77 bl[77] br[77] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_78 bl[78] br[78] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_79 bl[79] br[79] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_80 bl[80] br[80] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_81 bl[81] br[81] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_82 bl[82] br[82] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_83 bl[83] br[83] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_84 bl[84] br[84] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_85 bl[85] br[85] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_86 bl[86] br[86] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_87 bl[87] br[87] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_88 bl[88] br[88] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_89 bl[89] br[89] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_90 bl[90] br[90] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_91 bl[91] br[91] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_92 bl[92] br[92] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_93 bl[93] br[93] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_94 bl[94] br[94] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_95 bl[95] br[95] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_96 bl[96] br[96] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_97 bl[97] br[97] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_98 bl[98] br[98] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_99 bl[99] br[99] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_100 bl[100] br[100] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_101 bl[101] br[101] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_102 bl[102] br[102] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_103 bl[103] br[103] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_104 bl[104] br[104] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_105 bl[105] br[105] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_106 bl[106] br[106] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_107 bl[107] br[107] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_108 bl[108] br[108] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_109 bl[109] br[109] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_110 bl[110] br[110] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_111 bl[111] br[111] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_112 bl[112] br[112] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_113 bl[113] br[113] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_114 bl[114] br[114] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_115 bl[115] br[115] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_116 bl[116] br[116] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_117 bl[117] br[117] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_118 bl[118] br[118] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_119 bl[119] br[119] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_120 bl[120] br[120] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_121 bl[121] br[121] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_122 bl[122] br[122] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_123 bl[123] br[123] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_124 bl[124] br[124] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_125 bl[125] br[125] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_126 bl[126] br[126] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_127 bl[127] br[127] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_128 bl[128] br[128] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_129 bl[129] br[129] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_130 bl[130] br[130] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_131 bl[131] br[131] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_132 bl[132] br[132] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_133 bl[133] br[133] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_134 bl[134] br[134] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_135 bl[135] br[135] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_136 bl[136] br[136] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_137 bl[137] br[137] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_138 bl[138] br[138] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_139 bl[139] br[139] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_140 bl[140] br[140] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_141 bl[141] br[141] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_142 bl[142] br[142] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_143 bl[143] br[143] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_144 bl[144] br[144] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_145 bl[145] br[145] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_146 bl[146] br[146] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_147 bl[147] br[147] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_148 bl[148] br[148] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_149 bl[149] br[149] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_150 bl[150] br[150] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_151 bl[151] br[151] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_152 bl[152] br[152] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_153 bl[153] br[153] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_154 bl[154] br[154] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_155 bl[155] br[155] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_156 bl[156] br[156] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_157 bl[157] br[157] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_158 bl[158] br[158] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_159 bl[159] br[159] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_160 bl[160] br[160] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_161 bl[161] br[161] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_162 bl[162] br[162] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_163 bl[163] br[163] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_164 bl[164] br[164] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_165 bl[165] br[165] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_166 bl[166] br[166] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_167 bl[167] br[167] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_168 bl[168] br[168] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_169 bl[169] br[169] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_170 bl[170] br[170] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_171 bl[171] br[171] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_172 bl[172] br[172] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_173 bl[173] br[173] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_174 bl[174] br[174] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_175 bl[175] br[175] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_176 bl[176] br[176] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_177 bl[177] br[177] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_178 bl[178] br[178] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_179 bl[179] br[179] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_180 bl[180] br[180] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_181 bl[181] br[181] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_182 bl[182] br[182] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_183 bl[183] br[183] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_184 bl[184] br[184] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_185 bl[185] br[185] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_186 bl[186] br[186] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_187 bl[187] br[187] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_188 bl[188] br[188] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_189 bl[189] br[189] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_190 bl[190] br[190] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_191 bl[191] br[191] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_192 bl[192] br[192] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_193 bl[193] br[193] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_194 bl[194] br[194] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_195 bl[195] br[195] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_196 bl[196] br[196] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_197 bl[197] br[197] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_198 bl[198] br[198] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_199 bl[199] br[199] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_200 bl[200] br[200] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_201 bl[201] br[201] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_202 bl[202] br[202] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_203 bl[203] br[203] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_204 bl[204] br[204] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_205 bl[205] br[205] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_206 bl[206] br[206] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_207 bl[207] br[207] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_208 bl[208] br[208] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_209 bl[209] br[209] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_210 bl[210] br[210] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_211 bl[211] br[211] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_212 bl[212] br[212] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_213 bl[213] br[213] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_214 bl[214] br[214] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_215 bl[215] br[215] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_216 bl[216] br[216] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_217 bl[217] br[217] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_218 bl[218] br[218] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_219 bl[219] br[219] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_220 bl[220] br[220] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_221 bl[221] br[221] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_222 bl[222] br[222] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_223 bl[223] br[223] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_224 bl[224] br[224] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_225 bl[225] br[225] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_226 bl[226] br[226] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_227 bl[227] br[227] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_228 bl[228] br[228] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_229 bl[229] br[229] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_230 bl[230] br[230] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_231 bl[231] br[231] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_232 bl[232] br[232] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_233 bl[233] br[233] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_234 bl[234] br[234] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_235 bl[235] br[235] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_236 bl[236] br[236] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_237 bl[237] br[237] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_238 bl[238] br[238] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_239 bl[239] br[239] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_240 bl[240] br[240] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_241 bl[241] br[241] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_242 bl[242] br[242] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_243 bl[243] br[243] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_244 bl[244] br[244] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_245 bl[245] br[245] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_246 bl[246] br[246] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_247 bl[247] br[247] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_248 bl[248] br[248] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_249 bl[249] br[249] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_250 bl[250] br[250] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_251 bl[251] br[251] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_252 bl[252] br[252] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_253 bl[253] br[253] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_254 bl[254] br[254] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_255 bl[255] br[255] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_91_0 bl[0] br[0] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_1 bl[1] br[1] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_2 bl[2] br[2] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_3 bl[3] br[3] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_4 bl[4] br[4] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_5 bl[5] br[5] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_6 bl[6] br[6] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_7 bl[7] br[7] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_8 bl[8] br[8] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_9 bl[9] br[9] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_10 bl[10] br[10] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_11 bl[11] br[11] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_12 bl[12] br[12] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_13 bl[13] br[13] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_14 bl[14] br[14] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_15 bl[15] br[15] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_16 bl[16] br[16] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_17 bl[17] br[17] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_18 bl[18] br[18] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_19 bl[19] br[19] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_20 bl[20] br[20] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_21 bl[21] br[21] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_22 bl[22] br[22] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_23 bl[23] br[23] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_24 bl[24] br[24] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_25 bl[25] br[25] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_26 bl[26] br[26] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_27 bl[27] br[27] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_28 bl[28] br[28] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_29 bl[29] br[29] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_30 bl[30] br[30] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_31 bl[31] br[31] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_32 bl[32] br[32] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_33 bl[33] br[33] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_34 bl[34] br[34] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_35 bl[35] br[35] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_36 bl[36] br[36] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_37 bl[37] br[37] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_38 bl[38] br[38] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_39 bl[39] br[39] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_40 bl[40] br[40] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_41 bl[41] br[41] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_42 bl[42] br[42] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_43 bl[43] br[43] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_44 bl[44] br[44] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_45 bl[45] br[45] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_46 bl[46] br[46] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_47 bl[47] br[47] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_48 bl[48] br[48] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_49 bl[49] br[49] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_50 bl[50] br[50] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_51 bl[51] br[51] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_52 bl[52] br[52] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_53 bl[53] br[53] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_54 bl[54] br[54] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_55 bl[55] br[55] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_56 bl[56] br[56] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_57 bl[57] br[57] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_58 bl[58] br[58] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_59 bl[59] br[59] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_60 bl[60] br[60] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_61 bl[61] br[61] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_62 bl[62] br[62] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_63 bl[63] br[63] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_64 bl[64] br[64] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_65 bl[65] br[65] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_66 bl[66] br[66] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_67 bl[67] br[67] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_68 bl[68] br[68] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_69 bl[69] br[69] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_70 bl[70] br[70] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_71 bl[71] br[71] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_72 bl[72] br[72] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_73 bl[73] br[73] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_74 bl[74] br[74] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_75 bl[75] br[75] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_76 bl[76] br[76] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_77 bl[77] br[77] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_78 bl[78] br[78] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_79 bl[79] br[79] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_80 bl[80] br[80] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_81 bl[81] br[81] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_82 bl[82] br[82] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_83 bl[83] br[83] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_84 bl[84] br[84] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_85 bl[85] br[85] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_86 bl[86] br[86] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_87 bl[87] br[87] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_88 bl[88] br[88] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_89 bl[89] br[89] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_90 bl[90] br[90] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_91 bl[91] br[91] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_92 bl[92] br[92] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_93 bl[93] br[93] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_94 bl[94] br[94] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_95 bl[95] br[95] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_96 bl[96] br[96] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_97 bl[97] br[97] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_98 bl[98] br[98] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_99 bl[99] br[99] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_100 bl[100] br[100] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_101 bl[101] br[101] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_102 bl[102] br[102] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_103 bl[103] br[103] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_104 bl[104] br[104] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_105 bl[105] br[105] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_106 bl[106] br[106] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_107 bl[107] br[107] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_108 bl[108] br[108] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_109 bl[109] br[109] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_110 bl[110] br[110] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_111 bl[111] br[111] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_112 bl[112] br[112] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_113 bl[113] br[113] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_114 bl[114] br[114] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_115 bl[115] br[115] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_116 bl[116] br[116] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_117 bl[117] br[117] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_118 bl[118] br[118] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_119 bl[119] br[119] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_120 bl[120] br[120] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_121 bl[121] br[121] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_122 bl[122] br[122] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_123 bl[123] br[123] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_124 bl[124] br[124] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_125 bl[125] br[125] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_126 bl[126] br[126] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_127 bl[127] br[127] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_128 bl[128] br[128] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_129 bl[129] br[129] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_130 bl[130] br[130] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_131 bl[131] br[131] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_132 bl[132] br[132] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_133 bl[133] br[133] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_134 bl[134] br[134] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_135 bl[135] br[135] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_136 bl[136] br[136] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_137 bl[137] br[137] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_138 bl[138] br[138] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_139 bl[139] br[139] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_140 bl[140] br[140] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_141 bl[141] br[141] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_142 bl[142] br[142] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_143 bl[143] br[143] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_144 bl[144] br[144] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_145 bl[145] br[145] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_146 bl[146] br[146] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_147 bl[147] br[147] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_148 bl[148] br[148] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_149 bl[149] br[149] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_150 bl[150] br[150] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_151 bl[151] br[151] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_152 bl[152] br[152] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_153 bl[153] br[153] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_154 bl[154] br[154] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_155 bl[155] br[155] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_156 bl[156] br[156] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_157 bl[157] br[157] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_158 bl[158] br[158] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_159 bl[159] br[159] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_160 bl[160] br[160] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_161 bl[161] br[161] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_162 bl[162] br[162] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_163 bl[163] br[163] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_164 bl[164] br[164] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_165 bl[165] br[165] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_166 bl[166] br[166] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_167 bl[167] br[167] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_168 bl[168] br[168] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_169 bl[169] br[169] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_170 bl[170] br[170] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_171 bl[171] br[171] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_172 bl[172] br[172] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_173 bl[173] br[173] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_174 bl[174] br[174] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_175 bl[175] br[175] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_176 bl[176] br[176] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_177 bl[177] br[177] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_178 bl[178] br[178] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_179 bl[179] br[179] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_180 bl[180] br[180] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_181 bl[181] br[181] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_182 bl[182] br[182] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_183 bl[183] br[183] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_184 bl[184] br[184] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_185 bl[185] br[185] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_186 bl[186] br[186] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_187 bl[187] br[187] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_188 bl[188] br[188] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_189 bl[189] br[189] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_190 bl[190] br[190] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_191 bl[191] br[191] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_192 bl[192] br[192] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_193 bl[193] br[193] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_194 bl[194] br[194] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_195 bl[195] br[195] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_196 bl[196] br[196] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_197 bl[197] br[197] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_198 bl[198] br[198] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_199 bl[199] br[199] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_200 bl[200] br[200] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_201 bl[201] br[201] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_202 bl[202] br[202] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_203 bl[203] br[203] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_204 bl[204] br[204] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_205 bl[205] br[205] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_206 bl[206] br[206] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_207 bl[207] br[207] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_208 bl[208] br[208] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_209 bl[209] br[209] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_210 bl[210] br[210] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_211 bl[211] br[211] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_212 bl[212] br[212] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_213 bl[213] br[213] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_214 bl[214] br[214] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_215 bl[215] br[215] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_216 bl[216] br[216] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_217 bl[217] br[217] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_218 bl[218] br[218] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_219 bl[219] br[219] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_220 bl[220] br[220] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_221 bl[221] br[221] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_222 bl[222] br[222] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_223 bl[223] br[223] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_224 bl[224] br[224] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_225 bl[225] br[225] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_226 bl[226] br[226] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_227 bl[227] br[227] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_228 bl[228] br[228] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_229 bl[229] br[229] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_230 bl[230] br[230] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_231 bl[231] br[231] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_232 bl[232] br[232] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_233 bl[233] br[233] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_234 bl[234] br[234] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_235 bl[235] br[235] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_236 bl[236] br[236] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_237 bl[237] br[237] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_238 bl[238] br[238] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_239 bl[239] br[239] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_240 bl[240] br[240] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_241 bl[241] br[241] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_242 bl[242] br[242] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_243 bl[243] br[243] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_244 bl[244] br[244] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_245 bl[245] br[245] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_246 bl[246] br[246] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_247 bl[247] br[247] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_248 bl[248] br[248] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_249 bl[249] br[249] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_250 bl[250] br[250] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_251 bl[251] br[251] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_252 bl[252] br[252] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_253 bl[253] br[253] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_254 bl[254] br[254] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_255 bl[255] br[255] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_92_0 bl[0] br[0] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_1 bl[1] br[1] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_2 bl[2] br[2] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_3 bl[3] br[3] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_4 bl[4] br[4] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_5 bl[5] br[5] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_6 bl[6] br[6] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_7 bl[7] br[7] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_8 bl[8] br[8] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_9 bl[9] br[9] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_10 bl[10] br[10] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_11 bl[11] br[11] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_12 bl[12] br[12] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_13 bl[13] br[13] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_14 bl[14] br[14] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_15 bl[15] br[15] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_16 bl[16] br[16] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_17 bl[17] br[17] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_18 bl[18] br[18] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_19 bl[19] br[19] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_20 bl[20] br[20] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_21 bl[21] br[21] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_22 bl[22] br[22] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_23 bl[23] br[23] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_24 bl[24] br[24] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_25 bl[25] br[25] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_26 bl[26] br[26] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_27 bl[27] br[27] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_28 bl[28] br[28] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_29 bl[29] br[29] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_30 bl[30] br[30] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_31 bl[31] br[31] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_32 bl[32] br[32] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_33 bl[33] br[33] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_34 bl[34] br[34] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_35 bl[35] br[35] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_36 bl[36] br[36] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_37 bl[37] br[37] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_38 bl[38] br[38] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_39 bl[39] br[39] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_40 bl[40] br[40] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_41 bl[41] br[41] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_42 bl[42] br[42] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_43 bl[43] br[43] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_44 bl[44] br[44] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_45 bl[45] br[45] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_46 bl[46] br[46] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_47 bl[47] br[47] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_48 bl[48] br[48] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_49 bl[49] br[49] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_50 bl[50] br[50] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_51 bl[51] br[51] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_52 bl[52] br[52] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_53 bl[53] br[53] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_54 bl[54] br[54] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_55 bl[55] br[55] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_56 bl[56] br[56] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_57 bl[57] br[57] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_58 bl[58] br[58] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_59 bl[59] br[59] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_60 bl[60] br[60] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_61 bl[61] br[61] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_62 bl[62] br[62] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_63 bl[63] br[63] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_64 bl[64] br[64] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_65 bl[65] br[65] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_66 bl[66] br[66] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_67 bl[67] br[67] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_68 bl[68] br[68] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_69 bl[69] br[69] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_70 bl[70] br[70] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_71 bl[71] br[71] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_72 bl[72] br[72] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_73 bl[73] br[73] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_74 bl[74] br[74] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_75 bl[75] br[75] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_76 bl[76] br[76] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_77 bl[77] br[77] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_78 bl[78] br[78] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_79 bl[79] br[79] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_80 bl[80] br[80] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_81 bl[81] br[81] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_82 bl[82] br[82] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_83 bl[83] br[83] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_84 bl[84] br[84] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_85 bl[85] br[85] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_86 bl[86] br[86] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_87 bl[87] br[87] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_88 bl[88] br[88] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_89 bl[89] br[89] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_90 bl[90] br[90] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_91 bl[91] br[91] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_92 bl[92] br[92] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_93 bl[93] br[93] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_94 bl[94] br[94] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_95 bl[95] br[95] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_96 bl[96] br[96] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_97 bl[97] br[97] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_98 bl[98] br[98] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_99 bl[99] br[99] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_100 bl[100] br[100] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_101 bl[101] br[101] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_102 bl[102] br[102] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_103 bl[103] br[103] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_104 bl[104] br[104] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_105 bl[105] br[105] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_106 bl[106] br[106] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_107 bl[107] br[107] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_108 bl[108] br[108] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_109 bl[109] br[109] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_110 bl[110] br[110] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_111 bl[111] br[111] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_112 bl[112] br[112] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_113 bl[113] br[113] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_114 bl[114] br[114] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_115 bl[115] br[115] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_116 bl[116] br[116] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_117 bl[117] br[117] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_118 bl[118] br[118] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_119 bl[119] br[119] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_120 bl[120] br[120] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_121 bl[121] br[121] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_122 bl[122] br[122] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_123 bl[123] br[123] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_124 bl[124] br[124] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_125 bl[125] br[125] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_126 bl[126] br[126] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_127 bl[127] br[127] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_128 bl[128] br[128] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_129 bl[129] br[129] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_130 bl[130] br[130] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_131 bl[131] br[131] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_132 bl[132] br[132] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_133 bl[133] br[133] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_134 bl[134] br[134] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_135 bl[135] br[135] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_136 bl[136] br[136] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_137 bl[137] br[137] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_138 bl[138] br[138] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_139 bl[139] br[139] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_140 bl[140] br[140] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_141 bl[141] br[141] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_142 bl[142] br[142] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_143 bl[143] br[143] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_144 bl[144] br[144] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_145 bl[145] br[145] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_146 bl[146] br[146] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_147 bl[147] br[147] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_148 bl[148] br[148] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_149 bl[149] br[149] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_150 bl[150] br[150] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_151 bl[151] br[151] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_152 bl[152] br[152] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_153 bl[153] br[153] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_154 bl[154] br[154] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_155 bl[155] br[155] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_156 bl[156] br[156] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_157 bl[157] br[157] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_158 bl[158] br[158] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_159 bl[159] br[159] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_160 bl[160] br[160] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_161 bl[161] br[161] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_162 bl[162] br[162] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_163 bl[163] br[163] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_164 bl[164] br[164] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_165 bl[165] br[165] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_166 bl[166] br[166] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_167 bl[167] br[167] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_168 bl[168] br[168] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_169 bl[169] br[169] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_170 bl[170] br[170] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_171 bl[171] br[171] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_172 bl[172] br[172] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_173 bl[173] br[173] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_174 bl[174] br[174] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_175 bl[175] br[175] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_176 bl[176] br[176] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_177 bl[177] br[177] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_178 bl[178] br[178] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_179 bl[179] br[179] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_180 bl[180] br[180] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_181 bl[181] br[181] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_182 bl[182] br[182] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_183 bl[183] br[183] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_184 bl[184] br[184] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_185 bl[185] br[185] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_186 bl[186] br[186] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_187 bl[187] br[187] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_188 bl[188] br[188] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_189 bl[189] br[189] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_190 bl[190] br[190] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_191 bl[191] br[191] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_192 bl[192] br[192] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_193 bl[193] br[193] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_194 bl[194] br[194] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_195 bl[195] br[195] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_196 bl[196] br[196] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_197 bl[197] br[197] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_198 bl[198] br[198] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_199 bl[199] br[199] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_200 bl[200] br[200] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_201 bl[201] br[201] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_202 bl[202] br[202] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_203 bl[203] br[203] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_204 bl[204] br[204] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_205 bl[205] br[205] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_206 bl[206] br[206] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_207 bl[207] br[207] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_208 bl[208] br[208] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_209 bl[209] br[209] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_210 bl[210] br[210] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_211 bl[211] br[211] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_212 bl[212] br[212] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_213 bl[213] br[213] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_214 bl[214] br[214] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_215 bl[215] br[215] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_216 bl[216] br[216] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_217 bl[217] br[217] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_218 bl[218] br[218] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_219 bl[219] br[219] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_220 bl[220] br[220] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_221 bl[221] br[221] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_222 bl[222] br[222] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_223 bl[223] br[223] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_224 bl[224] br[224] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_225 bl[225] br[225] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_226 bl[226] br[226] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_227 bl[227] br[227] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_228 bl[228] br[228] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_229 bl[229] br[229] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_230 bl[230] br[230] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_231 bl[231] br[231] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_232 bl[232] br[232] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_233 bl[233] br[233] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_234 bl[234] br[234] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_235 bl[235] br[235] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_236 bl[236] br[236] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_237 bl[237] br[237] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_238 bl[238] br[238] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_239 bl[239] br[239] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_240 bl[240] br[240] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_241 bl[241] br[241] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_242 bl[242] br[242] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_243 bl[243] br[243] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_244 bl[244] br[244] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_245 bl[245] br[245] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_246 bl[246] br[246] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_247 bl[247] br[247] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_248 bl[248] br[248] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_249 bl[249] br[249] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_250 bl[250] br[250] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_251 bl[251] br[251] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_252 bl[252] br[252] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_253 bl[253] br[253] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_254 bl[254] br[254] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_255 bl[255] br[255] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_93_0 bl[0] br[0] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_1 bl[1] br[1] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_2 bl[2] br[2] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_3 bl[3] br[3] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_4 bl[4] br[4] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_5 bl[5] br[5] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_6 bl[6] br[6] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_7 bl[7] br[7] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_8 bl[8] br[8] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_9 bl[9] br[9] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_10 bl[10] br[10] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_11 bl[11] br[11] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_12 bl[12] br[12] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_13 bl[13] br[13] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_14 bl[14] br[14] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_15 bl[15] br[15] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_16 bl[16] br[16] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_17 bl[17] br[17] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_18 bl[18] br[18] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_19 bl[19] br[19] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_20 bl[20] br[20] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_21 bl[21] br[21] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_22 bl[22] br[22] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_23 bl[23] br[23] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_24 bl[24] br[24] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_25 bl[25] br[25] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_26 bl[26] br[26] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_27 bl[27] br[27] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_28 bl[28] br[28] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_29 bl[29] br[29] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_30 bl[30] br[30] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_31 bl[31] br[31] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_32 bl[32] br[32] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_33 bl[33] br[33] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_34 bl[34] br[34] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_35 bl[35] br[35] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_36 bl[36] br[36] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_37 bl[37] br[37] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_38 bl[38] br[38] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_39 bl[39] br[39] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_40 bl[40] br[40] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_41 bl[41] br[41] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_42 bl[42] br[42] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_43 bl[43] br[43] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_44 bl[44] br[44] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_45 bl[45] br[45] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_46 bl[46] br[46] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_47 bl[47] br[47] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_48 bl[48] br[48] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_49 bl[49] br[49] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_50 bl[50] br[50] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_51 bl[51] br[51] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_52 bl[52] br[52] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_53 bl[53] br[53] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_54 bl[54] br[54] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_55 bl[55] br[55] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_56 bl[56] br[56] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_57 bl[57] br[57] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_58 bl[58] br[58] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_59 bl[59] br[59] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_60 bl[60] br[60] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_61 bl[61] br[61] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_62 bl[62] br[62] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_63 bl[63] br[63] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_64 bl[64] br[64] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_65 bl[65] br[65] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_66 bl[66] br[66] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_67 bl[67] br[67] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_68 bl[68] br[68] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_69 bl[69] br[69] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_70 bl[70] br[70] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_71 bl[71] br[71] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_72 bl[72] br[72] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_73 bl[73] br[73] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_74 bl[74] br[74] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_75 bl[75] br[75] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_76 bl[76] br[76] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_77 bl[77] br[77] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_78 bl[78] br[78] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_79 bl[79] br[79] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_80 bl[80] br[80] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_81 bl[81] br[81] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_82 bl[82] br[82] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_83 bl[83] br[83] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_84 bl[84] br[84] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_85 bl[85] br[85] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_86 bl[86] br[86] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_87 bl[87] br[87] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_88 bl[88] br[88] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_89 bl[89] br[89] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_90 bl[90] br[90] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_91 bl[91] br[91] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_92 bl[92] br[92] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_93 bl[93] br[93] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_94 bl[94] br[94] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_95 bl[95] br[95] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_96 bl[96] br[96] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_97 bl[97] br[97] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_98 bl[98] br[98] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_99 bl[99] br[99] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_100 bl[100] br[100] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_101 bl[101] br[101] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_102 bl[102] br[102] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_103 bl[103] br[103] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_104 bl[104] br[104] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_105 bl[105] br[105] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_106 bl[106] br[106] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_107 bl[107] br[107] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_108 bl[108] br[108] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_109 bl[109] br[109] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_110 bl[110] br[110] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_111 bl[111] br[111] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_112 bl[112] br[112] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_113 bl[113] br[113] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_114 bl[114] br[114] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_115 bl[115] br[115] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_116 bl[116] br[116] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_117 bl[117] br[117] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_118 bl[118] br[118] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_119 bl[119] br[119] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_120 bl[120] br[120] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_121 bl[121] br[121] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_122 bl[122] br[122] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_123 bl[123] br[123] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_124 bl[124] br[124] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_125 bl[125] br[125] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_126 bl[126] br[126] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_127 bl[127] br[127] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_128 bl[128] br[128] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_129 bl[129] br[129] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_130 bl[130] br[130] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_131 bl[131] br[131] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_132 bl[132] br[132] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_133 bl[133] br[133] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_134 bl[134] br[134] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_135 bl[135] br[135] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_136 bl[136] br[136] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_137 bl[137] br[137] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_138 bl[138] br[138] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_139 bl[139] br[139] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_140 bl[140] br[140] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_141 bl[141] br[141] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_142 bl[142] br[142] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_143 bl[143] br[143] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_144 bl[144] br[144] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_145 bl[145] br[145] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_146 bl[146] br[146] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_147 bl[147] br[147] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_148 bl[148] br[148] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_149 bl[149] br[149] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_150 bl[150] br[150] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_151 bl[151] br[151] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_152 bl[152] br[152] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_153 bl[153] br[153] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_154 bl[154] br[154] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_155 bl[155] br[155] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_156 bl[156] br[156] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_157 bl[157] br[157] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_158 bl[158] br[158] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_159 bl[159] br[159] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_160 bl[160] br[160] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_161 bl[161] br[161] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_162 bl[162] br[162] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_163 bl[163] br[163] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_164 bl[164] br[164] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_165 bl[165] br[165] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_166 bl[166] br[166] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_167 bl[167] br[167] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_168 bl[168] br[168] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_169 bl[169] br[169] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_170 bl[170] br[170] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_171 bl[171] br[171] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_172 bl[172] br[172] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_173 bl[173] br[173] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_174 bl[174] br[174] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_175 bl[175] br[175] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_176 bl[176] br[176] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_177 bl[177] br[177] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_178 bl[178] br[178] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_179 bl[179] br[179] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_180 bl[180] br[180] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_181 bl[181] br[181] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_182 bl[182] br[182] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_183 bl[183] br[183] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_184 bl[184] br[184] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_185 bl[185] br[185] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_186 bl[186] br[186] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_187 bl[187] br[187] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_188 bl[188] br[188] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_189 bl[189] br[189] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_190 bl[190] br[190] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_191 bl[191] br[191] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_192 bl[192] br[192] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_193 bl[193] br[193] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_194 bl[194] br[194] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_195 bl[195] br[195] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_196 bl[196] br[196] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_197 bl[197] br[197] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_198 bl[198] br[198] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_199 bl[199] br[199] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_200 bl[200] br[200] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_201 bl[201] br[201] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_202 bl[202] br[202] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_203 bl[203] br[203] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_204 bl[204] br[204] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_205 bl[205] br[205] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_206 bl[206] br[206] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_207 bl[207] br[207] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_208 bl[208] br[208] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_209 bl[209] br[209] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_210 bl[210] br[210] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_211 bl[211] br[211] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_212 bl[212] br[212] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_213 bl[213] br[213] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_214 bl[214] br[214] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_215 bl[215] br[215] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_216 bl[216] br[216] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_217 bl[217] br[217] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_218 bl[218] br[218] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_219 bl[219] br[219] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_220 bl[220] br[220] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_221 bl[221] br[221] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_222 bl[222] br[222] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_223 bl[223] br[223] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_224 bl[224] br[224] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_225 bl[225] br[225] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_226 bl[226] br[226] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_227 bl[227] br[227] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_228 bl[228] br[228] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_229 bl[229] br[229] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_230 bl[230] br[230] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_231 bl[231] br[231] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_232 bl[232] br[232] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_233 bl[233] br[233] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_234 bl[234] br[234] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_235 bl[235] br[235] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_236 bl[236] br[236] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_237 bl[237] br[237] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_238 bl[238] br[238] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_239 bl[239] br[239] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_240 bl[240] br[240] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_241 bl[241] br[241] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_242 bl[242] br[242] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_243 bl[243] br[243] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_244 bl[244] br[244] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_245 bl[245] br[245] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_246 bl[246] br[246] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_247 bl[247] br[247] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_248 bl[248] br[248] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_249 bl[249] br[249] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_250 bl[250] br[250] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_251 bl[251] br[251] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_252 bl[252] br[252] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_253 bl[253] br[253] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_254 bl[254] br[254] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_255 bl[255] br[255] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_94_0 bl[0] br[0] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_1 bl[1] br[1] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_2 bl[2] br[2] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_3 bl[3] br[3] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_4 bl[4] br[4] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_5 bl[5] br[5] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_6 bl[6] br[6] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_7 bl[7] br[7] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_8 bl[8] br[8] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_9 bl[9] br[9] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_10 bl[10] br[10] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_11 bl[11] br[11] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_12 bl[12] br[12] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_13 bl[13] br[13] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_14 bl[14] br[14] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_15 bl[15] br[15] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_16 bl[16] br[16] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_17 bl[17] br[17] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_18 bl[18] br[18] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_19 bl[19] br[19] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_20 bl[20] br[20] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_21 bl[21] br[21] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_22 bl[22] br[22] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_23 bl[23] br[23] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_24 bl[24] br[24] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_25 bl[25] br[25] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_26 bl[26] br[26] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_27 bl[27] br[27] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_28 bl[28] br[28] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_29 bl[29] br[29] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_30 bl[30] br[30] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_31 bl[31] br[31] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_32 bl[32] br[32] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_33 bl[33] br[33] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_34 bl[34] br[34] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_35 bl[35] br[35] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_36 bl[36] br[36] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_37 bl[37] br[37] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_38 bl[38] br[38] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_39 bl[39] br[39] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_40 bl[40] br[40] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_41 bl[41] br[41] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_42 bl[42] br[42] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_43 bl[43] br[43] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_44 bl[44] br[44] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_45 bl[45] br[45] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_46 bl[46] br[46] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_47 bl[47] br[47] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_48 bl[48] br[48] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_49 bl[49] br[49] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_50 bl[50] br[50] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_51 bl[51] br[51] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_52 bl[52] br[52] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_53 bl[53] br[53] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_54 bl[54] br[54] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_55 bl[55] br[55] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_56 bl[56] br[56] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_57 bl[57] br[57] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_58 bl[58] br[58] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_59 bl[59] br[59] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_60 bl[60] br[60] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_61 bl[61] br[61] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_62 bl[62] br[62] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_63 bl[63] br[63] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_64 bl[64] br[64] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_65 bl[65] br[65] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_66 bl[66] br[66] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_67 bl[67] br[67] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_68 bl[68] br[68] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_69 bl[69] br[69] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_70 bl[70] br[70] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_71 bl[71] br[71] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_72 bl[72] br[72] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_73 bl[73] br[73] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_74 bl[74] br[74] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_75 bl[75] br[75] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_76 bl[76] br[76] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_77 bl[77] br[77] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_78 bl[78] br[78] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_79 bl[79] br[79] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_80 bl[80] br[80] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_81 bl[81] br[81] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_82 bl[82] br[82] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_83 bl[83] br[83] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_84 bl[84] br[84] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_85 bl[85] br[85] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_86 bl[86] br[86] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_87 bl[87] br[87] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_88 bl[88] br[88] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_89 bl[89] br[89] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_90 bl[90] br[90] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_91 bl[91] br[91] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_92 bl[92] br[92] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_93 bl[93] br[93] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_94 bl[94] br[94] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_95 bl[95] br[95] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_96 bl[96] br[96] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_97 bl[97] br[97] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_98 bl[98] br[98] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_99 bl[99] br[99] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_100 bl[100] br[100] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_101 bl[101] br[101] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_102 bl[102] br[102] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_103 bl[103] br[103] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_104 bl[104] br[104] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_105 bl[105] br[105] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_106 bl[106] br[106] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_107 bl[107] br[107] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_108 bl[108] br[108] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_109 bl[109] br[109] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_110 bl[110] br[110] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_111 bl[111] br[111] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_112 bl[112] br[112] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_113 bl[113] br[113] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_114 bl[114] br[114] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_115 bl[115] br[115] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_116 bl[116] br[116] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_117 bl[117] br[117] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_118 bl[118] br[118] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_119 bl[119] br[119] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_120 bl[120] br[120] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_121 bl[121] br[121] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_122 bl[122] br[122] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_123 bl[123] br[123] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_124 bl[124] br[124] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_125 bl[125] br[125] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_126 bl[126] br[126] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_127 bl[127] br[127] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_128 bl[128] br[128] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_129 bl[129] br[129] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_130 bl[130] br[130] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_131 bl[131] br[131] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_132 bl[132] br[132] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_133 bl[133] br[133] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_134 bl[134] br[134] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_135 bl[135] br[135] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_136 bl[136] br[136] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_137 bl[137] br[137] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_138 bl[138] br[138] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_139 bl[139] br[139] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_140 bl[140] br[140] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_141 bl[141] br[141] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_142 bl[142] br[142] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_143 bl[143] br[143] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_144 bl[144] br[144] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_145 bl[145] br[145] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_146 bl[146] br[146] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_147 bl[147] br[147] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_148 bl[148] br[148] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_149 bl[149] br[149] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_150 bl[150] br[150] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_151 bl[151] br[151] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_152 bl[152] br[152] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_153 bl[153] br[153] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_154 bl[154] br[154] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_155 bl[155] br[155] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_156 bl[156] br[156] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_157 bl[157] br[157] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_158 bl[158] br[158] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_159 bl[159] br[159] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_160 bl[160] br[160] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_161 bl[161] br[161] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_162 bl[162] br[162] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_163 bl[163] br[163] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_164 bl[164] br[164] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_165 bl[165] br[165] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_166 bl[166] br[166] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_167 bl[167] br[167] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_168 bl[168] br[168] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_169 bl[169] br[169] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_170 bl[170] br[170] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_171 bl[171] br[171] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_172 bl[172] br[172] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_173 bl[173] br[173] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_174 bl[174] br[174] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_175 bl[175] br[175] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_176 bl[176] br[176] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_177 bl[177] br[177] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_178 bl[178] br[178] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_179 bl[179] br[179] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_180 bl[180] br[180] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_181 bl[181] br[181] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_182 bl[182] br[182] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_183 bl[183] br[183] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_184 bl[184] br[184] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_185 bl[185] br[185] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_186 bl[186] br[186] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_187 bl[187] br[187] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_188 bl[188] br[188] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_189 bl[189] br[189] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_190 bl[190] br[190] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_191 bl[191] br[191] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_192 bl[192] br[192] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_193 bl[193] br[193] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_194 bl[194] br[194] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_195 bl[195] br[195] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_196 bl[196] br[196] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_197 bl[197] br[197] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_198 bl[198] br[198] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_199 bl[199] br[199] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_200 bl[200] br[200] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_201 bl[201] br[201] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_202 bl[202] br[202] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_203 bl[203] br[203] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_204 bl[204] br[204] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_205 bl[205] br[205] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_206 bl[206] br[206] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_207 bl[207] br[207] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_208 bl[208] br[208] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_209 bl[209] br[209] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_210 bl[210] br[210] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_211 bl[211] br[211] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_212 bl[212] br[212] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_213 bl[213] br[213] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_214 bl[214] br[214] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_215 bl[215] br[215] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_216 bl[216] br[216] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_217 bl[217] br[217] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_218 bl[218] br[218] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_219 bl[219] br[219] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_220 bl[220] br[220] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_221 bl[221] br[221] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_222 bl[222] br[222] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_223 bl[223] br[223] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_224 bl[224] br[224] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_225 bl[225] br[225] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_226 bl[226] br[226] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_227 bl[227] br[227] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_228 bl[228] br[228] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_229 bl[229] br[229] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_230 bl[230] br[230] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_231 bl[231] br[231] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_232 bl[232] br[232] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_233 bl[233] br[233] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_234 bl[234] br[234] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_235 bl[235] br[235] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_236 bl[236] br[236] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_237 bl[237] br[237] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_238 bl[238] br[238] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_239 bl[239] br[239] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_240 bl[240] br[240] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_241 bl[241] br[241] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_242 bl[242] br[242] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_243 bl[243] br[243] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_244 bl[244] br[244] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_245 bl[245] br[245] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_246 bl[246] br[246] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_247 bl[247] br[247] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_248 bl[248] br[248] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_249 bl[249] br[249] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_250 bl[250] br[250] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_251 bl[251] br[251] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_252 bl[252] br[252] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_253 bl[253] br[253] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_254 bl[254] br[254] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_255 bl[255] br[255] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_95_0 bl[0] br[0] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_1 bl[1] br[1] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_2 bl[2] br[2] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_3 bl[3] br[3] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_4 bl[4] br[4] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_5 bl[5] br[5] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_6 bl[6] br[6] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_7 bl[7] br[7] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_8 bl[8] br[8] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_9 bl[9] br[9] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_10 bl[10] br[10] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_11 bl[11] br[11] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_12 bl[12] br[12] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_13 bl[13] br[13] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_14 bl[14] br[14] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_15 bl[15] br[15] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_16 bl[16] br[16] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_17 bl[17] br[17] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_18 bl[18] br[18] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_19 bl[19] br[19] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_20 bl[20] br[20] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_21 bl[21] br[21] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_22 bl[22] br[22] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_23 bl[23] br[23] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_24 bl[24] br[24] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_25 bl[25] br[25] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_26 bl[26] br[26] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_27 bl[27] br[27] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_28 bl[28] br[28] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_29 bl[29] br[29] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_30 bl[30] br[30] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_31 bl[31] br[31] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_32 bl[32] br[32] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_33 bl[33] br[33] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_34 bl[34] br[34] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_35 bl[35] br[35] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_36 bl[36] br[36] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_37 bl[37] br[37] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_38 bl[38] br[38] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_39 bl[39] br[39] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_40 bl[40] br[40] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_41 bl[41] br[41] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_42 bl[42] br[42] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_43 bl[43] br[43] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_44 bl[44] br[44] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_45 bl[45] br[45] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_46 bl[46] br[46] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_47 bl[47] br[47] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_48 bl[48] br[48] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_49 bl[49] br[49] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_50 bl[50] br[50] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_51 bl[51] br[51] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_52 bl[52] br[52] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_53 bl[53] br[53] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_54 bl[54] br[54] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_55 bl[55] br[55] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_56 bl[56] br[56] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_57 bl[57] br[57] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_58 bl[58] br[58] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_59 bl[59] br[59] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_60 bl[60] br[60] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_61 bl[61] br[61] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_62 bl[62] br[62] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_63 bl[63] br[63] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_64 bl[64] br[64] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_65 bl[65] br[65] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_66 bl[66] br[66] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_67 bl[67] br[67] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_68 bl[68] br[68] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_69 bl[69] br[69] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_70 bl[70] br[70] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_71 bl[71] br[71] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_72 bl[72] br[72] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_73 bl[73] br[73] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_74 bl[74] br[74] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_75 bl[75] br[75] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_76 bl[76] br[76] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_77 bl[77] br[77] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_78 bl[78] br[78] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_79 bl[79] br[79] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_80 bl[80] br[80] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_81 bl[81] br[81] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_82 bl[82] br[82] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_83 bl[83] br[83] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_84 bl[84] br[84] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_85 bl[85] br[85] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_86 bl[86] br[86] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_87 bl[87] br[87] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_88 bl[88] br[88] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_89 bl[89] br[89] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_90 bl[90] br[90] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_91 bl[91] br[91] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_92 bl[92] br[92] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_93 bl[93] br[93] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_94 bl[94] br[94] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_95 bl[95] br[95] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_96 bl[96] br[96] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_97 bl[97] br[97] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_98 bl[98] br[98] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_99 bl[99] br[99] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_100 bl[100] br[100] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_101 bl[101] br[101] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_102 bl[102] br[102] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_103 bl[103] br[103] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_104 bl[104] br[104] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_105 bl[105] br[105] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_106 bl[106] br[106] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_107 bl[107] br[107] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_108 bl[108] br[108] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_109 bl[109] br[109] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_110 bl[110] br[110] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_111 bl[111] br[111] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_112 bl[112] br[112] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_113 bl[113] br[113] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_114 bl[114] br[114] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_115 bl[115] br[115] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_116 bl[116] br[116] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_117 bl[117] br[117] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_118 bl[118] br[118] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_119 bl[119] br[119] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_120 bl[120] br[120] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_121 bl[121] br[121] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_122 bl[122] br[122] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_123 bl[123] br[123] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_124 bl[124] br[124] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_125 bl[125] br[125] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_126 bl[126] br[126] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_127 bl[127] br[127] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_128 bl[128] br[128] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_129 bl[129] br[129] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_130 bl[130] br[130] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_131 bl[131] br[131] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_132 bl[132] br[132] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_133 bl[133] br[133] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_134 bl[134] br[134] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_135 bl[135] br[135] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_136 bl[136] br[136] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_137 bl[137] br[137] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_138 bl[138] br[138] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_139 bl[139] br[139] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_140 bl[140] br[140] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_141 bl[141] br[141] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_142 bl[142] br[142] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_143 bl[143] br[143] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_144 bl[144] br[144] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_145 bl[145] br[145] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_146 bl[146] br[146] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_147 bl[147] br[147] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_148 bl[148] br[148] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_149 bl[149] br[149] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_150 bl[150] br[150] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_151 bl[151] br[151] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_152 bl[152] br[152] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_153 bl[153] br[153] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_154 bl[154] br[154] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_155 bl[155] br[155] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_156 bl[156] br[156] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_157 bl[157] br[157] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_158 bl[158] br[158] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_159 bl[159] br[159] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_160 bl[160] br[160] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_161 bl[161] br[161] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_162 bl[162] br[162] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_163 bl[163] br[163] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_164 bl[164] br[164] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_165 bl[165] br[165] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_166 bl[166] br[166] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_167 bl[167] br[167] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_168 bl[168] br[168] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_169 bl[169] br[169] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_170 bl[170] br[170] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_171 bl[171] br[171] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_172 bl[172] br[172] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_173 bl[173] br[173] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_174 bl[174] br[174] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_175 bl[175] br[175] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_176 bl[176] br[176] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_177 bl[177] br[177] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_178 bl[178] br[178] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_179 bl[179] br[179] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_180 bl[180] br[180] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_181 bl[181] br[181] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_182 bl[182] br[182] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_183 bl[183] br[183] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_184 bl[184] br[184] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_185 bl[185] br[185] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_186 bl[186] br[186] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_187 bl[187] br[187] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_188 bl[188] br[188] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_189 bl[189] br[189] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_190 bl[190] br[190] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_191 bl[191] br[191] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_192 bl[192] br[192] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_193 bl[193] br[193] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_194 bl[194] br[194] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_195 bl[195] br[195] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_196 bl[196] br[196] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_197 bl[197] br[197] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_198 bl[198] br[198] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_199 bl[199] br[199] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_200 bl[200] br[200] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_201 bl[201] br[201] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_202 bl[202] br[202] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_203 bl[203] br[203] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_204 bl[204] br[204] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_205 bl[205] br[205] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_206 bl[206] br[206] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_207 bl[207] br[207] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_208 bl[208] br[208] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_209 bl[209] br[209] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_210 bl[210] br[210] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_211 bl[211] br[211] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_212 bl[212] br[212] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_213 bl[213] br[213] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_214 bl[214] br[214] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_215 bl[215] br[215] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_216 bl[216] br[216] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_217 bl[217] br[217] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_218 bl[218] br[218] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_219 bl[219] br[219] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_220 bl[220] br[220] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_221 bl[221] br[221] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_222 bl[222] br[222] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_223 bl[223] br[223] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_224 bl[224] br[224] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_225 bl[225] br[225] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_226 bl[226] br[226] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_227 bl[227] br[227] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_228 bl[228] br[228] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_229 bl[229] br[229] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_230 bl[230] br[230] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_231 bl[231] br[231] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_232 bl[232] br[232] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_233 bl[233] br[233] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_234 bl[234] br[234] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_235 bl[235] br[235] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_236 bl[236] br[236] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_237 bl[237] br[237] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_238 bl[238] br[238] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_239 bl[239] br[239] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_240 bl[240] br[240] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_241 bl[241] br[241] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_242 bl[242] br[242] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_243 bl[243] br[243] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_244 bl[244] br[244] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_245 bl[245] br[245] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_246 bl[246] br[246] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_247 bl[247] br[247] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_248 bl[248] br[248] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_249 bl[249] br[249] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_250 bl[250] br[250] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_251 bl[251] br[251] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_252 bl[252] br[252] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_253 bl[253] br[253] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_254 bl[254] br[254] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_255 bl[255] br[255] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_96_0 bl[0] br[0] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_1 bl[1] br[1] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_2 bl[2] br[2] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_3 bl[3] br[3] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_4 bl[4] br[4] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_5 bl[5] br[5] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_6 bl[6] br[6] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_7 bl[7] br[7] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_8 bl[8] br[8] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_9 bl[9] br[9] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_10 bl[10] br[10] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_11 bl[11] br[11] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_12 bl[12] br[12] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_13 bl[13] br[13] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_14 bl[14] br[14] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_15 bl[15] br[15] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_16 bl[16] br[16] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_17 bl[17] br[17] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_18 bl[18] br[18] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_19 bl[19] br[19] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_20 bl[20] br[20] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_21 bl[21] br[21] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_22 bl[22] br[22] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_23 bl[23] br[23] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_24 bl[24] br[24] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_25 bl[25] br[25] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_26 bl[26] br[26] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_27 bl[27] br[27] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_28 bl[28] br[28] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_29 bl[29] br[29] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_30 bl[30] br[30] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_31 bl[31] br[31] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_32 bl[32] br[32] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_33 bl[33] br[33] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_34 bl[34] br[34] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_35 bl[35] br[35] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_36 bl[36] br[36] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_37 bl[37] br[37] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_38 bl[38] br[38] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_39 bl[39] br[39] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_40 bl[40] br[40] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_41 bl[41] br[41] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_42 bl[42] br[42] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_43 bl[43] br[43] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_44 bl[44] br[44] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_45 bl[45] br[45] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_46 bl[46] br[46] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_47 bl[47] br[47] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_48 bl[48] br[48] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_49 bl[49] br[49] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_50 bl[50] br[50] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_51 bl[51] br[51] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_52 bl[52] br[52] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_53 bl[53] br[53] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_54 bl[54] br[54] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_55 bl[55] br[55] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_56 bl[56] br[56] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_57 bl[57] br[57] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_58 bl[58] br[58] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_59 bl[59] br[59] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_60 bl[60] br[60] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_61 bl[61] br[61] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_62 bl[62] br[62] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_63 bl[63] br[63] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_64 bl[64] br[64] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_65 bl[65] br[65] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_66 bl[66] br[66] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_67 bl[67] br[67] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_68 bl[68] br[68] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_69 bl[69] br[69] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_70 bl[70] br[70] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_71 bl[71] br[71] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_72 bl[72] br[72] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_73 bl[73] br[73] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_74 bl[74] br[74] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_75 bl[75] br[75] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_76 bl[76] br[76] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_77 bl[77] br[77] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_78 bl[78] br[78] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_79 bl[79] br[79] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_80 bl[80] br[80] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_81 bl[81] br[81] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_82 bl[82] br[82] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_83 bl[83] br[83] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_84 bl[84] br[84] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_85 bl[85] br[85] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_86 bl[86] br[86] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_87 bl[87] br[87] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_88 bl[88] br[88] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_89 bl[89] br[89] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_90 bl[90] br[90] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_91 bl[91] br[91] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_92 bl[92] br[92] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_93 bl[93] br[93] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_94 bl[94] br[94] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_95 bl[95] br[95] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_96 bl[96] br[96] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_97 bl[97] br[97] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_98 bl[98] br[98] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_99 bl[99] br[99] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_100 bl[100] br[100] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_101 bl[101] br[101] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_102 bl[102] br[102] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_103 bl[103] br[103] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_104 bl[104] br[104] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_105 bl[105] br[105] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_106 bl[106] br[106] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_107 bl[107] br[107] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_108 bl[108] br[108] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_109 bl[109] br[109] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_110 bl[110] br[110] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_111 bl[111] br[111] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_112 bl[112] br[112] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_113 bl[113] br[113] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_114 bl[114] br[114] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_115 bl[115] br[115] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_116 bl[116] br[116] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_117 bl[117] br[117] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_118 bl[118] br[118] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_119 bl[119] br[119] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_120 bl[120] br[120] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_121 bl[121] br[121] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_122 bl[122] br[122] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_123 bl[123] br[123] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_124 bl[124] br[124] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_125 bl[125] br[125] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_126 bl[126] br[126] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_127 bl[127] br[127] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_128 bl[128] br[128] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_129 bl[129] br[129] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_130 bl[130] br[130] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_131 bl[131] br[131] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_132 bl[132] br[132] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_133 bl[133] br[133] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_134 bl[134] br[134] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_135 bl[135] br[135] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_136 bl[136] br[136] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_137 bl[137] br[137] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_138 bl[138] br[138] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_139 bl[139] br[139] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_140 bl[140] br[140] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_141 bl[141] br[141] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_142 bl[142] br[142] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_143 bl[143] br[143] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_144 bl[144] br[144] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_145 bl[145] br[145] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_146 bl[146] br[146] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_147 bl[147] br[147] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_148 bl[148] br[148] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_149 bl[149] br[149] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_150 bl[150] br[150] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_151 bl[151] br[151] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_152 bl[152] br[152] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_153 bl[153] br[153] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_154 bl[154] br[154] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_155 bl[155] br[155] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_156 bl[156] br[156] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_157 bl[157] br[157] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_158 bl[158] br[158] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_159 bl[159] br[159] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_160 bl[160] br[160] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_161 bl[161] br[161] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_162 bl[162] br[162] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_163 bl[163] br[163] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_164 bl[164] br[164] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_165 bl[165] br[165] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_166 bl[166] br[166] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_167 bl[167] br[167] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_168 bl[168] br[168] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_169 bl[169] br[169] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_170 bl[170] br[170] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_171 bl[171] br[171] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_172 bl[172] br[172] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_173 bl[173] br[173] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_174 bl[174] br[174] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_175 bl[175] br[175] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_176 bl[176] br[176] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_177 bl[177] br[177] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_178 bl[178] br[178] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_179 bl[179] br[179] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_180 bl[180] br[180] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_181 bl[181] br[181] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_182 bl[182] br[182] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_183 bl[183] br[183] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_184 bl[184] br[184] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_185 bl[185] br[185] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_186 bl[186] br[186] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_187 bl[187] br[187] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_188 bl[188] br[188] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_189 bl[189] br[189] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_190 bl[190] br[190] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_191 bl[191] br[191] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_192 bl[192] br[192] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_193 bl[193] br[193] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_194 bl[194] br[194] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_195 bl[195] br[195] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_196 bl[196] br[196] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_197 bl[197] br[197] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_198 bl[198] br[198] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_199 bl[199] br[199] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_200 bl[200] br[200] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_201 bl[201] br[201] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_202 bl[202] br[202] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_203 bl[203] br[203] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_204 bl[204] br[204] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_205 bl[205] br[205] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_206 bl[206] br[206] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_207 bl[207] br[207] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_208 bl[208] br[208] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_209 bl[209] br[209] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_210 bl[210] br[210] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_211 bl[211] br[211] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_212 bl[212] br[212] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_213 bl[213] br[213] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_214 bl[214] br[214] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_215 bl[215] br[215] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_216 bl[216] br[216] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_217 bl[217] br[217] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_218 bl[218] br[218] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_219 bl[219] br[219] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_220 bl[220] br[220] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_221 bl[221] br[221] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_222 bl[222] br[222] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_223 bl[223] br[223] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_224 bl[224] br[224] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_225 bl[225] br[225] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_226 bl[226] br[226] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_227 bl[227] br[227] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_228 bl[228] br[228] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_229 bl[229] br[229] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_230 bl[230] br[230] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_231 bl[231] br[231] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_232 bl[232] br[232] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_233 bl[233] br[233] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_234 bl[234] br[234] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_235 bl[235] br[235] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_236 bl[236] br[236] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_237 bl[237] br[237] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_238 bl[238] br[238] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_239 bl[239] br[239] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_240 bl[240] br[240] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_241 bl[241] br[241] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_242 bl[242] br[242] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_243 bl[243] br[243] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_244 bl[244] br[244] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_245 bl[245] br[245] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_246 bl[246] br[246] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_247 bl[247] br[247] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_248 bl[248] br[248] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_249 bl[249] br[249] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_250 bl[250] br[250] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_251 bl[251] br[251] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_252 bl[252] br[252] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_253 bl[253] br[253] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_254 bl[254] br[254] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_255 bl[255] br[255] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_97_0 bl[0] br[0] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_1 bl[1] br[1] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_2 bl[2] br[2] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_3 bl[3] br[3] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_4 bl[4] br[4] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_5 bl[5] br[5] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_6 bl[6] br[6] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_7 bl[7] br[7] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_8 bl[8] br[8] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_9 bl[9] br[9] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_10 bl[10] br[10] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_11 bl[11] br[11] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_12 bl[12] br[12] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_13 bl[13] br[13] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_14 bl[14] br[14] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_15 bl[15] br[15] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_16 bl[16] br[16] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_17 bl[17] br[17] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_18 bl[18] br[18] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_19 bl[19] br[19] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_20 bl[20] br[20] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_21 bl[21] br[21] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_22 bl[22] br[22] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_23 bl[23] br[23] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_24 bl[24] br[24] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_25 bl[25] br[25] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_26 bl[26] br[26] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_27 bl[27] br[27] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_28 bl[28] br[28] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_29 bl[29] br[29] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_30 bl[30] br[30] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_31 bl[31] br[31] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_32 bl[32] br[32] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_33 bl[33] br[33] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_34 bl[34] br[34] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_35 bl[35] br[35] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_36 bl[36] br[36] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_37 bl[37] br[37] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_38 bl[38] br[38] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_39 bl[39] br[39] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_40 bl[40] br[40] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_41 bl[41] br[41] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_42 bl[42] br[42] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_43 bl[43] br[43] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_44 bl[44] br[44] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_45 bl[45] br[45] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_46 bl[46] br[46] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_47 bl[47] br[47] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_48 bl[48] br[48] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_49 bl[49] br[49] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_50 bl[50] br[50] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_51 bl[51] br[51] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_52 bl[52] br[52] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_53 bl[53] br[53] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_54 bl[54] br[54] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_55 bl[55] br[55] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_56 bl[56] br[56] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_57 bl[57] br[57] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_58 bl[58] br[58] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_59 bl[59] br[59] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_60 bl[60] br[60] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_61 bl[61] br[61] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_62 bl[62] br[62] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_63 bl[63] br[63] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_64 bl[64] br[64] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_65 bl[65] br[65] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_66 bl[66] br[66] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_67 bl[67] br[67] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_68 bl[68] br[68] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_69 bl[69] br[69] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_70 bl[70] br[70] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_71 bl[71] br[71] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_72 bl[72] br[72] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_73 bl[73] br[73] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_74 bl[74] br[74] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_75 bl[75] br[75] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_76 bl[76] br[76] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_77 bl[77] br[77] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_78 bl[78] br[78] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_79 bl[79] br[79] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_80 bl[80] br[80] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_81 bl[81] br[81] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_82 bl[82] br[82] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_83 bl[83] br[83] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_84 bl[84] br[84] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_85 bl[85] br[85] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_86 bl[86] br[86] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_87 bl[87] br[87] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_88 bl[88] br[88] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_89 bl[89] br[89] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_90 bl[90] br[90] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_91 bl[91] br[91] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_92 bl[92] br[92] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_93 bl[93] br[93] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_94 bl[94] br[94] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_95 bl[95] br[95] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_96 bl[96] br[96] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_97 bl[97] br[97] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_98 bl[98] br[98] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_99 bl[99] br[99] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_100 bl[100] br[100] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_101 bl[101] br[101] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_102 bl[102] br[102] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_103 bl[103] br[103] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_104 bl[104] br[104] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_105 bl[105] br[105] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_106 bl[106] br[106] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_107 bl[107] br[107] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_108 bl[108] br[108] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_109 bl[109] br[109] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_110 bl[110] br[110] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_111 bl[111] br[111] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_112 bl[112] br[112] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_113 bl[113] br[113] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_114 bl[114] br[114] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_115 bl[115] br[115] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_116 bl[116] br[116] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_117 bl[117] br[117] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_118 bl[118] br[118] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_119 bl[119] br[119] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_120 bl[120] br[120] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_121 bl[121] br[121] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_122 bl[122] br[122] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_123 bl[123] br[123] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_124 bl[124] br[124] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_125 bl[125] br[125] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_126 bl[126] br[126] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_127 bl[127] br[127] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_128 bl[128] br[128] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_129 bl[129] br[129] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_130 bl[130] br[130] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_131 bl[131] br[131] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_132 bl[132] br[132] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_133 bl[133] br[133] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_134 bl[134] br[134] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_135 bl[135] br[135] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_136 bl[136] br[136] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_137 bl[137] br[137] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_138 bl[138] br[138] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_139 bl[139] br[139] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_140 bl[140] br[140] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_141 bl[141] br[141] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_142 bl[142] br[142] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_143 bl[143] br[143] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_144 bl[144] br[144] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_145 bl[145] br[145] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_146 bl[146] br[146] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_147 bl[147] br[147] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_148 bl[148] br[148] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_149 bl[149] br[149] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_150 bl[150] br[150] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_151 bl[151] br[151] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_152 bl[152] br[152] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_153 bl[153] br[153] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_154 bl[154] br[154] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_155 bl[155] br[155] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_156 bl[156] br[156] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_157 bl[157] br[157] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_158 bl[158] br[158] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_159 bl[159] br[159] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_160 bl[160] br[160] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_161 bl[161] br[161] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_162 bl[162] br[162] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_163 bl[163] br[163] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_164 bl[164] br[164] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_165 bl[165] br[165] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_166 bl[166] br[166] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_167 bl[167] br[167] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_168 bl[168] br[168] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_169 bl[169] br[169] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_170 bl[170] br[170] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_171 bl[171] br[171] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_172 bl[172] br[172] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_173 bl[173] br[173] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_174 bl[174] br[174] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_175 bl[175] br[175] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_176 bl[176] br[176] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_177 bl[177] br[177] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_178 bl[178] br[178] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_179 bl[179] br[179] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_180 bl[180] br[180] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_181 bl[181] br[181] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_182 bl[182] br[182] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_183 bl[183] br[183] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_184 bl[184] br[184] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_185 bl[185] br[185] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_186 bl[186] br[186] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_187 bl[187] br[187] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_188 bl[188] br[188] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_189 bl[189] br[189] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_190 bl[190] br[190] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_191 bl[191] br[191] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_192 bl[192] br[192] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_193 bl[193] br[193] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_194 bl[194] br[194] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_195 bl[195] br[195] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_196 bl[196] br[196] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_197 bl[197] br[197] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_198 bl[198] br[198] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_199 bl[199] br[199] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_200 bl[200] br[200] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_201 bl[201] br[201] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_202 bl[202] br[202] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_203 bl[203] br[203] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_204 bl[204] br[204] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_205 bl[205] br[205] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_206 bl[206] br[206] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_207 bl[207] br[207] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_208 bl[208] br[208] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_209 bl[209] br[209] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_210 bl[210] br[210] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_211 bl[211] br[211] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_212 bl[212] br[212] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_213 bl[213] br[213] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_214 bl[214] br[214] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_215 bl[215] br[215] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_216 bl[216] br[216] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_217 bl[217] br[217] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_218 bl[218] br[218] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_219 bl[219] br[219] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_220 bl[220] br[220] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_221 bl[221] br[221] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_222 bl[222] br[222] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_223 bl[223] br[223] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_224 bl[224] br[224] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_225 bl[225] br[225] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_226 bl[226] br[226] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_227 bl[227] br[227] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_228 bl[228] br[228] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_229 bl[229] br[229] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_230 bl[230] br[230] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_231 bl[231] br[231] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_232 bl[232] br[232] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_233 bl[233] br[233] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_234 bl[234] br[234] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_235 bl[235] br[235] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_236 bl[236] br[236] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_237 bl[237] br[237] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_238 bl[238] br[238] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_239 bl[239] br[239] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_240 bl[240] br[240] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_241 bl[241] br[241] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_242 bl[242] br[242] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_243 bl[243] br[243] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_244 bl[244] br[244] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_245 bl[245] br[245] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_246 bl[246] br[246] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_247 bl[247] br[247] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_248 bl[248] br[248] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_249 bl[249] br[249] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_250 bl[250] br[250] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_251 bl[251] br[251] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_252 bl[252] br[252] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_253 bl[253] br[253] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_254 bl[254] br[254] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_255 bl[255] br[255] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_98_0 bl[0] br[0] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_1 bl[1] br[1] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_2 bl[2] br[2] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_3 bl[3] br[3] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_4 bl[4] br[4] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_5 bl[5] br[5] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_6 bl[6] br[6] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_7 bl[7] br[7] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_8 bl[8] br[8] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_9 bl[9] br[9] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_10 bl[10] br[10] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_11 bl[11] br[11] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_12 bl[12] br[12] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_13 bl[13] br[13] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_14 bl[14] br[14] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_15 bl[15] br[15] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_16 bl[16] br[16] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_17 bl[17] br[17] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_18 bl[18] br[18] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_19 bl[19] br[19] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_20 bl[20] br[20] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_21 bl[21] br[21] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_22 bl[22] br[22] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_23 bl[23] br[23] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_24 bl[24] br[24] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_25 bl[25] br[25] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_26 bl[26] br[26] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_27 bl[27] br[27] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_28 bl[28] br[28] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_29 bl[29] br[29] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_30 bl[30] br[30] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_31 bl[31] br[31] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_32 bl[32] br[32] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_33 bl[33] br[33] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_34 bl[34] br[34] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_35 bl[35] br[35] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_36 bl[36] br[36] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_37 bl[37] br[37] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_38 bl[38] br[38] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_39 bl[39] br[39] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_40 bl[40] br[40] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_41 bl[41] br[41] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_42 bl[42] br[42] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_43 bl[43] br[43] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_44 bl[44] br[44] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_45 bl[45] br[45] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_46 bl[46] br[46] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_47 bl[47] br[47] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_48 bl[48] br[48] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_49 bl[49] br[49] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_50 bl[50] br[50] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_51 bl[51] br[51] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_52 bl[52] br[52] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_53 bl[53] br[53] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_54 bl[54] br[54] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_55 bl[55] br[55] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_56 bl[56] br[56] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_57 bl[57] br[57] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_58 bl[58] br[58] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_59 bl[59] br[59] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_60 bl[60] br[60] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_61 bl[61] br[61] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_62 bl[62] br[62] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_63 bl[63] br[63] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_64 bl[64] br[64] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_65 bl[65] br[65] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_66 bl[66] br[66] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_67 bl[67] br[67] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_68 bl[68] br[68] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_69 bl[69] br[69] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_70 bl[70] br[70] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_71 bl[71] br[71] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_72 bl[72] br[72] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_73 bl[73] br[73] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_74 bl[74] br[74] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_75 bl[75] br[75] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_76 bl[76] br[76] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_77 bl[77] br[77] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_78 bl[78] br[78] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_79 bl[79] br[79] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_80 bl[80] br[80] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_81 bl[81] br[81] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_82 bl[82] br[82] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_83 bl[83] br[83] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_84 bl[84] br[84] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_85 bl[85] br[85] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_86 bl[86] br[86] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_87 bl[87] br[87] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_88 bl[88] br[88] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_89 bl[89] br[89] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_90 bl[90] br[90] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_91 bl[91] br[91] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_92 bl[92] br[92] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_93 bl[93] br[93] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_94 bl[94] br[94] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_95 bl[95] br[95] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_96 bl[96] br[96] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_97 bl[97] br[97] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_98 bl[98] br[98] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_99 bl[99] br[99] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_100 bl[100] br[100] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_101 bl[101] br[101] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_102 bl[102] br[102] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_103 bl[103] br[103] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_104 bl[104] br[104] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_105 bl[105] br[105] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_106 bl[106] br[106] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_107 bl[107] br[107] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_108 bl[108] br[108] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_109 bl[109] br[109] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_110 bl[110] br[110] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_111 bl[111] br[111] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_112 bl[112] br[112] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_113 bl[113] br[113] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_114 bl[114] br[114] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_115 bl[115] br[115] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_116 bl[116] br[116] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_117 bl[117] br[117] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_118 bl[118] br[118] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_119 bl[119] br[119] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_120 bl[120] br[120] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_121 bl[121] br[121] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_122 bl[122] br[122] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_123 bl[123] br[123] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_124 bl[124] br[124] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_125 bl[125] br[125] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_126 bl[126] br[126] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_127 bl[127] br[127] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_128 bl[128] br[128] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_129 bl[129] br[129] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_130 bl[130] br[130] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_131 bl[131] br[131] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_132 bl[132] br[132] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_133 bl[133] br[133] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_134 bl[134] br[134] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_135 bl[135] br[135] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_136 bl[136] br[136] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_137 bl[137] br[137] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_138 bl[138] br[138] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_139 bl[139] br[139] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_140 bl[140] br[140] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_141 bl[141] br[141] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_142 bl[142] br[142] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_143 bl[143] br[143] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_144 bl[144] br[144] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_145 bl[145] br[145] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_146 bl[146] br[146] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_147 bl[147] br[147] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_148 bl[148] br[148] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_149 bl[149] br[149] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_150 bl[150] br[150] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_151 bl[151] br[151] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_152 bl[152] br[152] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_153 bl[153] br[153] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_154 bl[154] br[154] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_155 bl[155] br[155] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_156 bl[156] br[156] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_157 bl[157] br[157] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_158 bl[158] br[158] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_159 bl[159] br[159] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_160 bl[160] br[160] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_161 bl[161] br[161] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_162 bl[162] br[162] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_163 bl[163] br[163] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_164 bl[164] br[164] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_165 bl[165] br[165] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_166 bl[166] br[166] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_167 bl[167] br[167] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_168 bl[168] br[168] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_169 bl[169] br[169] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_170 bl[170] br[170] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_171 bl[171] br[171] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_172 bl[172] br[172] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_173 bl[173] br[173] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_174 bl[174] br[174] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_175 bl[175] br[175] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_176 bl[176] br[176] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_177 bl[177] br[177] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_178 bl[178] br[178] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_179 bl[179] br[179] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_180 bl[180] br[180] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_181 bl[181] br[181] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_182 bl[182] br[182] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_183 bl[183] br[183] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_184 bl[184] br[184] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_185 bl[185] br[185] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_186 bl[186] br[186] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_187 bl[187] br[187] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_188 bl[188] br[188] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_189 bl[189] br[189] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_190 bl[190] br[190] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_191 bl[191] br[191] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_192 bl[192] br[192] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_193 bl[193] br[193] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_194 bl[194] br[194] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_195 bl[195] br[195] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_196 bl[196] br[196] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_197 bl[197] br[197] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_198 bl[198] br[198] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_199 bl[199] br[199] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_200 bl[200] br[200] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_201 bl[201] br[201] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_202 bl[202] br[202] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_203 bl[203] br[203] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_204 bl[204] br[204] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_205 bl[205] br[205] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_206 bl[206] br[206] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_207 bl[207] br[207] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_208 bl[208] br[208] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_209 bl[209] br[209] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_210 bl[210] br[210] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_211 bl[211] br[211] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_212 bl[212] br[212] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_213 bl[213] br[213] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_214 bl[214] br[214] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_215 bl[215] br[215] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_216 bl[216] br[216] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_217 bl[217] br[217] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_218 bl[218] br[218] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_219 bl[219] br[219] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_220 bl[220] br[220] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_221 bl[221] br[221] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_222 bl[222] br[222] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_223 bl[223] br[223] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_224 bl[224] br[224] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_225 bl[225] br[225] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_226 bl[226] br[226] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_227 bl[227] br[227] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_228 bl[228] br[228] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_229 bl[229] br[229] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_230 bl[230] br[230] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_231 bl[231] br[231] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_232 bl[232] br[232] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_233 bl[233] br[233] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_234 bl[234] br[234] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_235 bl[235] br[235] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_236 bl[236] br[236] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_237 bl[237] br[237] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_238 bl[238] br[238] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_239 bl[239] br[239] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_240 bl[240] br[240] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_241 bl[241] br[241] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_242 bl[242] br[242] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_243 bl[243] br[243] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_244 bl[244] br[244] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_245 bl[245] br[245] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_246 bl[246] br[246] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_247 bl[247] br[247] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_248 bl[248] br[248] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_249 bl[249] br[249] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_250 bl[250] br[250] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_251 bl[251] br[251] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_252 bl[252] br[252] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_253 bl[253] br[253] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_254 bl[254] br[254] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_255 bl[255] br[255] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_99_0 bl[0] br[0] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_1 bl[1] br[1] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_2 bl[2] br[2] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_3 bl[3] br[3] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_4 bl[4] br[4] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_5 bl[5] br[5] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_6 bl[6] br[6] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_7 bl[7] br[7] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_8 bl[8] br[8] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_9 bl[9] br[9] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_10 bl[10] br[10] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_11 bl[11] br[11] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_12 bl[12] br[12] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_13 bl[13] br[13] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_14 bl[14] br[14] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_15 bl[15] br[15] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_16 bl[16] br[16] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_17 bl[17] br[17] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_18 bl[18] br[18] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_19 bl[19] br[19] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_20 bl[20] br[20] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_21 bl[21] br[21] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_22 bl[22] br[22] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_23 bl[23] br[23] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_24 bl[24] br[24] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_25 bl[25] br[25] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_26 bl[26] br[26] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_27 bl[27] br[27] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_28 bl[28] br[28] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_29 bl[29] br[29] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_30 bl[30] br[30] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_31 bl[31] br[31] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_32 bl[32] br[32] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_33 bl[33] br[33] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_34 bl[34] br[34] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_35 bl[35] br[35] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_36 bl[36] br[36] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_37 bl[37] br[37] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_38 bl[38] br[38] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_39 bl[39] br[39] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_40 bl[40] br[40] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_41 bl[41] br[41] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_42 bl[42] br[42] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_43 bl[43] br[43] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_44 bl[44] br[44] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_45 bl[45] br[45] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_46 bl[46] br[46] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_47 bl[47] br[47] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_48 bl[48] br[48] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_49 bl[49] br[49] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_50 bl[50] br[50] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_51 bl[51] br[51] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_52 bl[52] br[52] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_53 bl[53] br[53] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_54 bl[54] br[54] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_55 bl[55] br[55] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_56 bl[56] br[56] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_57 bl[57] br[57] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_58 bl[58] br[58] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_59 bl[59] br[59] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_60 bl[60] br[60] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_61 bl[61] br[61] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_62 bl[62] br[62] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_63 bl[63] br[63] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_64 bl[64] br[64] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_65 bl[65] br[65] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_66 bl[66] br[66] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_67 bl[67] br[67] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_68 bl[68] br[68] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_69 bl[69] br[69] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_70 bl[70] br[70] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_71 bl[71] br[71] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_72 bl[72] br[72] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_73 bl[73] br[73] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_74 bl[74] br[74] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_75 bl[75] br[75] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_76 bl[76] br[76] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_77 bl[77] br[77] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_78 bl[78] br[78] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_79 bl[79] br[79] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_80 bl[80] br[80] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_81 bl[81] br[81] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_82 bl[82] br[82] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_83 bl[83] br[83] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_84 bl[84] br[84] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_85 bl[85] br[85] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_86 bl[86] br[86] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_87 bl[87] br[87] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_88 bl[88] br[88] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_89 bl[89] br[89] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_90 bl[90] br[90] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_91 bl[91] br[91] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_92 bl[92] br[92] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_93 bl[93] br[93] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_94 bl[94] br[94] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_95 bl[95] br[95] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_96 bl[96] br[96] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_97 bl[97] br[97] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_98 bl[98] br[98] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_99 bl[99] br[99] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_100 bl[100] br[100] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_101 bl[101] br[101] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_102 bl[102] br[102] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_103 bl[103] br[103] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_104 bl[104] br[104] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_105 bl[105] br[105] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_106 bl[106] br[106] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_107 bl[107] br[107] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_108 bl[108] br[108] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_109 bl[109] br[109] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_110 bl[110] br[110] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_111 bl[111] br[111] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_112 bl[112] br[112] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_113 bl[113] br[113] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_114 bl[114] br[114] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_115 bl[115] br[115] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_116 bl[116] br[116] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_117 bl[117] br[117] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_118 bl[118] br[118] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_119 bl[119] br[119] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_120 bl[120] br[120] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_121 bl[121] br[121] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_122 bl[122] br[122] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_123 bl[123] br[123] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_124 bl[124] br[124] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_125 bl[125] br[125] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_126 bl[126] br[126] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_127 bl[127] br[127] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_128 bl[128] br[128] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_129 bl[129] br[129] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_130 bl[130] br[130] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_131 bl[131] br[131] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_132 bl[132] br[132] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_133 bl[133] br[133] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_134 bl[134] br[134] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_135 bl[135] br[135] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_136 bl[136] br[136] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_137 bl[137] br[137] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_138 bl[138] br[138] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_139 bl[139] br[139] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_140 bl[140] br[140] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_141 bl[141] br[141] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_142 bl[142] br[142] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_143 bl[143] br[143] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_144 bl[144] br[144] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_145 bl[145] br[145] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_146 bl[146] br[146] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_147 bl[147] br[147] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_148 bl[148] br[148] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_149 bl[149] br[149] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_150 bl[150] br[150] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_151 bl[151] br[151] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_152 bl[152] br[152] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_153 bl[153] br[153] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_154 bl[154] br[154] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_155 bl[155] br[155] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_156 bl[156] br[156] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_157 bl[157] br[157] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_158 bl[158] br[158] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_159 bl[159] br[159] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_160 bl[160] br[160] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_161 bl[161] br[161] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_162 bl[162] br[162] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_163 bl[163] br[163] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_164 bl[164] br[164] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_165 bl[165] br[165] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_166 bl[166] br[166] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_167 bl[167] br[167] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_168 bl[168] br[168] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_169 bl[169] br[169] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_170 bl[170] br[170] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_171 bl[171] br[171] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_172 bl[172] br[172] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_173 bl[173] br[173] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_174 bl[174] br[174] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_175 bl[175] br[175] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_176 bl[176] br[176] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_177 bl[177] br[177] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_178 bl[178] br[178] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_179 bl[179] br[179] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_180 bl[180] br[180] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_181 bl[181] br[181] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_182 bl[182] br[182] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_183 bl[183] br[183] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_184 bl[184] br[184] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_185 bl[185] br[185] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_186 bl[186] br[186] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_187 bl[187] br[187] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_188 bl[188] br[188] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_189 bl[189] br[189] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_190 bl[190] br[190] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_191 bl[191] br[191] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_192 bl[192] br[192] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_193 bl[193] br[193] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_194 bl[194] br[194] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_195 bl[195] br[195] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_196 bl[196] br[196] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_197 bl[197] br[197] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_198 bl[198] br[198] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_199 bl[199] br[199] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_200 bl[200] br[200] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_201 bl[201] br[201] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_202 bl[202] br[202] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_203 bl[203] br[203] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_204 bl[204] br[204] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_205 bl[205] br[205] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_206 bl[206] br[206] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_207 bl[207] br[207] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_208 bl[208] br[208] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_209 bl[209] br[209] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_210 bl[210] br[210] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_211 bl[211] br[211] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_212 bl[212] br[212] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_213 bl[213] br[213] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_214 bl[214] br[214] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_215 bl[215] br[215] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_216 bl[216] br[216] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_217 bl[217] br[217] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_218 bl[218] br[218] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_219 bl[219] br[219] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_220 bl[220] br[220] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_221 bl[221] br[221] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_222 bl[222] br[222] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_223 bl[223] br[223] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_224 bl[224] br[224] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_225 bl[225] br[225] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_226 bl[226] br[226] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_227 bl[227] br[227] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_228 bl[228] br[228] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_229 bl[229] br[229] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_230 bl[230] br[230] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_231 bl[231] br[231] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_232 bl[232] br[232] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_233 bl[233] br[233] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_234 bl[234] br[234] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_235 bl[235] br[235] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_236 bl[236] br[236] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_237 bl[237] br[237] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_238 bl[238] br[238] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_239 bl[239] br[239] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_240 bl[240] br[240] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_241 bl[241] br[241] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_242 bl[242] br[242] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_243 bl[243] br[243] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_244 bl[244] br[244] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_245 bl[245] br[245] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_246 bl[246] br[246] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_247 bl[247] br[247] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_248 bl[248] br[248] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_249 bl[249] br[249] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_250 bl[250] br[250] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_251 bl[251] br[251] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_252 bl[252] br[252] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_253 bl[253] br[253] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_254 bl[254] br[254] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_255 bl[255] br[255] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_100_0 bl[0] br[0] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_1 bl[1] br[1] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_2 bl[2] br[2] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_3 bl[3] br[3] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_4 bl[4] br[4] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_5 bl[5] br[5] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_6 bl[6] br[6] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_7 bl[7] br[7] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_8 bl[8] br[8] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_9 bl[9] br[9] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_10 bl[10] br[10] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_11 bl[11] br[11] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_12 bl[12] br[12] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_13 bl[13] br[13] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_14 bl[14] br[14] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_15 bl[15] br[15] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_16 bl[16] br[16] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_17 bl[17] br[17] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_18 bl[18] br[18] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_19 bl[19] br[19] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_20 bl[20] br[20] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_21 bl[21] br[21] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_22 bl[22] br[22] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_23 bl[23] br[23] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_24 bl[24] br[24] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_25 bl[25] br[25] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_26 bl[26] br[26] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_27 bl[27] br[27] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_28 bl[28] br[28] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_29 bl[29] br[29] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_30 bl[30] br[30] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_31 bl[31] br[31] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_32 bl[32] br[32] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_33 bl[33] br[33] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_34 bl[34] br[34] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_35 bl[35] br[35] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_36 bl[36] br[36] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_37 bl[37] br[37] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_38 bl[38] br[38] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_39 bl[39] br[39] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_40 bl[40] br[40] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_41 bl[41] br[41] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_42 bl[42] br[42] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_43 bl[43] br[43] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_44 bl[44] br[44] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_45 bl[45] br[45] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_46 bl[46] br[46] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_47 bl[47] br[47] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_48 bl[48] br[48] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_49 bl[49] br[49] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_50 bl[50] br[50] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_51 bl[51] br[51] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_52 bl[52] br[52] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_53 bl[53] br[53] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_54 bl[54] br[54] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_55 bl[55] br[55] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_56 bl[56] br[56] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_57 bl[57] br[57] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_58 bl[58] br[58] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_59 bl[59] br[59] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_60 bl[60] br[60] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_61 bl[61] br[61] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_62 bl[62] br[62] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_63 bl[63] br[63] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_64 bl[64] br[64] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_65 bl[65] br[65] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_66 bl[66] br[66] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_67 bl[67] br[67] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_68 bl[68] br[68] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_69 bl[69] br[69] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_70 bl[70] br[70] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_71 bl[71] br[71] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_72 bl[72] br[72] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_73 bl[73] br[73] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_74 bl[74] br[74] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_75 bl[75] br[75] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_76 bl[76] br[76] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_77 bl[77] br[77] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_78 bl[78] br[78] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_79 bl[79] br[79] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_80 bl[80] br[80] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_81 bl[81] br[81] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_82 bl[82] br[82] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_83 bl[83] br[83] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_84 bl[84] br[84] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_85 bl[85] br[85] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_86 bl[86] br[86] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_87 bl[87] br[87] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_88 bl[88] br[88] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_89 bl[89] br[89] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_90 bl[90] br[90] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_91 bl[91] br[91] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_92 bl[92] br[92] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_93 bl[93] br[93] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_94 bl[94] br[94] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_95 bl[95] br[95] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_96 bl[96] br[96] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_97 bl[97] br[97] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_98 bl[98] br[98] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_99 bl[99] br[99] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_100 bl[100] br[100] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_101 bl[101] br[101] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_102 bl[102] br[102] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_103 bl[103] br[103] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_104 bl[104] br[104] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_105 bl[105] br[105] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_106 bl[106] br[106] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_107 bl[107] br[107] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_108 bl[108] br[108] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_109 bl[109] br[109] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_110 bl[110] br[110] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_111 bl[111] br[111] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_112 bl[112] br[112] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_113 bl[113] br[113] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_114 bl[114] br[114] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_115 bl[115] br[115] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_116 bl[116] br[116] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_117 bl[117] br[117] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_118 bl[118] br[118] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_119 bl[119] br[119] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_120 bl[120] br[120] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_121 bl[121] br[121] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_122 bl[122] br[122] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_123 bl[123] br[123] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_124 bl[124] br[124] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_125 bl[125] br[125] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_126 bl[126] br[126] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_127 bl[127] br[127] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_128 bl[128] br[128] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_129 bl[129] br[129] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_130 bl[130] br[130] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_131 bl[131] br[131] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_132 bl[132] br[132] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_133 bl[133] br[133] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_134 bl[134] br[134] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_135 bl[135] br[135] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_136 bl[136] br[136] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_137 bl[137] br[137] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_138 bl[138] br[138] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_139 bl[139] br[139] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_140 bl[140] br[140] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_141 bl[141] br[141] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_142 bl[142] br[142] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_143 bl[143] br[143] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_144 bl[144] br[144] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_145 bl[145] br[145] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_146 bl[146] br[146] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_147 bl[147] br[147] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_148 bl[148] br[148] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_149 bl[149] br[149] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_150 bl[150] br[150] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_151 bl[151] br[151] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_152 bl[152] br[152] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_153 bl[153] br[153] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_154 bl[154] br[154] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_155 bl[155] br[155] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_156 bl[156] br[156] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_157 bl[157] br[157] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_158 bl[158] br[158] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_159 bl[159] br[159] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_160 bl[160] br[160] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_161 bl[161] br[161] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_162 bl[162] br[162] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_163 bl[163] br[163] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_164 bl[164] br[164] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_165 bl[165] br[165] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_166 bl[166] br[166] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_167 bl[167] br[167] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_168 bl[168] br[168] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_169 bl[169] br[169] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_170 bl[170] br[170] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_171 bl[171] br[171] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_172 bl[172] br[172] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_173 bl[173] br[173] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_174 bl[174] br[174] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_175 bl[175] br[175] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_176 bl[176] br[176] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_177 bl[177] br[177] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_178 bl[178] br[178] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_179 bl[179] br[179] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_180 bl[180] br[180] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_181 bl[181] br[181] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_182 bl[182] br[182] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_183 bl[183] br[183] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_184 bl[184] br[184] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_185 bl[185] br[185] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_186 bl[186] br[186] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_187 bl[187] br[187] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_188 bl[188] br[188] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_189 bl[189] br[189] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_190 bl[190] br[190] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_191 bl[191] br[191] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_192 bl[192] br[192] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_193 bl[193] br[193] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_194 bl[194] br[194] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_195 bl[195] br[195] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_196 bl[196] br[196] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_197 bl[197] br[197] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_198 bl[198] br[198] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_199 bl[199] br[199] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_200 bl[200] br[200] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_201 bl[201] br[201] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_202 bl[202] br[202] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_203 bl[203] br[203] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_204 bl[204] br[204] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_205 bl[205] br[205] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_206 bl[206] br[206] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_207 bl[207] br[207] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_208 bl[208] br[208] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_209 bl[209] br[209] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_210 bl[210] br[210] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_211 bl[211] br[211] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_212 bl[212] br[212] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_213 bl[213] br[213] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_214 bl[214] br[214] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_215 bl[215] br[215] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_216 bl[216] br[216] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_217 bl[217] br[217] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_218 bl[218] br[218] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_219 bl[219] br[219] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_220 bl[220] br[220] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_221 bl[221] br[221] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_222 bl[222] br[222] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_223 bl[223] br[223] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_224 bl[224] br[224] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_225 bl[225] br[225] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_226 bl[226] br[226] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_227 bl[227] br[227] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_228 bl[228] br[228] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_229 bl[229] br[229] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_230 bl[230] br[230] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_231 bl[231] br[231] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_232 bl[232] br[232] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_233 bl[233] br[233] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_234 bl[234] br[234] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_235 bl[235] br[235] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_236 bl[236] br[236] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_237 bl[237] br[237] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_238 bl[238] br[238] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_239 bl[239] br[239] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_240 bl[240] br[240] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_241 bl[241] br[241] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_242 bl[242] br[242] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_243 bl[243] br[243] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_244 bl[244] br[244] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_245 bl[245] br[245] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_246 bl[246] br[246] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_247 bl[247] br[247] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_248 bl[248] br[248] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_249 bl[249] br[249] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_250 bl[250] br[250] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_251 bl[251] br[251] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_252 bl[252] br[252] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_253 bl[253] br[253] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_254 bl[254] br[254] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_255 bl[255] br[255] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_101_0 bl[0] br[0] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_1 bl[1] br[1] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_2 bl[2] br[2] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_3 bl[3] br[3] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_4 bl[4] br[4] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_5 bl[5] br[5] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_6 bl[6] br[6] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_7 bl[7] br[7] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_8 bl[8] br[8] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_9 bl[9] br[9] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_10 bl[10] br[10] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_11 bl[11] br[11] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_12 bl[12] br[12] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_13 bl[13] br[13] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_14 bl[14] br[14] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_15 bl[15] br[15] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_16 bl[16] br[16] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_17 bl[17] br[17] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_18 bl[18] br[18] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_19 bl[19] br[19] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_20 bl[20] br[20] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_21 bl[21] br[21] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_22 bl[22] br[22] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_23 bl[23] br[23] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_24 bl[24] br[24] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_25 bl[25] br[25] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_26 bl[26] br[26] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_27 bl[27] br[27] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_28 bl[28] br[28] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_29 bl[29] br[29] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_30 bl[30] br[30] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_31 bl[31] br[31] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_32 bl[32] br[32] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_33 bl[33] br[33] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_34 bl[34] br[34] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_35 bl[35] br[35] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_36 bl[36] br[36] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_37 bl[37] br[37] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_38 bl[38] br[38] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_39 bl[39] br[39] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_40 bl[40] br[40] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_41 bl[41] br[41] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_42 bl[42] br[42] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_43 bl[43] br[43] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_44 bl[44] br[44] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_45 bl[45] br[45] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_46 bl[46] br[46] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_47 bl[47] br[47] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_48 bl[48] br[48] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_49 bl[49] br[49] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_50 bl[50] br[50] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_51 bl[51] br[51] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_52 bl[52] br[52] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_53 bl[53] br[53] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_54 bl[54] br[54] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_55 bl[55] br[55] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_56 bl[56] br[56] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_57 bl[57] br[57] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_58 bl[58] br[58] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_59 bl[59] br[59] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_60 bl[60] br[60] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_61 bl[61] br[61] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_62 bl[62] br[62] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_63 bl[63] br[63] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_64 bl[64] br[64] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_65 bl[65] br[65] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_66 bl[66] br[66] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_67 bl[67] br[67] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_68 bl[68] br[68] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_69 bl[69] br[69] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_70 bl[70] br[70] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_71 bl[71] br[71] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_72 bl[72] br[72] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_73 bl[73] br[73] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_74 bl[74] br[74] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_75 bl[75] br[75] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_76 bl[76] br[76] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_77 bl[77] br[77] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_78 bl[78] br[78] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_79 bl[79] br[79] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_80 bl[80] br[80] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_81 bl[81] br[81] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_82 bl[82] br[82] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_83 bl[83] br[83] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_84 bl[84] br[84] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_85 bl[85] br[85] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_86 bl[86] br[86] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_87 bl[87] br[87] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_88 bl[88] br[88] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_89 bl[89] br[89] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_90 bl[90] br[90] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_91 bl[91] br[91] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_92 bl[92] br[92] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_93 bl[93] br[93] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_94 bl[94] br[94] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_95 bl[95] br[95] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_96 bl[96] br[96] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_97 bl[97] br[97] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_98 bl[98] br[98] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_99 bl[99] br[99] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_100 bl[100] br[100] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_101 bl[101] br[101] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_102 bl[102] br[102] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_103 bl[103] br[103] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_104 bl[104] br[104] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_105 bl[105] br[105] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_106 bl[106] br[106] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_107 bl[107] br[107] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_108 bl[108] br[108] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_109 bl[109] br[109] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_110 bl[110] br[110] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_111 bl[111] br[111] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_112 bl[112] br[112] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_113 bl[113] br[113] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_114 bl[114] br[114] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_115 bl[115] br[115] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_116 bl[116] br[116] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_117 bl[117] br[117] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_118 bl[118] br[118] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_119 bl[119] br[119] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_120 bl[120] br[120] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_121 bl[121] br[121] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_122 bl[122] br[122] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_123 bl[123] br[123] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_124 bl[124] br[124] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_125 bl[125] br[125] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_126 bl[126] br[126] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_127 bl[127] br[127] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_128 bl[128] br[128] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_129 bl[129] br[129] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_130 bl[130] br[130] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_131 bl[131] br[131] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_132 bl[132] br[132] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_133 bl[133] br[133] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_134 bl[134] br[134] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_135 bl[135] br[135] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_136 bl[136] br[136] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_137 bl[137] br[137] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_138 bl[138] br[138] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_139 bl[139] br[139] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_140 bl[140] br[140] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_141 bl[141] br[141] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_142 bl[142] br[142] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_143 bl[143] br[143] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_144 bl[144] br[144] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_145 bl[145] br[145] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_146 bl[146] br[146] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_147 bl[147] br[147] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_148 bl[148] br[148] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_149 bl[149] br[149] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_150 bl[150] br[150] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_151 bl[151] br[151] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_152 bl[152] br[152] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_153 bl[153] br[153] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_154 bl[154] br[154] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_155 bl[155] br[155] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_156 bl[156] br[156] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_157 bl[157] br[157] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_158 bl[158] br[158] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_159 bl[159] br[159] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_160 bl[160] br[160] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_161 bl[161] br[161] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_162 bl[162] br[162] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_163 bl[163] br[163] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_164 bl[164] br[164] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_165 bl[165] br[165] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_166 bl[166] br[166] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_167 bl[167] br[167] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_168 bl[168] br[168] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_169 bl[169] br[169] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_170 bl[170] br[170] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_171 bl[171] br[171] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_172 bl[172] br[172] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_173 bl[173] br[173] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_174 bl[174] br[174] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_175 bl[175] br[175] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_176 bl[176] br[176] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_177 bl[177] br[177] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_178 bl[178] br[178] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_179 bl[179] br[179] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_180 bl[180] br[180] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_181 bl[181] br[181] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_182 bl[182] br[182] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_183 bl[183] br[183] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_184 bl[184] br[184] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_185 bl[185] br[185] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_186 bl[186] br[186] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_187 bl[187] br[187] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_188 bl[188] br[188] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_189 bl[189] br[189] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_190 bl[190] br[190] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_191 bl[191] br[191] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_192 bl[192] br[192] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_193 bl[193] br[193] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_194 bl[194] br[194] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_195 bl[195] br[195] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_196 bl[196] br[196] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_197 bl[197] br[197] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_198 bl[198] br[198] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_199 bl[199] br[199] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_200 bl[200] br[200] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_201 bl[201] br[201] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_202 bl[202] br[202] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_203 bl[203] br[203] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_204 bl[204] br[204] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_205 bl[205] br[205] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_206 bl[206] br[206] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_207 bl[207] br[207] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_208 bl[208] br[208] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_209 bl[209] br[209] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_210 bl[210] br[210] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_211 bl[211] br[211] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_212 bl[212] br[212] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_213 bl[213] br[213] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_214 bl[214] br[214] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_215 bl[215] br[215] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_216 bl[216] br[216] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_217 bl[217] br[217] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_218 bl[218] br[218] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_219 bl[219] br[219] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_220 bl[220] br[220] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_221 bl[221] br[221] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_222 bl[222] br[222] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_223 bl[223] br[223] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_224 bl[224] br[224] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_225 bl[225] br[225] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_226 bl[226] br[226] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_227 bl[227] br[227] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_228 bl[228] br[228] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_229 bl[229] br[229] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_230 bl[230] br[230] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_231 bl[231] br[231] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_232 bl[232] br[232] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_233 bl[233] br[233] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_234 bl[234] br[234] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_235 bl[235] br[235] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_236 bl[236] br[236] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_237 bl[237] br[237] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_238 bl[238] br[238] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_239 bl[239] br[239] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_240 bl[240] br[240] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_241 bl[241] br[241] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_242 bl[242] br[242] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_243 bl[243] br[243] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_244 bl[244] br[244] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_245 bl[245] br[245] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_246 bl[246] br[246] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_247 bl[247] br[247] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_248 bl[248] br[248] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_249 bl[249] br[249] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_250 bl[250] br[250] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_251 bl[251] br[251] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_252 bl[252] br[252] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_253 bl[253] br[253] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_254 bl[254] br[254] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_255 bl[255] br[255] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_102_0 bl[0] br[0] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_1 bl[1] br[1] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_2 bl[2] br[2] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_3 bl[3] br[3] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_4 bl[4] br[4] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_5 bl[5] br[5] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_6 bl[6] br[6] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_7 bl[7] br[7] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_8 bl[8] br[8] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_9 bl[9] br[9] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_10 bl[10] br[10] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_11 bl[11] br[11] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_12 bl[12] br[12] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_13 bl[13] br[13] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_14 bl[14] br[14] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_15 bl[15] br[15] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_16 bl[16] br[16] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_17 bl[17] br[17] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_18 bl[18] br[18] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_19 bl[19] br[19] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_20 bl[20] br[20] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_21 bl[21] br[21] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_22 bl[22] br[22] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_23 bl[23] br[23] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_24 bl[24] br[24] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_25 bl[25] br[25] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_26 bl[26] br[26] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_27 bl[27] br[27] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_28 bl[28] br[28] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_29 bl[29] br[29] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_30 bl[30] br[30] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_31 bl[31] br[31] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_32 bl[32] br[32] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_33 bl[33] br[33] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_34 bl[34] br[34] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_35 bl[35] br[35] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_36 bl[36] br[36] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_37 bl[37] br[37] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_38 bl[38] br[38] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_39 bl[39] br[39] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_40 bl[40] br[40] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_41 bl[41] br[41] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_42 bl[42] br[42] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_43 bl[43] br[43] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_44 bl[44] br[44] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_45 bl[45] br[45] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_46 bl[46] br[46] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_47 bl[47] br[47] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_48 bl[48] br[48] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_49 bl[49] br[49] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_50 bl[50] br[50] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_51 bl[51] br[51] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_52 bl[52] br[52] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_53 bl[53] br[53] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_54 bl[54] br[54] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_55 bl[55] br[55] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_56 bl[56] br[56] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_57 bl[57] br[57] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_58 bl[58] br[58] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_59 bl[59] br[59] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_60 bl[60] br[60] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_61 bl[61] br[61] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_62 bl[62] br[62] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_63 bl[63] br[63] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_64 bl[64] br[64] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_65 bl[65] br[65] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_66 bl[66] br[66] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_67 bl[67] br[67] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_68 bl[68] br[68] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_69 bl[69] br[69] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_70 bl[70] br[70] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_71 bl[71] br[71] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_72 bl[72] br[72] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_73 bl[73] br[73] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_74 bl[74] br[74] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_75 bl[75] br[75] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_76 bl[76] br[76] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_77 bl[77] br[77] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_78 bl[78] br[78] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_79 bl[79] br[79] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_80 bl[80] br[80] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_81 bl[81] br[81] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_82 bl[82] br[82] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_83 bl[83] br[83] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_84 bl[84] br[84] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_85 bl[85] br[85] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_86 bl[86] br[86] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_87 bl[87] br[87] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_88 bl[88] br[88] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_89 bl[89] br[89] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_90 bl[90] br[90] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_91 bl[91] br[91] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_92 bl[92] br[92] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_93 bl[93] br[93] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_94 bl[94] br[94] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_95 bl[95] br[95] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_96 bl[96] br[96] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_97 bl[97] br[97] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_98 bl[98] br[98] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_99 bl[99] br[99] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_100 bl[100] br[100] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_101 bl[101] br[101] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_102 bl[102] br[102] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_103 bl[103] br[103] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_104 bl[104] br[104] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_105 bl[105] br[105] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_106 bl[106] br[106] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_107 bl[107] br[107] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_108 bl[108] br[108] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_109 bl[109] br[109] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_110 bl[110] br[110] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_111 bl[111] br[111] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_112 bl[112] br[112] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_113 bl[113] br[113] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_114 bl[114] br[114] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_115 bl[115] br[115] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_116 bl[116] br[116] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_117 bl[117] br[117] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_118 bl[118] br[118] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_119 bl[119] br[119] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_120 bl[120] br[120] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_121 bl[121] br[121] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_122 bl[122] br[122] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_123 bl[123] br[123] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_124 bl[124] br[124] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_125 bl[125] br[125] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_126 bl[126] br[126] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_127 bl[127] br[127] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_128 bl[128] br[128] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_129 bl[129] br[129] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_130 bl[130] br[130] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_131 bl[131] br[131] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_132 bl[132] br[132] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_133 bl[133] br[133] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_134 bl[134] br[134] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_135 bl[135] br[135] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_136 bl[136] br[136] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_137 bl[137] br[137] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_138 bl[138] br[138] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_139 bl[139] br[139] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_140 bl[140] br[140] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_141 bl[141] br[141] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_142 bl[142] br[142] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_143 bl[143] br[143] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_144 bl[144] br[144] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_145 bl[145] br[145] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_146 bl[146] br[146] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_147 bl[147] br[147] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_148 bl[148] br[148] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_149 bl[149] br[149] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_150 bl[150] br[150] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_151 bl[151] br[151] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_152 bl[152] br[152] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_153 bl[153] br[153] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_154 bl[154] br[154] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_155 bl[155] br[155] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_156 bl[156] br[156] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_157 bl[157] br[157] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_158 bl[158] br[158] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_159 bl[159] br[159] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_160 bl[160] br[160] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_161 bl[161] br[161] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_162 bl[162] br[162] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_163 bl[163] br[163] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_164 bl[164] br[164] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_165 bl[165] br[165] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_166 bl[166] br[166] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_167 bl[167] br[167] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_168 bl[168] br[168] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_169 bl[169] br[169] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_170 bl[170] br[170] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_171 bl[171] br[171] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_172 bl[172] br[172] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_173 bl[173] br[173] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_174 bl[174] br[174] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_175 bl[175] br[175] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_176 bl[176] br[176] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_177 bl[177] br[177] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_178 bl[178] br[178] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_179 bl[179] br[179] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_180 bl[180] br[180] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_181 bl[181] br[181] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_182 bl[182] br[182] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_183 bl[183] br[183] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_184 bl[184] br[184] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_185 bl[185] br[185] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_186 bl[186] br[186] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_187 bl[187] br[187] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_188 bl[188] br[188] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_189 bl[189] br[189] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_190 bl[190] br[190] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_191 bl[191] br[191] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_192 bl[192] br[192] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_193 bl[193] br[193] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_194 bl[194] br[194] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_195 bl[195] br[195] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_196 bl[196] br[196] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_197 bl[197] br[197] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_198 bl[198] br[198] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_199 bl[199] br[199] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_200 bl[200] br[200] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_201 bl[201] br[201] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_202 bl[202] br[202] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_203 bl[203] br[203] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_204 bl[204] br[204] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_205 bl[205] br[205] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_206 bl[206] br[206] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_207 bl[207] br[207] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_208 bl[208] br[208] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_209 bl[209] br[209] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_210 bl[210] br[210] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_211 bl[211] br[211] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_212 bl[212] br[212] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_213 bl[213] br[213] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_214 bl[214] br[214] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_215 bl[215] br[215] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_216 bl[216] br[216] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_217 bl[217] br[217] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_218 bl[218] br[218] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_219 bl[219] br[219] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_220 bl[220] br[220] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_221 bl[221] br[221] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_222 bl[222] br[222] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_223 bl[223] br[223] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_224 bl[224] br[224] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_225 bl[225] br[225] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_226 bl[226] br[226] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_227 bl[227] br[227] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_228 bl[228] br[228] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_229 bl[229] br[229] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_230 bl[230] br[230] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_231 bl[231] br[231] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_232 bl[232] br[232] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_233 bl[233] br[233] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_234 bl[234] br[234] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_235 bl[235] br[235] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_236 bl[236] br[236] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_237 bl[237] br[237] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_238 bl[238] br[238] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_239 bl[239] br[239] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_240 bl[240] br[240] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_241 bl[241] br[241] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_242 bl[242] br[242] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_243 bl[243] br[243] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_244 bl[244] br[244] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_245 bl[245] br[245] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_246 bl[246] br[246] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_247 bl[247] br[247] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_248 bl[248] br[248] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_249 bl[249] br[249] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_250 bl[250] br[250] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_251 bl[251] br[251] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_252 bl[252] br[252] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_253 bl[253] br[253] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_254 bl[254] br[254] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_255 bl[255] br[255] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_103_0 bl[0] br[0] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_1 bl[1] br[1] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_2 bl[2] br[2] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_3 bl[3] br[3] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_4 bl[4] br[4] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_5 bl[5] br[5] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_6 bl[6] br[6] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_7 bl[7] br[7] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_8 bl[8] br[8] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_9 bl[9] br[9] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_10 bl[10] br[10] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_11 bl[11] br[11] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_12 bl[12] br[12] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_13 bl[13] br[13] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_14 bl[14] br[14] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_15 bl[15] br[15] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_16 bl[16] br[16] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_17 bl[17] br[17] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_18 bl[18] br[18] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_19 bl[19] br[19] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_20 bl[20] br[20] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_21 bl[21] br[21] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_22 bl[22] br[22] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_23 bl[23] br[23] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_24 bl[24] br[24] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_25 bl[25] br[25] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_26 bl[26] br[26] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_27 bl[27] br[27] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_28 bl[28] br[28] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_29 bl[29] br[29] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_30 bl[30] br[30] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_31 bl[31] br[31] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_32 bl[32] br[32] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_33 bl[33] br[33] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_34 bl[34] br[34] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_35 bl[35] br[35] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_36 bl[36] br[36] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_37 bl[37] br[37] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_38 bl[38] br[38] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_39 bl[39] br[39] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_40 bl[40] br[40] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_41 bl[41] br[41] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_42 bl[42] br[42] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_43 bl[43] br[43] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_44 bl[44] br[44] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_45 bl[45] br[45] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_46 bl[46] br[46] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_47 bl[47] br[47] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_48 bl[48] br[48] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_49 bl[49] br[49] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_50 bl[50] br[50] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_51 bl[51] br[51] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_52 bl[52] br[52] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_53 bl[53] br[53] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_54 bl[54] br[54] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_55 bl[55] br[55] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_56 bl[56] br[56] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_57 bl[57] br[57] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_58 bl[58] br[58] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_59 bl[59] br[59] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_60 bl[60] br[60] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_61 bl[61] br[61] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_62 bl[62] br[62] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_63 bl[63] br[63] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_64 bl[64] br[64] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_65 bl[65] br[65] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_66 bl[66] br[66] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_67 bl[67] br[67] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_68 bl[68] br[68] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_69 bl[69] br[69] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_70 bl[70] br[70] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_71 bl[71] br[71] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_72 bl[72] br[72] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_73 bl[73] br[73] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_74 bl[74] br[74] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_75 bl[75] br[75] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_76 bl[76] br[76] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_77 bl[77] br[77] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_78 bl[78] br[78] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_79 bl[79] br[79] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_80 bl[80] br[80] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_81 bl[81] br[81] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_82 bl[82] br[82] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_83 bl[83] br[83] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_84 bl[84] br[84] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_85 bl[85] br[85] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_86 bl[86] br[86] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_87 bl[87] br[87] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_88 bl[88] br[88] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_89 bl[89] br[89] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_90 bl[90] br[90] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_91 bl[91] br[91] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_92 bl[92] br[92] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_93 bl[93] br[93] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_94 bl[94] br[94] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_95 bl[95] br[95] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_96 bl[96] br[96] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_97 bl[97] br[97] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_98 bl[98] br[98] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_99 bl[99] br[99] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_100 bl[100] br[100] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_101 bl[101] br[101] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_102 bl[102] br[102] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_103 bl[103] br[103] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_104 bl[104] br[104] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_105 bl[105] br[105] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_106 bl[106] br[106] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_107 bl[107] br[107] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_108 bl[108] br[108] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_109 bl[109] br[109] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_110 bl[110] br[110] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_111 bl[111] br[111] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_112 bl[112] br[112] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_113 bl[113] br[113] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_114 bl[114] br[114] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_115 bl[115] br[115] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_116 bl[116] br[116] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_117 bl[117] br[117] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_118 bl[118] br[118] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_119 bl[119] br[119] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_120 bl[120] br[120] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_121 bl[121] br[121] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_122 bl[122] br[122] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_123 bl[123] br[123] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_124 bl[124] br[124] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_125 bl[125] br[125] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_126 bl[126] br[126] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_127 bl[127] br[127] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_128 bl[128] br[128] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_129 bl[129] br[129] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_130 bl[130] br[130] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_131 bl[131] br[131] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_132 bl[132] br[132] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_133 bl[133] br[133] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_134 bl[134] br[134] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_135 bl[135] br[135] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_136 bl[136] br[136] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_137 bl[137] br[137] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_138 bl[138] br[138] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_139 bl[139] br[139] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_140 bl[140] br[140] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_141 bl[141] br[141] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_142 bl[142] br[142] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_143 bl[143] br[143] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_144 bl[144] br[144] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_145 bl[145] br[145] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_146 bl[146] br[146] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_147 bl[147] br[147] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_148 bl[148] br[148] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_149 bl[149] br[149] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_150 bl[150] br[150] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_151 bl[151] br[151] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_152 bl[152] br[152] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_153 bl[153] br[153] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_154 bl[154] br[154] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_155 bl[155] br[155] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_156 bl[156] br[156] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_157 bl[157] br[157] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_158 bl[158] br[158] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_159 bl[159] br[159] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_160 bl[160] br[160] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_161 bl[161] br[161] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_162 bl[162] br[162] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_163 bl[163] br[163] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_164 bl[164] br[164] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_165 bl[165] br[165] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_166 bl[166] br[166] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_167 bl[167] br[167] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_168 bl[168] br[168] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_169 bl[169] br[169] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_170 bl[170] br[170] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_171 bl[171] br[171] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_172 bl[172] br[172] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_173 bl[173] br[173] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_174 bl[174] br[174] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_175 bl[175] br[175] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_176 bl[176] br[176] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_177 bl[177] br[177] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_178 bl[178] br[178] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_179 bl[179] br[179] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_180 bl[180] br[180] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_181 bl[181] br[181] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_182 bl[182] br[182] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_183 bl[183] br[183] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_184 bl[184] br[184] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_185 bl[185] br[185] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_186 bl[186] br[186] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_187 bl[187] br[187] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_188 bl[188] br[188] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_189 bl[189] br[189] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_190 bl[190] br[190] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_191 bl[191] br[191] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_192 bl[192] br[192] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_193 bl[193] br[193] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_194 bl[194] br[194] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_195 bl[195] br[195] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_196 bl[196] br[196] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_197 bl[197] br[197] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_198 bl[198] br[198] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_199 bl[199] br[199] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_200 bl[200] br[200] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_201 bl[201] br[201] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_202 bl[202] br[202] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_203 bl[203] br[203] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_204 bl[204] br[204] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_205 bl[205] br[205] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_206 bl[206] br[206] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_207 bl[207] br[207] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_208 bl[208] br[208] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_209 bl[209] br[209] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_210 bl[210] br[210] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_211 bl[211] br[211] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_212 bl[212] br[212] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_213 bl[213] br[213] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_214 bl[214] br[214] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_215 bl[215] br[215] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_216 bl[216] br[216] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_217 bl[217] br[217] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_218 bl[218] br[218] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_219 bl[219] br[219] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_220 bl[220] br[220] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_221 bl[221] br[221] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_222 bl[222] br[222] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_223 bl[223] br[223] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_224 bl[224] br[224] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_225 bl[225] br[225] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_226 bl[226] br[226] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_227 bl[227] br[227] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_228 bl[228] br[228] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_229 bl[229] br[229] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_230 bl[230] br[230] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_231 bl[231] br[231] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_232 bl[232] br[232] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_233 bl[233] br[233] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_234 bl[234] br[234] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_235 bl[235] br[235] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_236 bl[236] br[236] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_237 bl[237] br[237] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_238 bl[238] br[238] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_239 bl[239] br[239] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_240 bl[240] br[240] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_241 bl[241] br[241] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_242 bl[242] br[242] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_243 bl[243] br[243] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_244 bl[244] br[244] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_245 bl[245] br[245] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_246 bl[246] br[246] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_247 bl[247] br[247] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_248 bl[248] br[248] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_249 bl[249] br[249] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_250 bl[250] br[250] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_251 bl[251] br[251] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_252 bl[252] br[252] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_253 bl[253] br[253] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_254 bl[254] br[254] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_255 bl[255] br[255] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_104_0 bl[0] br[0] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_1 bl[1] br[1] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_2 bl[2] br[2] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_3 bl[3] br[3] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_4 bl[4] br[4] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_5 bl[5] br[5] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_6 bl[6] br[6] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_7 bl[7] br[7] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_8 bl[8] br[8] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_9 bl[9] br[9] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_10 bl[10] br[10] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_11 bl[11] br[11] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_12 bl[12] br[12] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_13 bl[13] br[13] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_14 bl[14] br[14] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_15 bl[15] br[15] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_16 bl[16] br[16] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_17 bl[17] br[17] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_18 bl[18] br[18] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_19 bl[19] br[19] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_20 bl[20] br[20] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_21 bl[21] br[21] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_22 bl[22] br[22] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_23 bl[23] br[23] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_24 bl[24] br[24] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_25 bl[25] br[25] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_26 bl[26] br[26] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_27 bl[27] br[27] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_28 bl[28] br[28] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_29 bl[29] br[29] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_30 bl[30] br[30] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_31 bl[31] br[31] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_32 bl[32] br[32] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_33 bl[33] br[33] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_34 bl[34] br[34] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_35 bl[35] br[35] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_36 bl[36] br[36] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_37 bl[37] br[37] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_38 bl[38] br[38] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_39 bl[39] br[39] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_40 bl[40] br[40] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_41 bl[41] br[41] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_42 bl[42] br[42] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_43 bl[43] br[43] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_44 bl[44] br[44] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_45 bl[45] br[45] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_46 bl[46] br[46] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_47 bl[47] br[47] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_48 bl[48] br[48] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_49 bl[49] br[49] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_50 bl[50] br[50] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_51 bl[51] br[51] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_52 bl[52] br[52] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_53 bl[53] br[53] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_54 bl[54] br[54] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_55 bl[55] br[55] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_56 bl[56] br[56] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_57 bl[57] br[57] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_58 bl[58] br[58] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_59 bl[59] br[59] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_60 bl[60] br[60] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_61 bl[61] br[61] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_62 bl[62] br[62] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_63 bl[63] br[63] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_64 bl[64] br[64] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_65 bl[65] br[65] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_66 bl[66] br[66] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_67 bl[67] br[67] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_68 bl[68] br[68] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_69 bl[69] br[69] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_70 bl[70] br[70] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_71 bl[71] br[71] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_72 bl[72] br[72] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_73 bl[73] br[73] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_74 bl[74] br[74] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_75 bl[75] br[75] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_76 bl[76] br[76] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_77 bl[77] br[77] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_78 bl[78] br[78] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_79 bl[79] br[79] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_80 bl[80] br[80] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_81 bl[81] br[81] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_82 bl[82] br[82] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_83 bl[83] br[83] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_84 bl[84] br[84] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_85 bl[85] br[85] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_86 bl[86] br[86] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_87 bl[87] br[87] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_88 bl[88] br[88] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_89 bl[89] br[89] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_90 bl[90] br[90] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_91 bl[91] br[91] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_92 bl[92] br[92] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_93 bl[93] br[93] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_94 bl[94] br[94] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_95 bl[95] br[95] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_96 bl[96] br[96] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_97 bl[97] br[97] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_98 bl[98] br[98] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_99 bl[99] br[99] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_100 bl[100] br[100] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_101 bl[101] br[101] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_102 bl[102] br[102] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_103 bl[103] br[103] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_104 bl[104] br[104] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_105 bl[105] br[105] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_106 bl[106] br[106] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_107 bl[107] br[107] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_108 bl[108] br[108] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_109 bl[109] br[109] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_110 bl[110] br[110] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_111 bl[111] br[111] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_112 bl[112] br[112] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_113 bl[113] br[113] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_114 bl[114] br[114] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_115 bl[115] br[115] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_116 bl[116] br[116] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_117 bl[117] br[117] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_118 bl[118] br[118] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_119 bl[119] br[119] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_120 bl[120] br[120] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_121 bl[121] br[121] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_122 bl[122] br[122] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_123 bl[123] br[123] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_124 bl[124] br[124] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_125 bl[125] br[125] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_126 bl[126] br[126] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_127 bl[127] br[127] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_128 bl[128] br[128] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_129 bl[129] br[129] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_130 bl[130] br[130] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_131 bl[131] br[131] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_132 bl[132] br[132] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_133 bl[133] br[133] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_134 bl[134] br[134] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_135 bl[135] br[135] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_136 bl[136] br[136] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_137 bl[137] br[137] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_138 bl[138] br[138] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_139 bl[139] br[139] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_140 bl[140] br[140] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_141 bl[141] br[141] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_142 bl[142] br[142] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_143 bl[143] br[143] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_144 bl[144] br[144] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_145 bl[145] br[145] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_146 bl[146] br[146] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_147 bl[147] br[147] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_148 bl[148] br[148] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_149 bl[149] br[149] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_150 bl[150] br[150] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_151 bl[151] br[151] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_152 bl[152] br[152] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_153 bl[153] br[153] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_154 bl[154] br[154] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_155 bl[155] br[155] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_156 bl[156] br[156] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_157 bl[157] br[157] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_158 bl[158] br[158] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_159 bl[159] br[159] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_160 bl[160] br[160] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_161 bl[161] br[161] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_162 bl[162] br[162] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_163 bl[163] br[163] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_164 bl[164] br[164] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_165 bl[165] br[165] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_166 bl[166] br[166] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_167 bl[167] br[167] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_168 bl[168] br[168] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_169 bl[169] br[169] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_170 bl[170] br[170] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_171 bl[171] br[171] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_172 bl[172] br[172] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_173 bl[173] br[173] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_174 bl[174] br[174] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_175 bl[175] br[175] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_176 bl[176] br[176] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_177 bl[177] br[177] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_178 bl[178] br[178] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_179 bl[179] br[179] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_180 bl[180] br[180] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_181 bl[181] br[181] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_182 bl[182] br[182] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_183 bl[183] br[183] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_184 bl[184] br[184] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_185 bl[185] br[185] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_186 bl[186] br[186] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_187 bl[187] br[187] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_188 bl[188] br[188] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_189 bl[189] br[189] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_190 bl[190] br[190] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_191 bl[191] br[191] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_192 bl[192] br[192] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_193 bl[193] br[193] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_194 bl[194] br[194] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_195 bl[195] br[195] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_196 bl[196] br[196] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_197 bl[197] br[197] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_198 bl[198] br[198] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_199 bl[199] br[199] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_200 bl[200] br[200] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_201 bl[201] br[201] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_202 bl[202] br[202] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_203 bl[203] br[203] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_204 bl[204] br[204] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_205 bl[205] br[205] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_206 bl[206] br[206] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_207 bl[207] br[207] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_208 bl[208] br[208] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_209 bl[209] br[209] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_210 bl[210] br[210] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_211 bl[211] br[211] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_212 bl[212] br[212] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_213 bl[213] br[213] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_214 bl[214] br[214] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_215 bl[215] br[215] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_216 bl[216] br[216] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_217 bl[217] br[217] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_218 bl[218] br[218] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_219 bl[219] br[219] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_220 bl[220] br[220] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_221 bl[221] br[221] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_222 bl[222] br[222] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_223 bl[223] br[223] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_224 bl[224] br[224] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_225 bl[225] br[225] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_226 bl[226] br[226] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_227 bl[227] br[227] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_228 bl[228] br[228] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_229 bl[229] br[229] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_230 bl[230] br[230] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_231 bl[231] br[231] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_232 bl[232] br[232] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_233 bl[233] br[233] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_234 bl[234] br[234] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_235 bl[235] br[235] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_236 bl[236] br[236] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_237 bl[237] br[237] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_238 bl[238] br[238] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_239 bl[239] br[239] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_240 bl[240] br[240] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_241 bl[241] br[241] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_242 bl[242] br[242] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_243 bl[243] br[243] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_244 bl[244] br[244] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_245 bl[245] br[245] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_246 bl[246] br[246] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_247 bl[247] br[247] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_248 bl[248] br[248] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_249 bl[249] br[249] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_250 bl[250] br[250] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_251 bl[251] br[251] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_252 bl[252] br[252] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_253 bl[253] br[253] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_254 bl[254] br[254] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_255 bl[255] br[255] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_105_0 bl[0] br[0] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_1 bl[1] br[1] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_2 bl[2] br[2] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_3 bl[3] br[3] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_4 bl[4] br[4] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_5 bl[5] br[5] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_6 bl[6] br[6] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_7 bl[7] br[7] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_8 bl[8] br[8] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_9 bl[9] br[9] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_10 bl[10] br[10] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_11 bl[11] br[11] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_12 bl[12] br[12] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_13 bl[13] br[13] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_14 bl[14] br[14] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_15 bl[15] br[15] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_16 bl[16] br[16] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_17 bl[17] br[17] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_18 bl[18] br[18] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_19 bl[19] br[19] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_20 bl[20] br[20] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_21 bl[21] br[21] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_22 bl[22] br[22] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_23 bl[23] br[23] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_24 bl[24] br[24] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_25 bl[25] br[25] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_26 bl[26] br[26] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_27 bl[27] br[27] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_28 bl[28] br[28] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_29 bl[29] br[29] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_30 bl[30] br[30] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_31 bl[31] br[31] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_32 bl[32] br[32] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_33 bl[33] br[33] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_34 bl[34] br[34] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_35 bl[35] br[35] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_36 bl[36] br[36] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_37 bl[37] br[37] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_38 bl[38] br[38] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_39 bl[39] br[39] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_40 bl[40] br[40] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_41 bl[41] br[41] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_42 bl[42] br[42] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_43 bl[43] br[43] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_44 bl[44] br[44] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_45 bl[45] br[45] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_46 bl[46] br[46] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_47 bl[47] br[47] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_48 bl[48] br[48] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_49 bl[49] br[49] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_50 bl[50] br[50] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_51 bl[51] br[51] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_52 bl[52] br[52] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_53 bl[53] br[53] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_54 bl[54] br[54] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_55 bl[55] br[55] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_56 bl[56] br[56] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_57 bl[57] br[57] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_58 bl[58] br[58] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_59 bl[59] br[59] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_60 bl[60] br[60] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_61 bl[61] br[61] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_62 bl[62] br[62] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_63 bl[63] br[63] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_64 bl[64] br[64] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_65 bl[65] br[65] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_66 bl[66] br[66] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_67 bl[67] br[67] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_68 bl[68] br[68] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_69 bl[69] br[69] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_70 bl[70] br[70] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_71 bl[71] br[71] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_72 bl[72] br[72] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_73 bl[73] br[73] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_74 bl[74] br[74] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_75 bl[75] br[75] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_76 bl[76] br[76] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_77 bl[77] br[77] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_78 bl[78] br[78] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_79 bl[79] br[79] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_80 bl[80] br[80] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_81 bl[81] br[81] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_82 bl[82] br[82] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_83 bl[83] br[83] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_84 bl[84] br[84] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_85 bl[85] br[85] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_86 bl[86] br[86] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_87 bl[87] br[87] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_88 bl[88] br[88] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_89 bl[89] br[89] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_90 bl[90] br[90] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_91 bl[91] br[91] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_92 bl[92] br[92] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_93 bl[93] br[93] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_94 bl[94] br[94] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_95 bl[95] br[95] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_96 bl[96] br[96] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_97 bl[97] br[97] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_98 bl[98] br[98] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_99 bl[99] br[99] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_100 bl[100] br[100] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_101 bl[101] br[101] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_102 bl[102] br[102] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_103 bl[103] br[103] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_104 bl[104] br[104] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_105 bl[105] br[105] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_106 bl[106] br[106] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_107 bl[107] br[107] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_108 bl[108] br[108] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_109 bl[109] br[109] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_110 bl[110] br[110] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_111 bl[111] br[111] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_112 bl[112] br[112] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_113 bl[113] br[113] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_114 bl[114] br[114] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_115 bl[115] br[115] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_116 bl[116] br[116] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_117 bl[117] br[117] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_118 bl[118] br[118] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_119 bl[119] br[119] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_120 bl[120] br[120] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_121 bl[121] br[121] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_122 bl[122] br[122] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_123 bl[123] br[123] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_124 bl[124] br[124] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_125 bl[125] br[125] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_126 bl[126] br[126] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_127 bl[127] br[127] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_128 bl[128] br[128] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_129 bl[129] br[129] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_130 bl[130] br[130] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_131 bl[131] br[131] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_132 bl[132] br[132] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_133 bl[133] br[133] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_134 bl[134] br[134] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_135 bl[135] br[135] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_136 bl[136] br[136] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_137 bl[137] br[137] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_138 bl[138] br[138] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_139 bl[139] br[139] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_140 bl[140] br[140] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_141 bl[141] br[141] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_142 bl[142] br[142] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_143 bl[143] br[143] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_144 bl[144] br[144] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_145 bl[145] br[145] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_146 bl[146] br[146] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_147 bl[147] br[147] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_148 bl[148] br[148] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_149 bl[149] br[149] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_150 bl[150] br[150] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_151 bl[151] br[151] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_152 bl[152] br[152] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_153 bl[153] br[153] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_154 bl[154] br[154] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_155 bl[155] br[155] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_156 bl[156] br[156] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_157 bl[157] br[157] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_158 bl[158] br[158] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_159 bl[159] br[159] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_160 bl[160] br[160] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_161 bl[161] br[161] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_162 bl[162] br[162] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_163 bl[163] br[163] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_164 bl[164] br[164] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_165 bl[165] br[165] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_166 bl[166] br[166] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_167 bl[167] br[167] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_168 bl[168] br[168] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_169 bl[169] br[169] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_170 bl[170] br[170] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_171 bl[171] br[171] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_172 bl[172] br[172] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_173 bl[173] br[173] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_174 bl[174] br[174] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_175 bl[175] br[175] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_176 bl[176] br[176] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_177 bl[177] br[177] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_178 bl[178] br[178] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_179 bl[179] br[179] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_180 bl[180] br[180] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_181 bl[181] br[181] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_182 bl[182] br[182] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_183 bl[183] br[183] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_184 bl[184] br[184] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_185 bl[185] br[185] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_186 bl[186] br[186] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_187 bl[187] br[187] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_188 bl[188] br[188] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_189 bl[189] br[189] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_190 bl[190] br[190] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_191 bl[191] br[191] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_192 bl[192] br[192] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_193 bl[193] br[193] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_194 bl[194] br[194] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_195 bl[195] br[195] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_196 bl[196] br[196] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_197 bl[197] br[197] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_198 bl[198] br[198] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_199 bl[199] br[199] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_200 bl[200] br[200] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_201 bl[201] br[201] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_202 bl[202] br[202] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_203 bl[203] br[203] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_204 bl[204] br[204] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_205 bl[205] br[205] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_206 bl[206] br[206] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_207 bl[207] br[207] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_208 bl[208] br[208] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_209 bl[209] br[209] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_210 bl[210] br[210] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_211 bl[211] br[211] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_212 bl[212] br[212] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_213 bl[213] br[213] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_214 bl[214] br[214] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_215 bl[215] br[215] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_216 bl[216] br[216] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_217 bl[217] br[217] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_218 bl[218] br[218] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_219 bl[219] br[219] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_220 bl[220] br[220] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_221 bl[221] br[221] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_222 bl[222] br[222] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_223 bl[223] br[223] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_224 bl[224] br[224] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_225 bl[225] br[225] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_226 bl[226] br[226] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_227 bl[227] br[227] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_228 bl[228] br[228] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_229 bl[229] br[229] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_230 bl[230] br[230] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_231 bl[231] br[231] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_232 bl[232] br[232] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_233 bl[233] br[233] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_234 bl[234] br[234] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_235 bl[235] br[235] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_236 bl[236] br[236] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_237 bl[237] br[237] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_238 bl[238] br[238] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_239 bl[239] br[239] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_240 bl[240] br[240] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_241 bl[241] br[241] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_242 bl[242] br[242] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_243 bl[243] br[243] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_244 bl[244] br[244] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_245 bl[245] br[245] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_246 bl[246] br[246] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_247 bl[247] br[247] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_248 bl[248] br[248] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_249 bl[249] br[249] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_250 bl[250] br[250] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_251 bl[251] br[251] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_252 bl[252] br[252] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_253 bl[253] br[253] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_254 bl[254] br[254] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_255 bl[255] br[255] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_106_0 bl[0] br[0] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_1 bl[1] br[1] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_2 bl[2] br[2] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_3 bl[3] br[3] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_4 bl[4] br[4] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_5 bl[5] br[5] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_6 bl[6] br[6] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_7 bl[7] br[7] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_8 bl[8] br[8] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_9 bl[9] br[9] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_10 bl[10] br[10] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_11 bl[11] br[11] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_12 bl[12] br[12] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_13 bl[13] br[13] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_14 bl[14] br[14] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_15 bl[15] br[15] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_16 bl[16] br[16] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_17 bl[17] br[17] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_18 bl[18] br[18] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_19 bl[19] br[19] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_20 bl[20] br[20] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_21 bl[21] br[21] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_22 bl[22] br[22] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_23 bl[23] br[23] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_24 bl[24] br[24] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_25 bl[25] br[25] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_26 bl[26] br[26] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_27 bl[27] br[27] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_28 bl[28] br[28] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_29 bl[29] br[29] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_30 bl[30] br[30] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_31 bl[31] br[31] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_32 bl[32] br[32] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_33 bl[33] br[33] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_34 bl[34] br[34] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_35 bl[35] br[35] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_36 bl[36] br[36] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_37 bl[37] br[37] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_38 bl[38] br[38] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_39 bl[39] br[39] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_40 bl[40] br[40] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_41 bl[41] br[41] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_42 bl[42] br[42] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_43 bl[43] br[43] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_44 bl[44] br[44] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_45 bl[45] br[45] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_46 bl[46] br[46] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_47 bl[47] br[47] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_48 bl[48] br[48] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_49 bl[49] br[49] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_50 bl[50] br[50] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_51 bl[51] br[51] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_52 bl[52] br[52] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_53 bl[53] br[53] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_54 bl[54] br[54] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_55 bl[55] br[55] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_56 bl[56] br[56] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_57 bl[57] br[57] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_58 bl[58] br[58] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_59 bl[59] br[59] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_60 bl[60] br[60] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_61 bl[61] br[61] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_62 bl[62] br[62] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_63 bl[63] br[63] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_64 bl[64] br[64] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_65 bl[65] br[65] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_66 bl[66] br[66] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_67 bl[67] br[67] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_68 bl[68] br[68] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_69 bl[69] br[69] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_70 bl[70] br[70] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_71 bl[71] br[71] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_72 bl[72] br[72] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_73 bl[73] br[73] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_74 bl[74] br[74] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_75 bl[75] br[75] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_76 bl[76] br[76] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_77 bl[77] br[77] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_78 bl[78] br[78] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_79 bl[79] br[79] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_80 bl[80] br[80] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_81 bl[81] br[81] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_82 bl[82] br[82] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_83 bl[83] br[83] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_84 bl[84] br[84] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_85 bl[85] br[85] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_86 bl[86] br[86] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_87 bl[87] br[87] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_88 bl[88] br[88] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_89 bl[89] br[89] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_90 bl[90] br[90] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_91 bl[91] br[91] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_92 bl[92] br[92] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_93 bl[93] br[93] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_94 bl[94] br[94] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_95 bl[95] br[95] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_96 bl[96] br[96] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_97 bl[97] br[97] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_98 bl[98] br[98] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_99 bl[99] br[99] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_100 bl[100] br[100] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_101 bl[101] br[101] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_102 bl[102] br[102] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_103 bl[103] br[103] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_104 bl[104] br[104] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_105 bl[105] br[105] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_106 bl[106] br[106] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_107 bl[107] br[107] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_108 bl[108] br[108] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_109 bl[109] br[109] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_110 bl[110] br[110] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_111 bl[111] br[111] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_112 bl[112] br[112] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_113 bl[113] br[113] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_114 bl[114] br[114] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_115 bl[115] br[115] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_116 bl[116] br[116] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_117 bl[117] br[117] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_118 bl[118] br[118] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_119 bl[119] br[119] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_120 bl[120] br[120] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_121 bl[121] br[121] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_122 bl[122] br[122] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_123 bl[123] br[123] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_124 bl[124] br[124] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_125 bl[125] br[125] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_126 bl[126] br[126] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_127 bl[127] br[127] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_128 bl[128] br[128] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_129 bl[129] br[129] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_130 bl[130] br[130] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_131 bl[131] br[131] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_132 bl[132] br[132] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_133 bl[133] br[133] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_134 bl[134] br[134] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_135 bl[135] br[135] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_136 bl[136] br[136] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_137 bl[137] br[137] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_138 bl[138] br[138] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_139 bl[139] br[139] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_140 bl[140] br[140] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_141 bl[141] br[141] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_142 bl[142] br[142] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_143 bl[143] br[143] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_144 bl[144] br[144] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_145 bl[145] br[145] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_146 bl[146] br[146] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_147 bl[147] br[147] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_148 bl[148] br[148] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_149 bl[149] br[149] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_150 bl[150] br[150] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_151 bl[151] br[151] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_152 bl[152] br[152] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_153 bl[153] br[153] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_154 bl[154] br[154] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_155 bl[155] br[155] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_156 bl[156] br[156] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_157 bl[157] br[157] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_158 bl[158] br[158] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_159 bl[159] br[159] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_160 bl[160] br[160] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_161 bl[161] br[161] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_162 bl[162] br[162] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_163 bl[163] br[163] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_164 bl[164] br[164] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_165 bl[165] br[165] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_166 bl[166] br[166] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_167 bl[167] br[167] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_168 bl[168] br[168] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_169 bl[169] br[169] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_170 bl[170] br[170] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_171 bl[171] br[171] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_172 bl[172] br[172] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_173 bl[173] br[173] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_174 bl[174] br[174] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_175 bl[175] br[175] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_176 bl[176] br[176] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_177 bl[177] br[177] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_178 bl[178] br[178] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_179 bl[179] br[179] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_180 bl[180] br[180] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_181 bl[181] br[181] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_182 bl[182] br[182] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_183 bl[183] br[183] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_184 bl[184] br[184] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_185 bl[185] br[185] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_186 bl[186] br[186] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_187 bl[187] br[187] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_188 bl[188] br[188] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_189 bl[189] br[189] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_190 bl[190] br[190] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_191 bl[191] br[191] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_192 bl[192] br[192] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_193 bl[193] br[193] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_194 bl[194] br[194] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_195 bl[195] br[195] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_196 bl[196] br[196] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_197 bl[197] br[197] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_198 bl[198] br[198] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_199 bl[199] br[199] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_200 bl[200] br[200] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_201 bl[201] br[201] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_202 bl[202] br[202] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_203 bl[203] br[203] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_204 bl[204] br[204] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_205 bl[205] br[205] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_206 bl[206] br[206] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_207 bl[207] br[207] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_208 bl[208] br[208] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_209 bl[209] br[209] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_210 bl[210] br[210] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_211 bl[211] br[211] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_212 bl[212] br[212] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_213 bl[213] br[213] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_214 bl[214] br[214] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_215 bl[215] br[215] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_216 bl[216] br[216] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_217 bl[217] br[217] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_218 bl[218] br[218] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_219 bl[219] br[219] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_220 bl[220] br[220] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_221 bl[221] br[221] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_222 bl[222] br[222] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_223 bl[223] br[223] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_224 bl[224] br[224] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_225 bl[225] br[225] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_226 bl[226] br[226] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_227 bl[227] br[227] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_228 bl[228] br[228] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_229 bl[229] br[229] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_230 bl[230] br[230] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_231 bl[231] br[231] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_232 bl[232] br[232] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_233 bl[233] br[233] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_234 bl[234] br[234] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_235 bl[235] br[235] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_236 bl[236] br[236] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_237 bl[237] br[237] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_238 bl[238] br[238] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_239 bl[239] br[239] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_240 bl[240] br[240] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_241 bl[241] br[241] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_242 bl[242] br[242] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_243 bl[243] br[243] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_244 bl[244] br[244] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_245 bl[245] br[245] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_246 bl[246] br[246] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_247 bl[247] br[247] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_248 bl[248] br[248] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_249 bl[249] br[249] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_250 bl[250] br[250] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_251 bl[251] br[251] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_252 bl[252] br[252] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_253 bl[253] br[253] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_254 bl[254] br[254] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_255 bl[255] br[255] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_107_0 bl[0] br[0] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_1 bl[1] br[1] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_2 bl[2] br[2] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_3 bl[3] br[3] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_4 bl[4] br[4] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_5 bl[5] br[5] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_6 bl[6] br[6] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_7 bl[7] br[7] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_8 bl[8] br[8] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_9 bl[9] br[9] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_10 bl[10] br[10] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_11 bl[11] br[11] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_12 bl[12] br[12] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_13 bl[13] br[13] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_14 bl[14] br[14] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_15 bl[15] br[15] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_16 bl[16] br[16] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_17 bl[17] br[17] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_18 bl[18] br[18] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_19 bl[19] br[19] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_20 bl[20] br[20] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_21 bl[21] br[21] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_22 bl[22] br[22] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_23 bl[23] br[23] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_24 bl[24] br[24] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_25 bl[25] br[25] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_26 bl[26] br[26] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_27 bl[27] br[27] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_28 bl[28] br[28] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_29 bl[29] br[29] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_30 bl[30] br[30] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_31 bl[31] br[31] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_32 bl[32] br[32] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_33 bl[33] br[33] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_34 bl[34] br[34] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_35 bl[35] br[35] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_36 bl[36] br[36] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_37 bl[37] br[37] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_38 bl[38] br[38] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_39 bl[39] br[39] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_40 bl[40] br[40] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_41 bl[41] br[41] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_42 bl[42] br[42] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_43 bl[43] br[43] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_44 bl[44] br[44] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_45 bl[45] br[45] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_46 bl[46] br[46] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_47 bl[47] br[47] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_48 bl[48] br[48] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_49 bl[49] br[49] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_50 bl[50] br[50] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_51 bl[51] br[51] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_52 bl[52] br[52] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_53 bl[53] br[53] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_54 bl[54] br[54] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_55 bl[55] br[55] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_56 bl[56] br[56] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_57 bl[57] br[57] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_58 bl[58] br[58] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_59 bl[59] br[59] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_60 bl[60] br[60] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_61 bl[61] br[61] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_62 bl[62] br[62] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_63 bl[63] br[63] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_64 bl[64] br[64] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_65 bl[65] br[65] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_66 bl[66] br[66] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_67 bl[67] br[67] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_68 bl[68] br[68] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_69 bl[69] br[69] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_70 bl[70] br[70] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_71 bl[71] br[71] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_72 bl[72] br[72] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_73 bl[73] br[73] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_74 bl[74] br[74] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_75 bl[75] br[75] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_76 bl[76] br[76] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_77 bl[77] br[77] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_78 bl[78] br[78] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_79 bl[79] br[79] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_80 bl[80] br[80] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_81 bl[81] br[81] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_82 bl[82] br[82] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_83 bl[83] br[83] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_84 bl[84] br[84] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_85 bl[85] br[85] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_86 bl[86] br[86] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_87 bl[87] br[87] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_88 bl[88] br[88] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_89 bl[89] br[89] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_90 bl[90] br[90] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_91 bl[91] br[91] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_92 bl[92] br[92] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_93 bl[93] br[93] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_94 bl[94] br[94] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_95 bl[95] br[95] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_96 bl[96] br[96] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_97 bl[97] br[97] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_98 bl[98] br[98] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_99 bl[99] br[99] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_100 bl[100] br[100] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_101 bl[101] br[101] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_102 bl[102] br[102] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_103 bl[103] br[103] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_104 bl[104] br[104] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_105 bl[105] br[105] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_106 bl[106] br[106] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_107 bl[107] br[107] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_108 bl[108] br[108] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_109 bl[109] br[109] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_110 bl[110] br[110] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_111 bl[111] br[111] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_112 bl[112] br[112] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_113 bl[113] br[113] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_114 bl[114] br[114] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_115 bl[115] br[115] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_116 bl[116] br[116] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_117 bl[117] br[117] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_118 bl[118] br[118] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_119 bl[119] br[119] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_120 bl[120] br[120] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_121 bl[121] br[121] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_122 bl[122] br[122] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_123 bl[123] br[123] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_124 bl[124] br[124] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_125 bl[125] br[125] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_126 bl[126] br[126] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_127 bl[127] br[127] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_128 bl[128] br[128] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_129 bl[129] br[129] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_130 bl[130] br[130] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_131 bl[131] br[131] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_132 bl[132] br[132] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_133 bl[133] br[133] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_134 bl[134] br[134] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_135 bl[135] br[135] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_136 bl[136] br[136] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_137 bl[137] br[137] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_138 bl[138] br[138] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_139 bl[139] br[139] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_140 bl[140] br[140] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_141 bl[141] br[141] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_142 bl[142] br[142] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_143 bl[143] br[143] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_144 bl[144] br[144] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_145 bl[145] br[145] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_146 bl[146] br[146] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_147 bl[147] br[147] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_148 bl[148] br[148] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_149 bl[149] br[149] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_150 bl[150] br[150] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_151 bl[151] br[151] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_152 bl[152] br[152] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_153 bl[153] br[153] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_154 bl[154] br[154] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_155 bl[155] br[155] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_156 bl[156] br[156] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_157 bl[157] br[157] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_158 bl[158] br[158] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_159 bl[159] br[159] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_160 bl[160] br[160] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_161 bl[161] br[161] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_162 bl[162] br[162] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_163 bl[163] br[163] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_164 bl[164] br[164] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_165 bl[165] br[165] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_166 bl[166] br[166] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_167 bl[167] br[167] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_168 bl[168] br[168] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_169 bl[169] br[169] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_170 bl[170] br[170] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_171 bl[171] br[171] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_172 bl[172] br[172] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_173 bl[173] br[173] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_174 bl[174] br[174] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_175 bl[175] br[175] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_176 bl[176] br[176] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_177 bl[177] br[177] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_178 bl[178] br[178] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_179 bl[179] br[179] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_180 bl[180] br[180] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_181 bl[181] br[181] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_182 bl[182] br[182] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_183 bl[183] br[183] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_184 bl[184] br[184] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_185 bl[185] br[185] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_186 bl[186] br[186] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_187 bl[187] br[187] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_188 bl[188] br[188] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_189 bl[189] br[189] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_190 bl[190] br[190] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_191 bl[191] br[191] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_192 bl[192] br[192] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_193 bl[193] br[193] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_194 bl[194] br[194] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_195 bl[195] br[195] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_196 bl[196] br[196] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_197 bl[197] br[197] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_198 bl[198] br[198] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_199 bl[199] br[199] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_200 bl[200] br[200] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_201 bl[201] br[201] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_202 bl[202] br[202] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_203 bl[203] br[203] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_204 bl[204] br[204] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_205 bl[205] br[205] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_206 bl[206] br[206] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_207 bl[207] br[207] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_208 bl[208] br[208] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_209 bl[209] br[209] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_210 bl[210] br[210] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_211 bl[211] br[211] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_212 bl[212] br[212] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_213 bl[213] br[213] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_214 bl[214] br[214] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_215 bl[215] br[215] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_216 bl[216] br[216] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_217 bl[217] br[217] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_218 bl[218] br[218] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_219 bl[219] br[219] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_220 bl[220] br[220] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_221 bl[221] br[221] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_222 bl[222] br[222] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_223 bl[223] br[223] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_224 bl[224] br[224] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_225 bl[225] br[225] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_226 bl[226] br[226] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_227 bl[227] br[227] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_228 bl[228] br[228] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_229 bl[229] br[229] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_230 bl[230] br[230] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_231 bl[231] br[231] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_232 bl[232] br[232] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_233 bl[233] br[233] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_234 bl[234] br[234] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_235 bl[235] br[235] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_236 bl[236] br[236] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_237 bl[237] br[237] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_238 bl[238] br[238] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_239 bl[239] br[239] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_240 bl[240] br[240] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_241 bl[241] br[241] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_242 bl[242] br[242] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_243 bl[243] br[243] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_244 bl[244] br[244] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_245 bl[245] br[245] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_246 bl[246] br[246] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_247 bl[247] br[247] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_248 bl[248] br[248] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_249 bl[249] br[249] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_250 bl[250] br[250] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_251 bl[251] br[251] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_252 bl[252] br[252] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_253 bl[253] br[253] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_254 bl[254] br[254] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_255 bl[255] br[255] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_108_0 bl[0] br[0] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_1 bl[1] br[1] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_2 bl[2] br[2] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_3 bl[3] br[3] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_4 bl[4] br[4] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_5 bl[5] br[5] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_6 bl[6] br[6] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_7 bl[7] br[7] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_8 bl[8] br[8] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_9 bl[9] br[9] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_10 bl[10] br[10] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_11 bl[11] br[11] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_12 bl[12] br[12] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_13 bl[13] br[13] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_14 bl[14] br[14] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_15 bl[15] br[15] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_16 bl[16] br[16] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_17 bl[17] br[17] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_18 bl[18] br[18] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_19 bl[19] br[19] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_20 bl[20] br[20] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_21 bl[21] br[21] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_22 bl[22] br[22] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_23 bl[23] br[23] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_24 bl[24] br[24] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_25 bl[25] br[25] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_26 bl[26] br[26] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_27 bl[27] br[27] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_28 bl[28] br[28] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_29 bl[29] br[29] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_30 bl[30] br[30] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_31 bl[31] br[31] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_32 bl[32] br[32] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_33 bl[33] br[33] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_34 bl[34] br[34] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_35 bl[35] br[35] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_36 bl[36] br[36] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_37 bl[37] br[37] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_38 bl[38] br[38] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_39 bl[39] br[39] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_40 bl[40] br[40] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_41 bl[41] br[41] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_42 bl[42] br[42] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_43 bl[43] br[43] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_44 bl[44] br[44] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_45 bl[45] br[45] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_46 bl[46] br[46] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_47 bl[47] br[47] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_48 bl[48] br[48] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_49 bl[49] br[49] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_50 bl[50] br[50] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_51 bl[51] br[51] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_52 bl[52] br[52] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_53 bl[53] br[53] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_54 bl[54] br[54] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_55 bl[55] br[55] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_56 bl[56] br[56] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_57 bl[57] br[57] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_58 bl[58] br[58] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_59 bl[59] br[59] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_60 bl[60] br[60] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_61 bl[61] br[61] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_62 bl[62] br[62] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_63 bl[63] br[63] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_64 bl[64] br[64] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_65 bl[65] br[65] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_66 bl[66] br[66] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_67 bl[67] br[67] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_68 bl[68] br[68] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_69 bl[69] br[69] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_70 bl[70] br[70] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_71 bl[71] br[71] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_72 bl[72] br[72] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_73 bl[73] br[73] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_74 bl[74] br[74] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_75 bl[75] br[75] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_76 bl[76] br[76] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_77 bl[77] br[77] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_78 bl[78] br[78] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_79 bl[79] br[79] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_80 bl[80] br[80] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_81 bl[81] br[81] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_82 bl[82] br[82] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_83 bl[83] br[83] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_84 bl[84] br[84] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_85 bl[85] br[85] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_86 bl[86] br[86] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_87 bl[87] br[87] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_88 bl[88] br[88] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_89 bl[89] br[89] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_90 bl[90] br[90] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_91 bl[91] br[91] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_92 bl[92] br[92] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_93 bl[93] br[93] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_94 bl[94] br[94] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_95 bl[95] br[95] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_96 bl[96] br[96] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_97 bl[97] br[97] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_98 bl[98] br[98] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_99 bl[99] br[99] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_100 bl[100] br[100] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_101 bl[101] br[101] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_102 bl[102] br[102] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_103 bl[103] br[103] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_104 bl[104] br[104] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_105 bl[105] br[105] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_106 bl[106] br[106] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_107 bl[107] br[107] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_108 bl[108] br[108] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_109 bl[109] br[109] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_110 bl[110] br[110] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_111 bl[111] br[111] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_112 bl[112] br[112] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_113 bl[113] br[113] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_114 bl[114] br[114] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_115 bl[115] br[115] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_116 bl[116] br[116] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_117 bl[117] br[117] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_118 bl[118] br[118] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_119 bl[119] br[119] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_120 bl[120] br[120] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_121 bl[121] br[121] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_122 bl[122] br[122] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_123 bl[123] br[123] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_124 bl[124] br[124] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_125 bl[125] br[125] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_126 bl[126] br[126] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_127 bl[127] br[127] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_128 bl[128] br[128] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_129 bl[129] br[129] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_130 bl[130] br[130] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_131 bl[131] br[131] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_132 bl[132] br[132] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_133 bl[133] br[133] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_134 bl[134] br[134] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_135 bl[135] br[135] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_136 bl[136] br[136] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_137 bl[137] br[137] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_138 bl[138] br[138] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_139 bl[139] br[139] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_140 bl[140] br[140] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_141 bl[141] br[141] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_142 bl[142] br[142] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_143 bl[143] br[143] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_144 bl[144] br[144] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_145 bl[145] br[145] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_146 bl[146] br[146] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_147 bl[147] br[147] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_148 bl[148] br[148] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_149 bl[149] br[149] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_150 bl[150] br[150] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_151 bl[151] br[151] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_152 bl[152] br[152] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_153 bl[153] br[153] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_154 bl[154] br[154] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_155 bl[155] br[155] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_156 bl[156] br[156] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_157 bl[157] br[157] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_158 bl[158] br[158] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_159 bl[159] br[159] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_160 bl[160] br[160] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_161 bl[161] br[161] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_162 bl[162] br[162] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_163 bl[163] br[163] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_164 bl[164] br[164] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_165 bl[165] br[165] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_166 bl[166] br[166] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_167 bl[167] br[167] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_168 bl[168] br[168] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_169 bl[169] br[169] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_170 bl[170] br[170] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_171 bl[171] br[171] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_172 bl[172] br[172] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_173 bl[173] br[173] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_174 bl[174] br[174] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_175 bl[175] br[175] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_176 bl[176] br[176] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_177 bl[177] br[177] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_178 bl[178] br[178] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_179 bl[179] br[179] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_180 bl[180] br[180] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_181 bl[181] br[181] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_182 bl[182] br[182] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_183 bl[183] br[183] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_184 bl[184] br[184] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_185 bl[185] br[185] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_186 bl[186] br[186] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_187 bl[187] br[187] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_188 bl[188] br[188] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_189 bl[189] br[189] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_190 bl[190] br[190] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_191 bl[191] br[191] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_192 bl[192] br[192] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_193 bl[193] br[193] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_194 bl[194] br[194] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_195 bl[195] br[195] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_196 bl[196] br[196] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_197 bl[197] br[197] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_198 bl[198] br[198] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_199 bl[199] br[199] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_200 bl[200] br[200] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_201 bl[201] br[201] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_202 bl[202] br[202] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_203 bl[203] br[203] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_204 bl[204] br[204] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_205 bl[205] br[205] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_206 bl[206] br[206] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_207 bl[207] br[207] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_208 bl[208] br[208] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_209 bl[209] br[209] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_210 bl[210] br[210] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_211 bl[211] br[211] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_212 bl[212] br[212] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_213 bl[213] br[213] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_214 bl[214] br[214] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_215 bl[215] br[215] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_216 bl[216] br[216] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_217 bl[217] br[217] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_218 bl[218] br[218] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_219 bl[219] br[219] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_220 bl[220] br[220] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_221 bl[221] br[221] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_222 bl[222] br[222] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_223 bl[223] br[223] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_224 bl[224] br[224] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_225 bl[225] br[225] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_226 bl[226] br[226] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_227 bl[227] br[227] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_228 bl[228] br[228] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_229 bl[229] br[229] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_230 bl[230] br[230] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_231 bl[231] br[231] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_232 bl[232] br[232] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_233 bl[233] br[233] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_234 bl[234] br[234] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_235 bl[235] br[235] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_236 bl[236] br[236] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_237 bl[237] br[237] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_238 bl[238] br[238] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_239 bl[239] br[239] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_240 bl[240] br[240] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_241 bl[241] br[241] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_242 bl[242] br[242] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_243 bl[243] br[243] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_244 bl[244] br[244] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_245 bl[245] br[245] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_246 bl[246] br[246] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_247 bl[247] br[247] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_248 bl[248] br[248] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_249 bl[249] br[249] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_250 bl[250] br[250] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_251 bl[251] br[251] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_252 bl[252] br[252] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_253 bl[253] br[253] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_254 bl[254] br[254] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_255 bl[255] br[255] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_109_0 bl[0] br[0] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_1 bl[1] br[1] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_2 bl[2] br[2] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_3 bl[3] br[3] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_4 bl[4] br[4] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_5 bl[5] br[5] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_6 bl[6] br[6] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_7 bl[7] br[7] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_8 bl[8] br[8] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_9 bl[9] br[9] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_10 bl[10] br[10] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_11 bl[11] br[11] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_12 bl[12] br[12] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_13 bl[13] br[13] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_14 bl[14] br[14] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_15 bl[15] br[15] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_16 bl[16] br[16] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_17 bl[17] br[17] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_18 bl[18] br[18] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_19 bl[19] br[19] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_20 bl[20] br[20] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_21 bl[21] br[21] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_22 bl[22] br[22] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_23 bl[23] br[23] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_24 bl[24] br[24] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_25 bl[25] br[25] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_26 bl[26] br[26] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_27 bl[27] br[27] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_28 bl[28] br[28] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_29 bl[29] br[29] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_30 bl[30] br[30] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_31 bl[31] br[31] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_32 bl[32] br[32] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_33 bl[33] br[33] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_34 bl[34] br[34] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_35 bl[35] br[35] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_36 bl[36] br[36] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_37 bl[37] br[37] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_38 bl[38] br[38] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_39 bl[39] br[39] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_40 bl[40] br[40] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_41 bl[41] br[41] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_42 bl[42] br[42] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_43 bl[43] br[43] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_44 bl[44] br[44] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_45 bl[45] br[45] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_46 bl[46] br[46] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_47 bl[47] br[47] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_48 bl[48] br[48] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_49 bl[49] br[49] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_50 bl[50] br[50] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_51 bl[51] br[51] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_52 bl[52] br[52] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_53 bl[53] br[53] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_54 bl[54] br[54] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_55 bl[55] br[55] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_56 bl[56] br[56] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_57 bl[57] br[57] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_58 bl[58] br[58] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_59 bl[59] br[59] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_60 bl[60] br[60] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_61 bl[61] br[61] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_62 bl[62] br[62] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_63 bl[63] br[63] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_64 bl[64] br[64] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_65 bl[65] br[65] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_66 bl[66] br[66] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_67 bl[67] br[67] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_68 bl[68] br[68] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_69 bl[69] br[69] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_70 bl[70] br[70] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_71 bl[71] br[71] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_72 bl[72] br[72] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_73 bl[73] br[73] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_74 bl[74] br[74] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_75 bl[75] br[75] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_76 bl[76] br[76] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_77 bl[77] br[77] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_78 bl[78] br[78] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_79 bl[79] br[79] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_80 bl[80] br[80] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_81 bl[81] br[81] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_82 bl[82] br[82] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_83 bl[83] br[83] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_84 bl[84] br[84] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_85 bl[85] br[85] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_86 bl[86] br[86] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_87 bl[87] br[87] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_88 bl[88] br[88] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_89 bl[89] br[89] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_90 bl[90] br[90] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_91 bl[91] br[91] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_92 bl[92] br[92] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_93 bl[93] br[93] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_94 bl[94] br[94] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_95 bl[95] br[95] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_96 bl[96] br[96] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_97 bl[97] br[97] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_98 bl[98] br[98] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_99 bl[99] br[99] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_100 bl[100] br[100] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_101 bl[101] br[101] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_102 bl[102] br[102] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_103 bl[103] br[103] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_104 bl[104] br[104] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_105 bl[105] br[105] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_106 bl[106] br[106] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_107 bl[107] br[107] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_108 bl[108] br[108] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_109 bl[109] br[109] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_110 bl[110] br[110] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_111 bl[111] br[111] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_112 bl[112] br[112] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_113 bl[113] br[113] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_114 bl[114] br[114] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_115 bl[115] br[115] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_116 bl[116] br[116] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_117 bl[117] br[117] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_118 bl[118] br[118] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_119 bl[119] br[119] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_120 bl[120] br[120] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_121 bl[121] br[121] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_122 bl[122] br[122] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_123 bl[123] br[123] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_124 bl[124] br[124] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_125 bl[125] br[125] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_126 bl[126] br[126] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_127 bl[127] br[127] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_128 bl[128] br[128] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_129 bl[129] br[129] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_130 bl[130] br[130] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_131 bl[131] br[131] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_132 bl[132] br[132] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_133 bl[133] br[133] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_134 bl[134] br[134] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_135 bl[135] br[135] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_136 bl[136] br[136] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_137 bl[137] br[137] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_138 bl[138] br[138] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_139 bl[139] br[139] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_140 bl[140] br[140] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_141 bl[141] br[141] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_142 bl[142] br[142] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_143 bl[143] br[143] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_144 bl[144] br[144] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_145 bl[145] br[145] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_146 bl[146] br[146] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_147 bl[147] br[147] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_148 bl[148] br[148] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_149 bl[149] br[149] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_150 bl[150] br[150] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_151 bl[151] br[151] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_152 bl[152] br[152] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_153 bl[153] br[153] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_154 bl[154] br[154] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_155 bl[155] br[155] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_156 bl[156] br[156] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_157 bl[157] br[157] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_158 bl[158] br[158] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_159 bl[159] br[159] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_160 bl[160] br[160] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_161 bl[161] br[161] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_162 bl[162] br[162] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_163 bl[163] br[163] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_164 bl[164] br[164] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_165 bl[165] br[165] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_166 bl[166] br[166] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_167 bl[167] br[167] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_168 bl[168] br[168] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_169 bl[169] br[169] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_170 bl[170] br[170] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_171 bl[171] br[171] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_172 bl[172] br[172] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_173 bl[173] br[173] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_174 bl[174] br[174] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_175 bl[175] br[175] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_176 bl[176] br[176] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_177 bl[177] br[177] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_178 bl[178] br[178] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_179 bl[179] br[179] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_180 bl[180] br[180] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_181 bl[181] br[181] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_182 bl[182] br[182] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_183 bl[183] br[183] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_184 bl[184] br[184] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_185 bl[185] br[185] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_186 bl[186] br[186] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_187 bl[187] br[187] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_188 bl[188] br[188] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_189 bl[189] br[189] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_190 bl[190] br[190] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_191 bl[191] br[191] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_192 bl[192] br[192] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_193 bl[193] br[193] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_194 bl[194] br[194] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_195 bl[195] br[195] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_196 bl[196] br[196] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_197 bl[197] br[197] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_198 bl[198] br[198] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_199 bl[199] br[199] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_200 bl[200] br[200] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_201 bl[201] br[201] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_202 bl[202] br[202] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_203 bl[203] br[203] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_204 bl[204] br[204] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_205 bl[205] br[205] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_206 bl[206] br[206] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_207 bl[207] br[207] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_208 bl[208] br[208] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_209 bl[209] br[209] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_210 bl[210] br[210] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_211 bl[211] br[211] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_212 bl[212] br[212] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_213 bl[213] br[213] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_214 bl[214] br[214] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_215 bl[215] br[215] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_216 bl[216] br[216] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_217 bl[217] br[217] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_218 bl[218] br[218] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_219 bl[219] br[219] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_220 bl[220] br[220] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_221 bl[221] br[221] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_222 bl[222] br[222] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_223 bl[223] br[223] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_224 bl[224] br[224] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_225 bl[225] br[225] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_226 bl[226] br[226] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_227 bl[227] br[227] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_228 bl[228] br[228] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_229 bl[229] br[229] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_230 bl[230] br[230] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_231 bl[231] br[231] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_232 bl[232] br[232] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_233 bl[233] br[233] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_234 bl[234] br[234] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_235 bl[235] br[235] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_236 bl[236] br[236] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_237 bl[237] br[237] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_238 bl[238] br[238] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_239 bl[239] br[239] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_240 bl[240] br[240] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_241 bl[241] br[241] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_242 bl[242] br[242] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_243 bl[243] br[243] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_244 bl[244] br[244] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_245 bl[245] br[245] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_246 bl[246] br[246] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_247 bl[247] br[247] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_248 bl[248] br[248] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_249 bl[249] br[249] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_250 bl[250] br[250] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_251 bl[251] br[251] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_252 bl[252] br[252] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_253 bl[253] br[253] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_254 bl[254] br[254] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_255 bl[255] br[255] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_110_0 bl[0] br[0] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_1 bl[1] br[1] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_2 bl[2] br[2] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_3 bl[3] br[3] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_4 bl[4] br[4] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_5 bl[5] br[5] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_6 bl[6] br[6] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_7 bl[7] br[7] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_8 bl[8] br[8] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_9 bl[9] br[9] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_10 bl[10] br[10] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_11 bl[11] br[11] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_12 bl[12] br[12] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_13 bl[13] br[13] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_14 bl[14] br[14] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_15 bl[15] br[15] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_16 bl[16] br[16] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_17 bl[17] br[17] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_18 bl[18] br[18] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_19 bl[19] br[19] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_20 bl[20] br[20] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_21 bl[21] br[21] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_22 bl[22] br[22] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_23 bl[23] br[23] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_24 bl[24] br[24] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_25 bl[25] br[25] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_26 bl[26] br[26] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_27 bl[27] br[27] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_28 bl[28] br[28] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_29 bl[29] br[29] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_30 bl[30] br[30] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_31 bl[31] br[31] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_32 bl[32] br[32] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_33 bl[33] br[33] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_34 bl[34] br[34] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_35 bl[35] br[35] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_36 bl[36] br[36] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_37 bl[37] br[37] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_38 bl[38] br[38] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_39 bl[39] br[39] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_40 bl[40] br[40] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_41 bl[41] br[41] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_42 bl[42] br[42] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_43 bl[43] br[43] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_44 bl[44] br[44] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_45 bl[45] br[45] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_46 bl[46] br[46] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_47 bl[47] br[47] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_48 bl[48] br[48] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_49 bl[49] br[49] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_50 bl[50] br[50] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_51 bl[51] br[51] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_52 bl[52] br[52] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_53 bl[53] br[53] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_54 bl[54] br[54] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_55 bl[55] br[55] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_56 bl[56] br[56] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_57 bl[57] br[57] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_58 bl[58] br[58] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_59 bl[59] br[59] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_60 bl[60] br[60] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_61 bl[61] br[61] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_62 bl[62] br[62] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_63 bl[63] br[63] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_64 bl[64] br[64] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_65 bl[65] br[65] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_66 bl[66] br[66] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_67 bl[67] br[67] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_68 bl[68] br[68] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_69 bl[69] br[69] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_70 bl[70] br[70] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_71 bl[71] br[71] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_72 bl[72] br[72] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_73 bl[73] br[73] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_74 bl[74] br[74] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_75 bl[75] br[75] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_76 bl[76] br[76] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_77 bl[77] br[77] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_78 bl[78] br[78] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_79 bl[79] br[79] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_80 bl[80] br[80] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_81 bl[81] br[81] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_82 bl[82] br[82] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_83 bl[83] br[83] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_84 bl[84] br[84] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_85 bl[85] br[85] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_86 bl[86] br[86] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_87 bl[87] br[87] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_88 bl[88] br[88] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_89 bl[89] br[89] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_90 bl[90] br[90] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_91 bl[91] br[91] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_92 bl[92] br[92] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_93 bl[93] br[93] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_94 bl[94] br[94] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_95 bl[95] br[95] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_96 bl[96] br[96] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_97 bl[97] br[97] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_98 bl[98] br[98] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_99 bl[99] br[99] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_100 bl[100] br[100] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_101 bl[101] br[101] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_102 bl[102] br[102] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_103 bl[103] br[103] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_104 bl[104] br[104] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_105 bl[105] br[105] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_106 bl[106] br[106] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_107 bl[107] br[107] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_108 bl[108] br[108] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_109 bl[109] br[109] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_110 bl[110] br[110] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_111 bl[111] br[111] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_112 bl[112] br[112] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_113 bl[113] br[113] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_114 bl[114] br[114] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_115 bl[115] br[115] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_116 bl[116] br[116] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_117 bl[117] br[117] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_118 bl[118] br[118] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_119 bl[119] br[119] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_120 bl[120] br[120] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_121 bl[121] br[121] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_122 bl[122] br[122] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_123 bl[123] br[123] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_124 bl[124] br[124] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_125 bl[125] br[125] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_126 bl[126] br[126] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_127 bl[127] br[127] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_128 bl[128] br[128] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_129 bl[129] br[129] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_130 bl[130] br[130] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_131 bl[131] br[131] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_132 bl[132] br[132] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_133 bl[133] br[133] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_134 bl[134] br[134] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_135 bl[135] br[135] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_136 bl[136] br[136] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_137 bl[137] br[137] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_138 bl[138] br[138] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_139 bl[139] br[139] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_140 bl[140] br[140] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_141 bl[141] br[141] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_142 bl[142] br[142] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_143 bl[143] br[143] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_144 bl[144] br[144] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_145 bl[145] br[145] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_146 bl[146] br[146] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_147 bl[147] br[147] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_148 bl[148] br[148] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_149 bl[149] br[149] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_150 bl[150] br[150] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_151 bl[151] br[151] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_152 bl[152] br[152] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_153 bl[153] br[153] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_154 bl[154] br[154] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_155 bl[155] br[155] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_156 bl[156] br[156] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_157 bl[157] br[157] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_158 bl[158] br[158] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_159 bl[159] br[159] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_160 bl[160] br[160] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_161 bl[161] br[161] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_162 bl[162] br[162] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_163 bl[163] br[163] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_164 bl[164] br[164] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_165 bl[165] br[165] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_166 bl[166] br[166] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_167 bl[167] br[167] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_168 bl[168] br[168] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_169 bl[169] br[169] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_170 bl[170] br[170] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_171 bl[171] br[171] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_172 bl[172] br[172] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_173 bl[173] br[173] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_174 bl[174] br[174] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_175 bl[175] br[175] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_176 bl[176] br[176] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_177 bl[177] br[177] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_178 bl[178] br[178] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_179 bl[179] br[179] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_180 bl[180] br[180] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_181 bl[181] br[181] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_182 bl[182] br[182] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_183 bl[183] br[183] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_184 bl[184] br[184] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_185 bl[185] br[185] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_186 bl[186] br[186] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_187 bl[187] br[187] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_188 bl[188] br[188] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_189 bl[189] br[189] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_190 bl[190] br[190] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_191 bl[191] br[191] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_192 bl[192] br[192] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_193 bl[193] br[193] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_194 bl[194] br[194] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_195 bl[195] br[195] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_196 bl[196] br[196] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_197 bl[197] br[197] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_198 bl[198] br[198] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_199 bl[199] br[199] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_200 bl[200] br[200] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_201 bl[201] br[201] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_202 bl[202] br[202] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_203 bl[203] br[203] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_204 bl[204] br[204] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_205 bl[205] br[205] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_206 bl[206] br[206] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_207 bl[207] br[207] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_208 bl[208] br[208] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_209 bl[209] br[209] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_210 bl[210] br[210] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_211 bl[211] br[211] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_212 bl[212] br[212] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_213 bl[213] br[213] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_214 bl[214] br[214] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_215 bl[215] br[215] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_216 bl[216] br[216] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_217 bl[217] br[217] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_218 bl[218] br[218] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_219 bl[219] br[219] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_220 bl[220] br[220] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_221 bl[221] br[221] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_222 bl[222] br[222] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_223 bl[223] br[223] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_224 bl[224] br[224] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_225 bl[225] br[225] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_226 bl[226] br[226] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_227 bl[227] br[227] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_228 bl[228] br[228] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_229 bl[229] br[229] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_230 bl[230] br[230] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_231 bl[231] br[231] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_232 bl[232] br[232] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_233 bl[233] br[233] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_234 bl[234] br[234] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_235 bl[235] br[235] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_236 bl[236] br[236] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_237 bl[237] br[237] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_238 bl[238] br[238] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_239 bl[239] br[239] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_240 bl[240] br[240] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_241 bl[241] br[241] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_242 bl[242] br[242] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_243 bl[243] br[243] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_244 bl[244] br[244] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_245 bl[245] br[245] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_246 bl[246] br[246] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_247 bl[247] br[247] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_248 bl[248] br[248] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_249 bl[249] br[249] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_250 bl[250] br[250] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_251 bl[251] br[251] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_252 bl[252] br[252] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_253 bl[253] br[253] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_254 bl[254] br[254] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_255 bl[255] br[255] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_111_0 bl[0] br[0] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_1 bl[1] br[1] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_2 bl[2] br[2] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_3 bl[3] br[3] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_4 bl[4] br[4] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_5 bl[5] br[5] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_6 bl[6] br[6] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_7 bl[7] br[7] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_8 bl[8] br[8] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_9 bl[9] br[9] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_10 bl[10] br[10] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_11 bl[11] br[11] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_12 bl[12] br[12] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_13 bl[13] br[13] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_14 bl[14] br[14] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_15 bl[15] br[15] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_16 bl[16] br[16] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_17 bl[17] br[17] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_18 bl[18] br[18] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_19 bl[19] br[19] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_20 bl[20] br[20] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_21 bl[21] br[21] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_22 bl[22] br[22] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_23 bl[23] br[23] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_24 bl[24] br[24] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_25 bl[25] br[25] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_26 bl[26] br[26] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_27 bl[27] br[27] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_28 bl[28] br[28] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_29 bl[29] br[29] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_30 bl[30] br[30] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_31 bl[31] br[31] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_32 bl[32] br[32] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_33 bl[33] br[33] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_34 bl[34] br[34] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_35 bl[35] br[35] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_36 bl[36] br[36] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_37 bl[37] br[37] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_38 bl[38] br[38] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_39 bl[39] br[39] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_40 bl[40] br[40] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_41 bl[41] br[41] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_42 bl[42] br[42] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_43 bl[43] br[43] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_44 bl[44] br[44] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_45 bl[45] br[45] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_46 bl[46] br[46] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_47 bl[47] br[47] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_48 bl[48] br[48] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_49 bl[49] br[49] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_50 bl[50] br[50] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_51 bl[51] br[51] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_52 bl[52] br[52] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_53 bl[53] br[53] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_54 bl[54] br[54] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_55 bl[55] br[55] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_56 bl[56] br[56] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_57 bl[57] br[57] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_58 bl[58] br[58] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_59 bl[59] br[59] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_60 bl[60] br[60] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_61 bl[61] br[61] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_62 bl[62] br[62] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_63 bl[63] br[63] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_64 bl[64] br[64] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_65 bl[65] br[65] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_66 bl[66] br[66] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_67 bl[67] br[67] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_68 bl[68] br[68] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_69 bl[69] br[69] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_70 bl[70] br[70] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_71 bl[71] br[71] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_72 bl[72] br[72] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_73 bl[73] br[73] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_74 bl[74] br[74] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_75 bl[75] br[75] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_76 bl[76] br[76] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_77 bl[77] br[77] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_78 bl[78] br[78] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_79 bl[79] br[79] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_80 bl[80] br[80] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_81 bl[81] br[81] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_82 bl[82] br[82] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_83 bl[83] br[83] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_84 bl[84] br[84] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_85 bl[85] br[85] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_86 bl[86] br[86] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_87 bl[87] br[87] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_88 bl[88] br[88] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_89 bl[89] br[89] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_90 bl[90] br[90] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_91 bl[91] br[91] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_92 bl[92] br[92] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_93 bl[93] br[93] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_94 bl[94] br[94] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_95 bl[95] br[95] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_96 bl[96] br[96] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_97 bl[97] br[97] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_98 bl[98] br[98] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_99 bl[99] br[99] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_100 bl[100] br[100] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_101 bl[101] br[101] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_102 bl[102] br[102] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_103 bl[103] br[103] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_104 bl[104] br[104] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_105 bl[105] br[105] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_106 bl[106] br[106] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_107 bl[107] br[107] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_108 bl[108] br[108] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_109 bl[109] br[109] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_110 bl[110] br[110] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_111 bl[111] br[111] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_112 bl[112] br[112] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_113 bl[113] br[113] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_114 bl[114] br[114] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_115 bl[115] br[115] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_116 bl[116] br[116] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_117 bl[117] br[117] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_118 bl[118] br[118] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_119 bl[119] br[119] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_120 bl[120] br[120] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_121 bl[121] br[121] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_122 bl[122] br[122] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_123 bl[123] br[123] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_124 bl[124] br[124] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_125 bl[125] br[125] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_126 bl[126] br[126] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_127 bl[127] br[127] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_128 bl[128] br[128] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_129 bl[129] br[129] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_130 bl[130] br[130] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_131 bl[131] br[131] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_132 bl[132] br[132] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_133 bl[133] br[133] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_134 bl[134] br[134] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_135 bl[135] br[135] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_136 bl[136] br[136] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_137 bl[137] br[137] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_138 bl[138] br[138] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_139 bl[139] br[139] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_140 bl[140] br[140] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_141 bl[141] br[141] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_142 bl[142] br[142] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_143 bl[143] br[143] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_144 bl[144] br[144] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_145 bl[145] br[145] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_146 bl[146] br[146] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_147 bl[147] br[147] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_148 bl[148] br[148] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_149 bl[149] br[149] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_150 bl[150] br[150] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_151 bl[151] br[151] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_152 bl[152] br[152] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_153 bl[153] br[153] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_154 bl[154] br[154] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_155 bl[155] br[155] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_156 bl[156] br[156] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_157 bl[157] br[157] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_158 bl[158] br[158] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_159 bl[159] br[159] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_160 bl[160] br[160] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_161 bl[161] br[161] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_162 bl[162] br[162] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_163 bl[163] br[163] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_164 bl[164] br[164] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_165 bl[165] br[165] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_166 bl[166] br[166] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_167 bl[167] br[167] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_168 bl[168] br[168] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_169 bl[169] br[169] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_170 bl[170] br[170] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_171 bl[171] br[171] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_172 bl[172] br[172] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_173 bl[173] br[173] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_174 bl[174] br[174] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_175 bl[175] br[175] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_176 bl[176] br[176] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_177 bl[177] br[177] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_178 bl[178] br[178] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_179 bl[179] br[179] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_180 bl[180] br[180] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_181 bl[181] br[181] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_182 bl[182] br[182] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_183 bl[183] br[183] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_184 bl[184] br[184] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_185 bl[185] br[185] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_186 bl[186] br[186] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_187 bl[187] br[187] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_188 bl[188] br[188] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_189 bl[189] br[189] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_190 bl[190] br[190] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_191 bl[191] br[191] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_192 bl[192] br[192] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_193 bl[193] br[193] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_194 bl[194] br[194] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_195 bl[195] br[195] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_196 bl[196] br[196] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_197 bl[197] br[197] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_198 bl[198] br[198] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_199 bl[199] br[199] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_200 bl[200] br[200] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_201 bl[201] br[201] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_202 bl[202] br[202] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_203 bl[203] br[203] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_204 bl[204] br[204] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_205 bl[205] br[205] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_206 bl[206] br[206] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_207 bl[207] br[207] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_208 bl[208] br[208] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_209 bl[209] br[209] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_210 bl[210] br[210] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_211 bl[211] br[211] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_212 bl[212] br[212] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_213 bl[213] br[213] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_214 bl[214] br[214] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_215 bl[215] br[215] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_216 bl[216] br[216] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_217 bl[217] br[217] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_218 bl[218] br[218] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_219 bl[219] br[219] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_220 bl[220] br[220] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_221 bl[221] br[221] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_222 bl[222] br[222] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_223 bl[223] br[223] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_224 bl[224] br[224] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_225 bl[225] br[225] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_226 bl[226] br[226] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_227 bl[227] br[227] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_228 bl[228] br[228] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_229 bl[229] br[229] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_230 bl[230] br[230] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_231 bl[231] br[231] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_232 bl[232] br[232] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_233 bl[233] br[233] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_234 bl[234] br[234] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_235 bl[235] br[235] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_236 bl[236] br[236] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_237 bl[237] br[237] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_238 bl[238] br[238] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_239 bl[239] br[239] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_240 bl[240] br[240] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_241 bl[241] br[241] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_242 bl[242] br[242] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_243 bl[243] br[243] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_244 bl[244] br[244] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_245 bl[245] br[245] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_246 bl[246] br[246] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_247 bl[247] br[247] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_248 bl[248] br[248] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_249 bl[249] br[249] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_250 bl[250] br[250] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_251 bl[251] br[251] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_252 bl[252] br[252] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_253 bl[253] br[253] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_254 bl[254] br[254] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_255 bl[255] br[255] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_112_0 bl[0] br[0] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_1 bl[1] br[1] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_2 bl[2] br[2] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_3 bl[3] br[3] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_4 bl[4] br[4] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_5 bl[5] br[5] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_6 bl[6] br[6] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_7 bl[7] br[7] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_8 bl[8] br[8] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_9 bl[9] br[9] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_10 bl[10] br[10] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_11 bl[11] br[11] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_12 bl[12] br[12] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_13 bl[13] br[13] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_14 bl[14] br[14] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_15 bl[15] br[15] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_16 bl[16] br[16] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_17 bl[17] br[17] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_18 bl[18] br[18] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_19 bl[19] br[19] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_20 bl[20] br[20] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_21 bl[21] br[21] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_22 bl[22] br[22] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_23 bl[23] br[23] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_24 bl[24] br[24] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_25 bl[25] br[25] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_26 bl[26] br[26] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_27 bl[27] br[27] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_28 bl[28] br[28] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_29 bl[29] br[29] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_30 bl[30] br[30] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_31 bl[31] br[31] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_32 bl[32] br[32] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_33 bl[33] br[33] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_34 bl[34] br[34] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_35 bl[35] br[35] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_36 bl[36] br[36] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_37 bl[37] br[37] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_38 bl[38] br[38] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_39 bl[39] br[39] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_40 bl[40] br[40] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_41 bl[41] br[41] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_42 bl[42] br[42] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_43 bl[43] br[43] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_44 bl[44] br[44] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_45 bl[45] br[45] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_46 bl[46] br[46] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_47 bl[47] br[47] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_48 bl[48] br[48] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_49 bl[49] br[49] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_50 bl[50] br[50] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_51 bl[51] br[51] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_52 bl[52] br[52] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_53 bl[53] br[53] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_54 bl[54] br[54] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_55 bl[55] br[55] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_56 bl[56] br[56] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_57 bl[57] br[57] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_58 bl[58] br[58] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_59 bl[59] br[59] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_60 bl[60] br[60] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_61 bl[61] br[61] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_62 bl[62] br[62] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_63 bl[63] br[63] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_64 bl[64] br[64] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_65 bl[65] br[65] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_66 bl[66] br[66] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_67 bl[67] br[67] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_68 bl[68] br[68] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_69 bl[69] br[69] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_70 bl[70] br[70] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_71 bl[71] br[71] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_72 bl[72] br[72] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_73 bl[73] br[73] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_74 bl[74] br[74] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_75 bl[75] br[75] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_76 bl[76] br[76] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_77 bl[77] br[77] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_78 bl[78] br[78] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_79 bl[79] br[79] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_80 bl[80] br[80] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_81 bl[81] br[81] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_82 bl[82] br[82] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_83 bl[83] br[83] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_84 bl[84] br[84] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_85 bl[85] br[85] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_86 bl[86] br[86] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_87 bl[87] br[87] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_88 bl[88] br[88] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_89 bl[89] br[89] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_90 bl[90] br[90] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_91 bl[91] br[91] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_92 bl[92] br[92] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_93 bl[93] br[93] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_94 bl[94] br[94] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_95 bl[95] br[95] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_96 bl[96] br[96] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_97 bl[97] br[97] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_98 bl[98] br[98] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_99 bl[99] br[99] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_100 bl[100] br[100] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_101 bl[101] br[101] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_102 bl[102] br[102] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_103 bl[103] br[103] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_104 bl[104] br[104] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_105 bl[105] br[105] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_106 bl[106] br[106] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_107 bl[107] br[107] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_108 bl[108] br[108] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_109 bl[109] br[109] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_110 bl[110] br[110] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_111 bl[111] br[111] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_112 bl[112] br[112] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_113 bl[113] br[113] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_114 bl[114] br[114] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_115 bl[115] br[115] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_116 bl[116] br[116] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_117 bl[117] br[117] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_118 bl[118] br[118] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_119 bl[119] br[119] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_120 bl[120] br[120] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_121 bl[121] br[121] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_122 bl[122] br[122] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_123 bl[123] br[123] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_124 bl[124] br[124] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_125 bl[125] br[125] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_126 bl[126] br[126] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_127 bl[127] br[127] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_128 bl[128] br[128] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_129 bl[129] br[129] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_130 bl[130] br[130] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_131 bl[131] br[131] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_132 bl[132] br[132] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_133 bl[133] br[133] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_134 bl[134] br[134] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_135 bl[135] br[135] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_136 bl[136] br[136] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_137 bl[137] br[137] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_138 bl[138] br[138] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_139 bl[139] br[139] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_140 bl[140] br[140] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_141 bl[141] br[141] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_142 bl[142] br[142] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_143 bl[143] br[143] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_144 bl[144] br[144] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_145 bl[145] br[145] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_146 bl[146] br[146] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_147 bl[147] br[147] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_148 bl[148] br[148] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_149 bl[149] br[149] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_150 bl[150] br[150] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_151 bl[151] br[151] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_152 bl[152] br[152] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_153 bl[153] br[153] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_154 bl[154] br[154] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_155 bl[155] br[155] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_156 bl[156] br[156] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_157 bl[157] br[157] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_158 bl[158] br[158] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_159 bl[159] br[159] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_160 bl[160] br[160] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_161 bl[161] br[161] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_162 bl[162] br[162] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_163 bl[163] br[163] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_164 bl[164] br[164] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_165 bl[165] br[165] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_166 bl[166] br[166] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_167 bl[167] br[167] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_168 bl[168] br[168] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_169 bl[169] br[169] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_170 bl[170] br[170] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_171 bl[171] br[171] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_172 bl[172] br[172] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_173 bl[173] br[173] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_174 bl[174] br[174] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_175 bl[175] br[175] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_176 bl[176] br[176] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_177 bl[177] br[177] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_178 bl[178] br[178] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_179 bl[179] br[179] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_180 bl[180] br[180] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_181 bl[181] br[181] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_182 bl[182] br[182] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_183 bl[183] br[183] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_184 bl[184] br[184] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_185 bl[185] br[185] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_186 bl[186] br[186] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_187 bl[187] br[187] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_188 bl[188] br[188] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_189 bl[189] br[189] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_190 bl[190] br[190] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_191 bl[191] br[191] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_192 bl[192] br[192] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_193 bl[193] br[193] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_194 bl[194] br[194] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_195 bl[195] br[195] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_196 bl[196] br[196] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_197 bl[197] br[197] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_198 bl[198] br[198] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_199 bl[199] br[199] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_200 bl[200] br[200] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_201 bl[201] br[201] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_202 bl[202] br[202] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_203 bl[203] br[203] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_204 bl[204] br[204] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_205 bl[205] br[205] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_206 bl[206] br[206] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_207 bl[207] br[207] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_208 bl[208] br[208] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_209 bl[209] br[209] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_210 bl[210] br[210] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_211 bl[211] br[211] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_212 bl[212] br[212] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_213 bl[213] br[213] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_214 bl[214] br[214] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_215 bl[215] br[215] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_216 bl[216] br[216] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_217 bl[217] br[217] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_218 bl[218] br[218] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_219 bl[219] br[219] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_220 bl[220] br[220] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_221 bl[221] br[221] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_222 bl[222] br[222] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_223 bl[223] br[223] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_224 bl[224] br[224] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_225 bl[225] br[225] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_226 bl[226] br[226] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_227 bl[227] br[227] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_228 bl[228] br[228] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_229 bl[229] br[229] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_230 bl[230] br[230] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_231 bl[231] br[231] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_232 bl[232] br[232] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_233 bl[233] br[233] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_234 bl[234] br[234] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_235 bl[235] br[235] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_236 bl[236] br[236] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_237 bl[237] br[237] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_238 bl[238] br[238] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_239 bl[239] br[239] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_240 bl[240] br[240] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_241 bl[241] br[241] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_242 bl[242] br[242] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_243 bl[243] br[243] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_244 bl[244] br[244] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_245 bl[245] br[245] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_246 bl[246] br[246] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_247 bl[247] br[247] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_248 bl[248] br[248] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_249 bl[249] br[249] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_250 bl[250] br[250] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_251 bl[251] br[251] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_252 bl[252] br[252] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_253 bl[253] br[253] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_254 bl[254] br[254] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_255 bl[255] br[255] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_113_0 bl[0] br[0] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_1 bl[1] br[1] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_2 bl[2] br[2] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_3 bl[3] br[3] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_4 bl[4] br[4] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_5 bl[5] br[5] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_6 bl[6] br[6] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_7 bl[7] br[7] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_8 bl[8] br[8] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_9 bl[9] br[9] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_10 bl[10] br[10] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_11 bl[11] br[11] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_12 bl[12] br[12] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_13 bl[13] br[13] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_14 bl[14] br[14] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_15 bl[15] br[15] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_16 bl[16] br[16] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_17 bl[17] br[17] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_18 bl[18] br[18] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_19 bl[19] br[19] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_20 bl[20] br[20] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_21 bl[21] br[21] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_22 bl[22] br[22] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_23 bl[23] br[23] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_24 bl[24] br[24] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_25 bl[25] br[25] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_26 bl[26] br[26] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_27 bl[27] br[27] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_28 bl[28] br[28] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_29 bl[29] br[29] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_30 bl[30] br[30] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_31 bl[31] br[31] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_32 bl[32] br[32] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_33 bl[33] br[33] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_34 bl[34] br[34] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_35 bl[35] br[35] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_36 bl[36] br[36] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_37 bl[37] br[37] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_38 bl[38] br[38] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_39 bl[39] br[39] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_40 bl[40] br[40] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_41 bl[41] br[41] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_42 bl[42] br[42] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_43 bl[43] br[43] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_44 bl[44] br[44] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_45 bl[45] br[45] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_46 bl[46] br[46] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_47 bl[47] br[47] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_48 bl[48] br[48] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_49 bl[49] br[49] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_50 bl[50] br[50] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_51 bl[51] br[51] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_52 bl[52] br[52] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_53 bl[53] br[53] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_54 bl[54] br[54] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_55 bl[55] br[55] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_56 bl[56] br[56] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_57 bl[57] br[57] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_58 bl[58] br[58] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_59 bl[59] br[59] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_60 bl[60] br[60] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_61 bl[61] br[61] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_62 bl[62] br[62] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_63 bl[63] br[63] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_64 bl[64] br[64] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_65 bl[65] br[65] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_66 bl[66] br[66] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_67 bl[67] br[67] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_68 bl[68] br[68] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_69 bl[69] br[69] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_70 bl[70] br[70] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_71 bl[71] br[71] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_72 bl[72] br[72] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_73 bl[73] br[73] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_74 bl[74] br[74] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_75 bl[75] br[75] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_76 bl[76] br[76] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_77 bl[77] br[77] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_78 bl[78] br[78] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_79 bl[79] br[79] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_80 bl[80] br[80] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_81 bl[81] br[81] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_82 bl[82] br[82] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_83 bl[83] br[83] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_84 bl[84] br[84] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_85 bl[85] br[85] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_86 bl[86] br[86] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_87 bl[87] br[87] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_88 bl[88] br[88] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_89 bl[89] br[89] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_90 bl[90] br[90] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_91 bl[91] br[91] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_92 bl[92] br[92] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_93 bl[93] br[93] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_94 bl[94] br[94] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_95 bl[95] br[95] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_96 bl[96] br[96] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_97 bl[97] br[97] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_98 bl[98] br[98] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_99 bl[99] br[99] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_100 bl[100] br[100] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_101 bl[101] br[101] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_102 bl[102] br[102] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_103 bl[103] br[103] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_104 bl[104] br[104] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_105 bl[105] br[105] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_106 bl[106] br[106] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_107 bl[107] br[107] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_108 bl[108] br[108] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_109 bl[109] br[109] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_110 bl[110] br[110] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_111 bl[111] br[111] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_112 bl[112] br[112] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_113 bl[113] br[113] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_114 bl[114] br[114] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_115 bl[115] br[115] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_116 bl[116] br[116] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_117 bl[117] br[117] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_118 bl[118] br[118] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_119 bl[119] br[119] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_120 bl[120] br[120] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_121 bl[121] br[121] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_122 bl[122] br[122] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_123 bl[123] br[123] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_124 bl[124] br[124] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_125 bl[125] br[125] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_126 bl[126] br[126] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_127 bl[127] br[127] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_128 bl[128] br[128] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_129 bl[129] br[129] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_130 bl[130] br[130] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_131 bl[131] br[131] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_132 bl[132] br[132] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_133 bl[133] br[133] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_134 bl[134] br[134] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_135 bl[135] br[135] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_136 bl[136] br[136] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_137 bl[137] br[137] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_138 bl[138] br[138] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_139 bl[139] br[139] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_140 bl[140] br[140] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_141 bl[141] br[141] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_142 bl[142] br[142] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_143 bl[143] br[143] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_144 bl[144] br[144] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_145 bl[145] br[145] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_146 bl[146] br[146] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_147 bl[147] br[147] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_148 bl[148] br[148] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_149 bl[149] br[149] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_150 bl[150] br[150] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_151 bl[151] br[151] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_152 bl[152] br[152] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_153 bl[153] br[153] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_154 bl[154] br[154] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_155 bl[155] br[155] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_156 bl[156] br[156] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_157 bl[157] br[157] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_158 bl[158] br[158] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_159 bl[159] br[159] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_160 bl[160] br[160] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_161 bl[161] br[161] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_162 bl[162] br[162] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_163 bl[163] br[163] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_164 bl[164] br[164] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_165 bl[165] br[165] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_166 bl[166] br[166] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_167 bl[167] br[167] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_168 bl[168] br[168] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_169 bl[169] br[169] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_170 bl[170] br[170] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_171 bl[171] br[171] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_172 bl[172] br[172] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_173 bl[173] br[173] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_174 bl[174] br[174] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_175 bl[175] br[175] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_176 bl[176] br[176] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_177 bl[177] br[177] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_178 bl[178] br[178] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_179 bl[179] br[179] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_180 bl[180] br[180] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_181 bl[181] br[181] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_182 bl[182] br[182] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_183 bl[183] br[183] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_184 bl[184] br[184] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_185 bl[185] br[185] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_186 bl[186] br[186] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_187 bl[187] br[187] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_188 bl[188] br[188] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_189 bl[189] br[189] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_190 bl[190] br[190] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_191 bl[191] br[191] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_192 bl[192] br[192] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_193 bl[193] br[193] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_194 bl[194] br[194] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_195 bl[195] br[195] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_196 bl[196] br[196] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_197 bl[197] br[197] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_198 bl[198] br[198] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_199 bl[199] br[199] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_200 bl[200] br[200] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_201 bl[201] br[201] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_202 bl[202] br[202] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_203 bl[203] br[203] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_204 bl[204] br[204] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_205 bl[205] br[205] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_206 bl[206] br[206] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_207 bl[207] br[207] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_208 bl[208] br[208] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_209 bl[209] br[209] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_210 bl[210] br[210] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_211 bl[211] br[211] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_212 bl[212] br[212] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_213 bl[213] br[213] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_214 bl[214] br[214] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_215 bl[215] br[215] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_216 bl[216] br[216] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_217 bl[217] br[217] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_218 bl[218] br[218] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_219 bl[219] br[219] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_220 bl[220] br[220] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_221 bl[221] br[221] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_222 bl[222] br[222] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_223 bl[223] br[223] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_224 bl[224] br[224] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_225 bl[225] br[225] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_226 bl[226] br[226] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_227 bl[227] br[227] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_228 bl[228] br[228] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_229 bl[229] br[229] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_230 bl[230] br[230] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_231 bl[231] br[231] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_232 bl[232] br[232] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_233 bl[233] br[233] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_234 bl[234] br[234] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_235 bl[235] br[235] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_236 bl[236] br[236] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_237 bl[237] br[237] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_238 bl[238] br[238] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_239 bl[239] br[239] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_240 bl[240] br[240] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_241 bl[241] br[241] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_242 bl[242] br[242] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_243 bl[243] br[243] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_244 bl[244] br[244] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_245 bl[245] br[245] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_246 bl[246] br[246] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_247 bl[247] br[247] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_248 bl[248] br[248] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_249 bl[249] br[249] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_250 bl[250] br[250] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_251 bl[251] br[251] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_252 bl[252] br[252] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_253 bl[253] br[253] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_254 bl[254] br[254] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_255 bl[255] br[255] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_114_0 bl[0] br[0] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_1 bl[1] br[1] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_2 bl[2] br[2] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_3 bl[3] br[3] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_4 bl[4] br[4] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_5 bl[5] br[5] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_6 bl[6] br[6] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_7 bl[7] br[7] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_8 bl[8] br[8] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_9 bl[9] br[9] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_10 bl[10] br[10] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_11 bl[11] br[11] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_12 bl[12] br[12] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_13 bl[13] br[13] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_14 bl[14] br[14] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_15 bl[15] br[15] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_16 bl[16] br[16] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_17 bl[17] br[17] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_18 bl[18] br[18] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_19 bl[19] br[19] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_20 bl[20] br[20] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_21 bl[21] br[21] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_22 bl[22] br[22] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_23 bl[23] br[23] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_24 bl[24] br[24] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_25 bl[25] br[25] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_26 bl[26] br[26] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_27 bl[27] br[27] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_28 bl[28] br[28] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_29 bl[29] br[29] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_30 bl[30] br[30] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_31 bl[31] br[31] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_32 bl[32] br[32] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_33 bl[33] br[33] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_34 bl[34] br[34] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_35 bl[35] br[35] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_36 bl[36] br[36] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_37 bl[37] br[37] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_38 bl[38] br[38] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_39 bl[39] br[39] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_40 bl[40] br[40] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_41 bl[41] br[41] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_42 bl[42] br[42] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_43 bl[43] br[43] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_44 bl[44] br[44] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_45 bl[45] br[45] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_46 bl[46] br[46] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_47 bl[47] br[47] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_48 bl[48] br[48] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_49 bl[49] br[49] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_50 bl[50] br[50] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_51 bl[51] br[51] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_52 bl[52] br[52] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_53 bl[53] br[53] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_54 bl[54] br[54] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_55 bl[55] br[55] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_56 bl[56] br[56] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_57 bl[57] br[57] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_58 bl[58] br[58] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_59 bl[59] br[59] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_60 bl[60] br[60] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_61 bl[61] br[61] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_62 bl[62] br[62] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_63 bl[63] br[63] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_64 bl[64] br[64] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_65 bl[65] br[65] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_66 bl[66] br[66] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_67 bl[67] br[67] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_68 bl[68] br[68] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_69 bl[69] br[69] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_70 bl[70] br[70] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_71 bl[71] br[71] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_72 bl[72] br[72] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_73 bl[73] br[73] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_74 bl[74] br[74] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_75 bl[75] br[75] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_76 bl[76] br[76] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_77 bl[77] br[77] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_78 bl[78] br[78] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_79 bl[79] br[79] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_80 bl[80] br[80] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_81 bl[81] br[81] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_82 bl[82] br[82] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_83 bl[83] br[83] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_84 bl[84] br[84] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_85 bl[85] br[85] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_86 bl[86] br[86] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_87 bl[87] br[87] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_88 bl[88] br[88] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_89 bl[89] br[89] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_90 bl[90] br[90] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_91 bl[91] br[91] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_92 bl[92] br[92] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_93 bl[93] br[93] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_94 bl[94] br[94] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_95 bl[95] br[95] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_96 bl[96] br[96] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_97 bl[97] br[97] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_98 bl[98] br[98] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_99 bl[99] br[99] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_100 bl[100] br[100] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_101 bl[101] br[101] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_102 bl[102] br[102] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_103 bl[103] br[103] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_104 bl[104] br[104] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_105 bl[105] br[105] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_106 bl[106] br[106] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_107 bl[107] br[107] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_108 bl[108] br[108] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_109 bl[109] br[109] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_110 bl[110] br[110] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_111 bl[111] br[111] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_112 bl[112] br[112] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_113 bl[113] br[113] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_114 bl[114] br[114] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_115 bl[115] br[115] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_116 bl[116] br[116] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_117 bl[117] br[117] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_118 bl[118] br[118] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_119 bl[119] br[119] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_120 bl[120] br[120] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_121 bl[121] br[121] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_122 bl[122] br[122] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_123 bl[123] br[123] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_124 bl[124] br[124] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_125 bl[125] br[125] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_126 bl[126] br[126] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_127 bl[127] br[127] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_128 bl[128] br[128] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_129 bl[129] br[129] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_130 bl[130] br[130] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_131 bl[131] br[131] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_132 bl[132] br[132] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_133 bl[133] br[133] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_134 bl[134] br[134] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_135 bl[135] br[135] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_136 bl[136] br[136] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_137 bl[137] br[137] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_138 bl[138] br[138] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_139 bl[139] br[139] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_140 bl[140] br[140] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_141 bl[141] br[141] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_142 bl[142] br[142] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_143 bl[143] br[143] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_144 bl[144] br[144] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_145 bl[145] br[145] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_146 bl[146] br[146] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_147 bl[147] br[147] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_148 bl[148] br[148] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_149 bl[149] br[149] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_150 bl[150] br[150] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_151 bl[151] br[151] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_152 bl[152] br[152] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_153 bl[153] br[153] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_154 bl[154] br[154] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_155 bl[155] br[155] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_156 bl[156] br[156] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_157 bl[157] br[157] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_158 bl[158] br[158] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_159 bl[159] br[159] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_160 bl[160] br[160] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_161 bl[161] br[161] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_162 bl[162] br[162] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_163 bl[163] br[163] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_164 bl[164] br[164] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_165 bl[165] br[165] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_166 bl[166] br[166] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_167 bl[167] br[167] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_168 bl[168] br[168] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_169 bl[169] br[169] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_170 bl[170] br[170] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_171 bl[171] br[171] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_172 bl[172] br[172] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_173 bl[173] br[173] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_174 bl[174] br[174] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_175 bl[175] br[175] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_176 bl[176] br[176] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_177 bl[177] br[177] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_178 bl[178] br[178] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_179 bl[179] br[179] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_180 bl[180] br[180] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_181 bl[181] br[181] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_182 bl[182] br[182] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_183 bl[183] br[183] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_184 bl[184] br[184] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_185 bl[185] br[185] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_186 bl[186] br[186] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_187 bl[187] br[187] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_188 bl[188] br[188] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_189 bl[189] br[189] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_190 bl[190] br[190] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_191 bl[191] br[191] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_192 bl[192] br[192] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_193 bl[193] br[193] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_194 bl[194] br[194] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_195 bl[195] br[195] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_196 bl[196] br[196] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_197 bl[197] br[197] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_198 bl[198] br[198] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_199 bl[199] br[199] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_200 bl[200] br[200] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_201 bl[201] br[201] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_202 bl[202] br[202] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_203 bl[203] br[203] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_204 bl[204] br[204] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_205 bl[205] br[205] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_206 bl[206] br[206] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_207 bl[207] br[207] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_208 bl[208] br[208] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_209 bl[209] br[209] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_210 bl[210] br[210] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_211 bl[211] br[211] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_212 bl[212] br[212] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_213 bl[213] br[213] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_214 bl[214] br[214] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_215 bl[215] br[215] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_216 bl[216] br[216] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_217 bl[217] br[217] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_218 bl[218] br[218] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_219 bl[219] br[219] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_220 bl[220] br[220] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_221 bl[221] br[221] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_222 bl[222] br[222] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_223 bl[223] br[223] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_224 bl[224] br[224] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_225 bl[225] br[225] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_226 bl[226] br[226] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_227 bl[227] br[227] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_228 bl[228] br[228] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_229 bl[229] br[229] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_230 bl[230] br[230] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_231 bl[231] br[231] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_232 bl[232] br[232] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_233 bl[233] br[233] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_234 bl[234] br[234] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_235 bl[235] br[235] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_236 bl[236] br[236] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_237 bl[237] br[237] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_238 bl[238] br[238] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_239 bl[239] br[239] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_240 bl[240] br[240] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_241 bl[241] br[241] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_242 bl[242] br[242] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_243 bl[243] br[243] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_244 bl[244] br[244] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_245 bl[245] br[245] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_246 bl[246] br[246] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_247 bl[247] br[247] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_248 bl[248] br[248] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_249 bl[249] br[249] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_250 bl[250] br[250] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_251 bl[251] br[251] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_252 bl[252] br[252] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_253 bl[253] br[253] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_254 bl[254] br[254] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_255 bl[255] br[255] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_115_0 bl[0] br[0] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_1 bl[1] br[1] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_2 bl[2] br[2] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_3 bl[3] br[3] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_4 bl[4] br[4] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_5 bl[5] br[5] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_6 bl[6] br[6] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_7 bl[7] br[7] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_8 bl[8] br[8] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_9 bl[9] br[9] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_10 bl[10] br[10] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_11 bl[11] br[11] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_12 bl[12] br[12] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_13 bl[13] br[13] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_14 bl[14] br[14] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_15 bl[15] br[15] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_16 bl[16] br[16] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_17 bl[17] br[17] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_18 bl[18] br[18] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_19 bl[19] br[19] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_20 bl[20] br[20] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_21 bl[21] br[21] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_22 bl[22] br[22] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_23 bl[23] br[23] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_24 bl[24] br[24] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_25 bl[25] br[25] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_26 bl[26] br[26] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_27 bl[27] br[27] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_28 bl[28] br[28] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_29 bl[29] br[29] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_30 bl[30] br[30] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_31 bl[31] br[31] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_32 bl[32] br[32] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_33 bl[33] br[33] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_34 bl[34] br[34] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_35 bl[35] br[35] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_36 bl[36] br[36] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_37 bl[37] br[37] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_38 bl[38] br[38] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_39 bl[39] br[39] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_40 bl[40] br[40] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_41 bl[41] br[41] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_42 bl[42] br[42] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_43 bl[43] br[43] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_44 bl[44] br[44] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_45 bl[45] br[45] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_46 bl[46] br[46] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_47 bl[47] br[47] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_48 bl[48] br[48] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_49 bl[49] br[49] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_50 bl[50] br[50] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_51 bl[51] br[51] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_52 bl[52] br[52] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_53 bl[53] br[53] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_54 bl[54] br[54] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_55 bl[55] br[55] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_56 bl[56] br[56] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_57 bl[57] br[57] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_58 bl[58] br[58] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_59 bl[59] br[59] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_60 bl[60] br[60] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_61 bl[61] br[61] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_62 bl[62] br[62] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_63 bl[63] br[63] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_64 bl[64] br[64] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_65 bl[65] br[65] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_66 bl[66] br[66] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_67 bl[67] br[67] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_68 bl[68] br[68] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_69 bl[69] br[69] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_70 bl[70] br[70] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_71 bl[71] br[71] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_72 bl[72] br[72] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_73 bl[73] br[73] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_74 bl[74] br[74] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_75 bl[75] br[75] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_76 bl[76] br[76] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_77 bl[77] br[77] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_78 bl[78] br[78] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_79 bl[79] br[79] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_80 bl[80] br[80] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_81 bl[81] br[81] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_82 bl[82] br[82] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_83 bl[83] br[83] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_84 bl[84] br[84] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_85 bl[85] br[85] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_86 bl[86] br[86] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_87 bl[87] br[87] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_88 bl[88] br[88] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_89 bl[89] br[89] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_90 bl[90] br[90] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_91 bl[91] br[91] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_92 bl[92] br[92] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_93 bl[93] br[93] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_94 bl[94] br[94] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_95 bl[95] br[95] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_96 bl[96] br[96] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_97 bl[97] br[97] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_98 bl[98] br[98] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_99 bl[99] br[99] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_100 bl[100] br[100] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_101 bl[101] br[101] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_102 bl[102] br[102] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_103 bl[103] br[103] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_104 bl[104] br[104] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_105 bl[105] br[105] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_106 bl[106] br[106] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_107 bl[107] br[107] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_108 bl[108] br[108] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_109 bl[109] br[109] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_110 bl[110] br[110] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_111 bl[111] br[111] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_112 bl[112] br[112] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_113 bl[113] br[113] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_114 bl[114] br[114] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_115 bl[115] br[115] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_116 bl[116] br[116] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_117 bl[117] br[117] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_118 bl[118] br[118] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_119 bl[119] br[119] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_120 bl[120] br[120] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_121 bl[121] br[121] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_122 bl[122] br[122] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_123 bl[123] br[123] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_124 bl[124] br[124] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_125 bl[125] br[125] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_126 bl[126] br[126] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_127 bl[127] br[127] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_128 bl[128] br[128] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_129 bl[129] br[129] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_130 bl[130] br[130] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_131 bl[131] br[131] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_132 bl[132] br[132] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_133 bl[133] br[133] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_134 bl[134] br[134] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_135 bl[135] br[135] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_136 bl[136] br[136] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_137 bl[137] br[137] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_138 bl[138] br[138] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_139 bl[139] br[139] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_140 bl[140] br[140] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_141 bl[141] br[141] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_142 bl[142] br[142] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_143 bl[143] br[143] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_144 bl[144] br[144] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_145 bl[145] br[145] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_146 bl[146] br[146] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_147 bl[147] br[147] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_148 bl[148] br[148] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_149 bl[149] br[149] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_150 bl[150] br[150] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_151 bl[151] br[151] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_152 bl[152] br[152] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_153 bl[153] br[153] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_154 bl[154] br[154] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_155 bl[155] br[155] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_156 bl[156] br[156] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_157 bl[157] br[157] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_158 bl[158] br[158] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_159 bl[159] br[159] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_160 bl[160] br[160] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_161 bl[161] br[161] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_162 bl[162] br[162] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_163 bl[163] br[163] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_164 bl[164] br[164] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_165 bl[165] br[165] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_166 bl[166] br[166] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_167 bl[167] br[167] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_168 bl[168] br[168] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_169 bl[169] br[169] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_170 bl[170] br[170] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_171 bl[171] br[171] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_172 bl[172] br[172] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_173 bl[173] br[173] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_174 bl[174] br[174] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_175 bl[175] br[175] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_176 bl[176] br[176] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_177 bl[177] br[177] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_178 bl[178] br[178] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_179 bl[179] br[179] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_180 bl[180] br[180] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_181 bl[181] br[181] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_182 bl[182] br[182] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_183 bl[183] br[183] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_184 bl[184] br[184] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_185 bl[185] br[185] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_186 bl[186] br[186] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_187 bl[187] br[187] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_188 bl[188] br[188] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_189 bl[189] br[189] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_190 bl[190] br[190] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_191 bl[191] br[191] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_192 bl[192] br[192] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_193 bl[193] br[193] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_194 bl[194] br[194] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_195 bl[195] br[195] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_196 bl[196] br[196] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_197 bl[197] br[197] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_198 bl[198] br[198] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_199 bl[199] br[199] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_200 bl[200] br[200] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_201 bl[201] br[201] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_202 bl[202] br[202] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_203 bl[203] br[203] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_204 bl[204] br[204] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_205 bl[205] br[205] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_206 bl[206] br[206] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_207 bl[207] br[207] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_208 bl[208] br[208] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_209 bl[209] br[209] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_210 bl[210] br[210] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_211 bl[211] br[211] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_212 bl[212] br[212] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_213 bl[213] br[213] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_214 bl[214] br[214] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_215 bl[215] br[215] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_216 bl[216] br[216] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_217 bl[217] br[217] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_218 bl[218] br[218] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_219 bl[219] br[219] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_220 bl[220] br[220] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_221 bl[221] br[221] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_222 bl[222] br[222] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_223 bl[223] br[223] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_224 bl[224] br[224] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_225 bl[225] br[225] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_226 bl[226] br[226] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_227 bl[227] br[227] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_228 bl[228] br[228] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_229 bl[229] br[229] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_230 bl[230] br[230] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_231 bl[231] br[231] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_232 bl[232] br[232] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_233 bl[233] br[233] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_234 bl[234] br[234] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_235 bl[235] br[235] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_236 bl[236] br[236] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_237 bl[237] br[237] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_238 bl[238] br[238] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_239 bl[239] br[239] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_240 bl[240] br[240] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_241 bl[241] br[241] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_242 bl[242] br[242] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_243 bl[243] br[243] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_244 bl[244] br[244] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_245 bl[245] br[245] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_246 bl[246] br[246] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_247 bl[247] br[247] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_248 bl[248] br[248] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_249 bl[249] br[249] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_250 bl[250] br[250] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_251 bl[251] br[251] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_252 bl[252] br[252] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_253 bl[253] br[253] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_254 bl[254] br[254] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_255 bl[255] br[255] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_116_0 bl[0] br[0] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_1 bl[1] br[1] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_2 bl[2] br[2] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_3 bl[3] br[3] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_4 bl[4] br[4] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_5 bl[5] br[5] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_6 bl[6] br[6] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_7 bl[7] br[7] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_8 bl[8] br[8] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_9 bl[9] br[9] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_10 bl[10] br[10] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_11 bl[11] br[11] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_12 bl[12] br[12] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_13 bl[13] br[13] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_14 bl[14] br[14] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_15 bl[15] br[15] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_16 bl[16] br[16] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_17 bl[17] br[17] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_18 bl[18] br[18] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_19 bl[19] br[19] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_20 bl[20] br[20] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_21 bl[21] br[21] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_22 bl[22] br[22] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_23 bl[23] br[23] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_24 bl[24] br[24] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_25 bl[25] br[25] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_26 bl[26] br[26] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_27 bl[27] br[27] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_28 bl[28] br[28] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_29 bl[29] br[29] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_30 bl[30] br[30] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_31 bl[31] br[31] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_32 bl[32] br[32] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_33 bl[33] br[33] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_34 bl[34] br[34] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_35 bl[35] br[35] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_36 bl[36] br[36] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_37 bl[37] br[37] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_38 bl[38] br[38] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_39 bl[39] br[39] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_40 bl[40] br[40] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_41 bl[41] br[41] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_42 bl[42] br[42] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_43 bl[43] br[43] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_44 bl[44] br[44] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_45 bl[45] br[45] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_46 bl[46] br[46] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_47 bl[47] br[47] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_48 bl[48] br[48] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_49 bl[49] br[49] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_50 bl[50] br[50] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_51 bl[51] br[51] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_52 bl[52] br[52] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_53 bl[53] br[53] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_54 bl[54] br[54] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_55 bl[55] br[55] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_56 bl[56] br[56] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_57 bl[57] br[57] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_58 bl[58] br[58] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_59 bl[59] br[59] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_60 bl[60] br[60] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_61 bl[61] br[61] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_62 bl[62] br[62] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_63 bl[63] br[63] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_64 bl[64] br[64] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_65 bl[65] br[65] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_66 bl[66] br[66] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_67 bl[67] br[67] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_68 bl[68] br[68] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_69 bl[69] br[69] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_70 bl[70] br[70] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_71 bl[71] br[71] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_72 bl[72] br[72] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_73 bl[73] br[73] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_74 bl[74] br[74] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_75 bl[75] br[75] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_76 bl[76] br[76] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_77 bl[77] br[77] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_78 bl[78] br[78] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_79 bl[79] br[79] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_80 bl[80] br[80] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_81 bl[81] br[81] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_82 bl[82] br[82] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_83 bl[83] br[83] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_84 bl[84] br[84] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_85 bl[85] br[85] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_86 bl[86] br[86] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_87 bl[87] br[87] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_88 bl[88] br[88] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_89 bl[89] br[89] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_90 bl[90] br[90] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_91 bl[91] br[91] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_92 bl[92] br[92] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_93 bl[93] br[93] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_94 bl[94] br[94] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_95 bl[95] br[95] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_96 bl[96] br[96] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_97 bl[97] br[97] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_98 bl[98] br[98] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_99 bl[99] br[99] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_100 bl[100] br[100] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_101 bl[101] br[101] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_102 bl[102] br[102] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_103 bl[103] br[103] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_104 bl[104] br[104] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_105 bl[105] br[105] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_106 bl[106] br[106] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_107 bl[107] br[107] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_108 bl[108] br[108] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_109 bl[109] br[109] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_110 bl[110] br[110] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_111 bl[111] br[111] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_112 bl[112] br[112] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_113 bl[113] br[113] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_114 bl[114] br[114] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_115 bl[115] br[115] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_116 bl[116] br[116] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_117 bl[117] br[117] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_118 bl[118] br[118] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_119 bl[119] br[119] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_120 bl[120] br[120] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_121 bl[121] br[121] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_122 bl[122] br[122] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_123 bl[123] br[123] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_124 bl[124] br[124] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_125 bl[125] br[125] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_126 bl[126] br[126] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_127 bl[127] br[127] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_128 bl[128] br[128] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_129 bl[129] br[129] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_130 bl[130] br[130] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_131 bl[131] br[131] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_132 bl[132] br[132] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_133 bl[133] br[133] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_134 bl[134] br[134] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_135 bl[135] br[135] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_136 bl[136] br[136] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_137 bl[137] br[137] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_138 bl[138] br[138] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_139 bl[139] br[139] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_140 bl[140] br[140] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_141 bl[141] br[141] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_142 bl[142] br[142] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_143 bl[143] br[143] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_144 bl[144] br[144] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_145 bl[145] br[145] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_146 bl[146] br[146] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_147 bl[147] br[147] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_148 bl[148] br[148] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_149 bl[149] br[149] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_150 bl[150] br[150] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_151 bl[151] br[151] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_152 bl[152] br[152] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_153 bl[153] br[153] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_154 bl[154] br[154] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_155 bl[155] br[155] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_156 bl[156] br[156] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_157 bl[157] br[157] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_158 bl[158] br[158] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_159 bl[159] br[159] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_160 bl[160] br[160] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_161 bl[161] br[161] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_162 bl[162] br[162] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_163 bl[163] br[163] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_164 bl[164] br[164] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_165 bl[165] br[165] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_166 bl[166] br[166] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_167 bl[167] br[167] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_168 bl[168] br[168] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_169 bl[169] br[169] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_170 bl[170] br[170] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_171 bl[171] br[171] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_172 bl[172] br[172] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_173 bl[173] br[173] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_174 bl[174] br[174] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_175 bl[175] br[175] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_176 bl[176] br[176] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_177 bl[177] br[177] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_178 bl[178] br[178] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_179 bl[179] br[179] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_180 bl[180] br[180] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_181 bl[181] br[181] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_182 bl[182] br[182] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_183 bl[183] br[183] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_184 bl[184] br[184] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_185 bl[185] br[185] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_186 bl[186] br[186] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_187 bl[187] br[187] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_188 bl[188] br[188] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_189 bl[189] br[189] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_190 bl[190] br[190] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_191 bl[191] br[191] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_192 bl[192] br[192] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_193 bl[193] br[193] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_194 bl[194] br[194] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_195 bl[195] br[195] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_196 bl[196] br[196] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_197 bl[197] br[197] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_198 bl[198] br[198] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_199 bl[199] br[199] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_200 bl[200] br[200] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_201 bl[201] br[201] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_202 bl[202] br[202] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_203 bl[203] br[203] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_204 bl[204] br[204] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_205 bl[205] br[205] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_206 bl[206] br[206] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_207 bl[207] br[207] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_208 bl[208] br[208] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_209 bl[209] br[209] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_210 bl[210] br[210] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_211 bl[211] br[211] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_212 bl[212] br[212] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_213 bl[213] br[213] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_214 bl[214] br[214] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_215 bl[215] br[215] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_216 bl[216] br[216] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_217 bl[217] br[217] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_218 bl[218] br[218] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_219 bl[219] br[219] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_220 bl[220] br[220] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_221 bl[221] br[221] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_222 bl[222] br[222] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_223 bl[223] br[223] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_224 bl[224] br[224] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_225 bl[225] br[225] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_226 bl[226] br[226] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_227 bl[227] br[227] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_228 bl[228] br[228] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_229 bl[229] br[229] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_230 bl[230] br[230] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_231 bl[231] br[231] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_232 bl[232] br[232] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_233 bl[233] br[233] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_234 bl[234] br[234] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_235 bl[235] br[235] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_236 bl[236] br[236] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_237 bl[237] br[237] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_238 bl[238] br[238] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_239 bl[239] br[239] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_240 bl[240] br[240] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_241 bl[241] br[241] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_242 bl[242] br[242] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_243 bl[243] br[243] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_244 bl[244] br[244] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_245 bl[245] br[245] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_246 bl[246] br[246] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_247 bl[247] br[247] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_248 bl[248] br[248] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_249 bl[249] br[249] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_250 bl[250] br[250] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_251 bl[251] br[251] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_252 bl[252] br[252] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_253 bl[253] br[253] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_254 bl[254] br[254] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_255 bl[255] br[255] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_117_0 bl[0] br[0] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_1 bl[1] br[1] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_2 bl[2] br[2] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_3 bl[3] br[3] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_4 bl[4] br[4] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_5 bl[5] br[5] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_6 bl[6] br[6] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_7 bl[7] br[7] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_8 bl[8] br[8] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_9 bl[9] br[9] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_10 bl[10] br[10] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_11 bl[11] br[11] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_12 bl[12] br[12] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_13 bl[13] br[13] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_14 bl[14] br[14] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_15 bl[15] br[15] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_16 bl[16] br[16] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_17 bl[17] br[17] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_18 bl[18] br[18] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_19 bl[19] br[19] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_20 bl[20] br[20] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_21 bl[21] br[21] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_22 bl[22] br[22] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_23 bl[23] br[23] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_24 bl[24] br[24] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_25 bl[25] br[25] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_26 bl[26] br[26] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_27 bl[27] br[27] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_28 bl[28] br[28] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_29 bl[29] br[29] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_30 bl[30] br[30] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_31 bl[31] br[31] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_32 bl[32] br[32] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_33 bl[33] br[33] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_34 bl[34] br[34] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_35 bl[35] br[35] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_36 bl[36] br[36] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_37 bl[37] br[37] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_38 bl[38] br[38] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_39 bl[39] br[39] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_40 bl[40] br[40] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_41 bl[41] br[41] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_42 bl[42] br[42] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_43 bl[43] br[43] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_44 bl[44] br[44] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_45 bl[45] br[45] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_46 bl[46] br[46] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_47 bl[47] br[47] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_48 bl[48] br[48] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_49 bl[49] br[49] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_50 bl[50] br[50] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_51 bl[51] br[51] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_52 bl[52] br[52] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_53 bl[53] br[53] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_54 bl[54] br[54] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_55 bl[55] br[55] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_56 bl[56] br[56] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_57 bl[57] br[57] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_58 bl[58] br[58] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_59 bl[59] br[59] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_60 bl[60] br[60] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_61 bl[61] br[61] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_62 bl[62] br[62] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_63 bl[63] br[63] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_64 bl[64] br[64] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_65 bl[65] br[65] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_66 bl[66] br[66] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_67 bl[67] br[67] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_68 bl[68] br[68] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_69 bl[69] br[69] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_70 bl[70] br[70] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_71 bl[71] br[71] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_72 bl[72] br[72] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_73 bl[73] br[73] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_74 bl[74] br[74] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_75 bl[75] br[75] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_76 bl[76] br[76] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_77 bl[77] br[77] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_78 bl[78] br[78] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_79 bl[79] br[79] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_80 bl[80] br[80] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_81 bl[81] br[81] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_82 bl[82] br[82] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_83 bl[83] br[83] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_84 bl[84] br[84] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_85 bl[85] br[85] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_86 bl[86] br[86] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_87 bl[87] br[87] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_88 bl[88] br[88] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_89 bl[89] br[89] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_90 bl[90] br[90] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_91 bl[91] br[91] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_92 bl[92] br[92] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_93 bl[93] br[93] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_94 bl[94] br[94] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_95 bl[95] br[95] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_96 bl[96] br[96] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_97 bl[97] br[97] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_98 bl[98] br[98] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_99 bl[99] br[99] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_100 bl[100] br[100] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_101 bl[101] br[101] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_102 bl[102] br[102] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_103 bl[103] br[103] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_104 bl[104] br[104] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_105 bl[105] br[105] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_106 bl[106] br[106] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_107 bl[107] br[107] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_108 bl[108] br[108] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_109 bl[109] br[109] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_110 bl[110] br[110] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_111 bl[111] br[111] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_112 bl[112] br[112] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_113 bl[113] br[113] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_114 bl[114] br[114] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_115 bl[115] br[115] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_116 bl[116] br[116] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_117 bl[117] br[117] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_118 bl[118] br[118] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_119 bl[119] br[119] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_120 bl[120] br[120] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_121 bl[121] br[121] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_122 bl[122] br[122] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_123 bl[123] br[123] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_124 bl[124] br[124] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_125 bl[125] br[125] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_126 bl[126] br[126] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_127 bl[127] br[127] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_128 bl[128] br[128] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_129 bl[129] br[129] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_130 bl[130] br[130] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_131 bl[131] br[131] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_132 bl[132] br[132] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_133 bl[133] br[133] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_134 bl[134] br[134] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_135 bl[135] br[135] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_136 bl[136] br[136] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_137 bl[137] br[137] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_138 bl[138] br[138] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_139 bl[139] br[139] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_140 bl[140] br[140] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_141 bl[141] br[141] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_142 bl[142] br[142] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_143 bl[143] br[143] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_144 bl[144] br[144] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_145 bl[145] br[145] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_146 bl[146] br[146] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_147 bl[147] br[147] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_148 bl[148] br[148] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_149 bl[149] br[149] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_150 bl[150] br[150] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_151 bl[151] br[151] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_152 bl[152] br[152] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_153 bl[153] br[153] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_154 bl[154] br[154] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_155 bl[155] br[155] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_156 bl[156] br[156] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_157 bl[157] br[157] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_158 bl[158] br[158] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_159 bl[159] br[159] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_160 bl[160] br[160] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_161 bl[161] br[161] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_162 bl[162] br[162] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_163 bl[163] br[163] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_164 bl[164] br[164] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_165 bl[165] br[165] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_166 bl[166] br[166] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_167 bl[167] br[167] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_168 bl[168] br[168] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_169 bl[169] br[169] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_170 bl[170] br[170] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_171 bl[171] br[171] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_172 bl[172] br[172] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_173 bl[173] br[173] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_174 bl[174] br[174] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_175 bl[175] br[175] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_176 bl[176] br[176] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_177 bl[177] br[177] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_178 bl[178] br[178] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_179 bl[179] br[179] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_180 bl[180] br[180] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_181 bl[181] br[181] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_182 bl[182] br[182] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_183 bl[183] br[183] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_184 bl[184] br[184] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_185 bl[185] br[185] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_186 bl[186] br[186] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_187 bl[187] br[187] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_188 bl[188] br[188] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_189 bl[189] br[189] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_190 bl[190] br[190] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_191 bl[191] br[191] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_192 bl[192] br[192] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_193 bl[193] br[193] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_194 bl[194] br[194] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_195 bl[195] br[195] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_196 bl[196] br[196] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_197 bl[197] br[197] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_198 bl[198] br[198] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_199 bl[199] br[199] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_200 bl[200] br[200] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_201 bl[201] br[201] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_202 bl[202] br[202] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_203 bl[203] br[203] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_204 bl[204] br[204] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_205 bl[205] br[205] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_206 bl[206] br[206] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_207 bl[207] br[207] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_208 bl[208] br[208] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_209 bl[209] br[209] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_210 bl[210] br[210] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_211 bl[211] br[211] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_212 bl[212] br[212] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_213 bl[213] br[213] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_214 bl[214] br[214] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_215 bl[215] br[215] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_216 bl[216] br[216] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_217 bl[217] br[217] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_218 bl[218] br[218] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_219 bl[219] br[219] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_220 bl[220] br[220] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_221 bl[221] br[221] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_222 bl[222] br[222] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_223 bl[223] br[223] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_224 bl[224] br[224] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_225 bl[225] br[225] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_226 bl[226] br[226] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_227 bl[227] br[227] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_228 bl[228] br[228] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_229 bl[229] br[229] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_230 bl[230] br[230] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_231 bl[231] br[231] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_232 bl[232] br[232] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_233 bl[233] br[233] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_234 bl[234] br[234] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_235 bl[235] br[235] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_236 bl[236] br[236] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_237 bl[237] br[237] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_238 bl[238] br[238] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_239 bl[239] br[239] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_240 bl[240] br[240] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_241 bl[241] br[241] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_242 bl[242] br[242] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_243 bl[243] br[243] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_244 bl[244] br[244] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_245 bl[245] br[245] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_246 bl[246] br[246] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_247 bl[247] br[247] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_248 bl[248] br[248] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_249 bl[249] br[249] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_250 bl[250] br[250] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_251 bl[251] br[251] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_252 bl[252] br[252] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_253 bl[253] br[253] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_254 bl[254] br[254] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_255 bl[255] br[255] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_118_0 bl[0] br[0] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_1 bl[1] br[1] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_2 bl[2] br[2] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_3 bl[3] br[3] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_4 bl[4] br[4] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_5 bl[5] br[5] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_6 bl[6] br[6] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_7 bl[7] br[7] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_8 bl[8] br[8] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_9 bl[9] br[9] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_10 bl[10] br[10] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_11 bl[11] br[11] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_12 bl[12] br[12] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_13 bl[13] br[13] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_14 bl[14] br[14] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_15 bl[15] br[15] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_16 bl[16] br[16] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_17 bl[17] br[17] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_18 bl[18] br[18] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_19 bl[19] br[19] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_20 bl[20] br[20] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_21 bl[21] br[21] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_22 bl[22] br[22] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_23 bl[23] br[23] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_24 bl[24] br[24] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_25 bl[25] br[25] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_26 bl[26] br[26] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_27 bl[27] br[27] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_28 bl[28] br[28] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_29 bl[29] br[29] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_30 bl[30] br[30] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_31 bl[31] br[31] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_32 bl[32] br[32] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_33 bl[33] br[33] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_34 bl[34] br[34] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_35 bl[35] br[35] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_36 bl[36] br[36] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_37 bl[37] br[37] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_38 bl[38] br[38] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_39 bl[39] br[39] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_40 bl[40] br[40] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_41 bl[41] br[41] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_42 bl[42] br[42] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_43 bl[43] br[43] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_44 bl[44] br[44] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_45 bl[45] br[45] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_46 bl[46] br[46] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_47 bl[47] br[47] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_48 bl[48] br[48] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_49 bl[49] br[49] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_50 bl[50] br[50] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_51 bl[51] br[51] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_52 bl[52] br[52] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_53 bl[53] br[53] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_54 bl[54] br[54] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_55 bl[55] br[55] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_56 bl[56] br[56] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_57 bl[57] br[57] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_58 bl[58] br[58] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_59 bl[59] br[59] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_60 bl[60] br[60] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_61 bl[61] br[61] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_62 bl[62] br[62] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_63 bl[63] br[63] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_64 bl[64] br[64] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_65 bl[65] br[65] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_66 bl[66] br[66] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_67 bl[67] br[67] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_68 bl[68] br[68] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_69 bl[69] br[69] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_70 bl[70] br[70] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_71 bl[71] br[71] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_72 bl[72] br[72] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_73 bl[73] br[73] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_74 bl[74] br[74] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_75 bl[75] br[75] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_76 bl[76] br[76] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_77 bl[77] br[77] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_78 bl[78] br[78] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_79 bl[79] br[79] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_80 bl[80] br[80] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_81 bl[81] br[81] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_82 bl[82] br[82] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_83 bl[83] br[83] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_84 bl[84] br[84] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_85 bl[85] br[85] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_86 bl[86] br[86] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_87 bl[87] br[87] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_88 bl[88] br[88] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_89 bl[89] br[89] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_90 bl[90] br[90] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_91 bl[91] br[91] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_92 bl[92] br[92] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_93 bl[93] br[93] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_94 bl[94] br[94] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_95 bl[95] br[95] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_96 bl[96] br[96] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_97 bl[97] br[97] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_98 bl[98] br[98] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_99 bl[99] br[99] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_100 bl[100] br[100] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_101 bl[101] br[101] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_102 bl[102] br[102] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_103 bl[103] br[103] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_104 bl[104] br[104] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_105 bl[105] br[105] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_106 bl[106] br[106] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_107 bl[107] br[107] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_108 bl[108] br[108] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_109 bl[109] br[109] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_110 bl[110] br[110] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_111 bl[111] br[111] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_112 bl[112] br[112] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_113 bl[113] br[113] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_114 bl[114] br[114] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_115 bl[115] br[115] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_116 bl[116] br[116] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_117 bl[117] br[117] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_118 bl[118] br[118] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_119 bl[119] br[119] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_120 bl[120] br[120] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_121 bl[121] br[121] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_122 bl[122] br[122] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_123 bl[123] br[123] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_124 bl[124] br[124] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_125 bl[125] br[125] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_126 bl[126] br[126] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_127 bl[127] br[127] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_128 bl[128] br[128] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_129 bl[129] br[129] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_130 bl[130] br[130] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_131 bl[131] br[131] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_132 bl[132] br[132] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_133 bl[133] br[133] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_134 bl[134] br[134] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_135 bl[135] br[135] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_136 bl[136] br[136] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_137 bl[137] br[137] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_138 bl[138] br[138] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_139 bl[139] br[139] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_140 bl[140] br[140] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_141 bl[141] br[141] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_142 bl[142] br[142] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_143 bl[143] br[143] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_144 bl[144] br[144] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_145 bl[145] br[145] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_146 bl[146] br[146] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_147 bl[147] br[147] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_148 bl[148] br[148] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_149 bl[149] br[149] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_150 bl[150] br[150] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_151 bl[151] br[151] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_152 bl[152] br[152] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_153 bl[153] br[153] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_154 bl[154] br[154] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_155 bl[155] br[155] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_156 bl[156] br[156] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_157 bl[157] br[157] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_158 bl[158] br[158] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_159 bl[159] br[159] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_160 bl[160] br[160] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_161 bl[161] br[161] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_162 bl[162] br[162] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_163 bl[163] br[163] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_164 bl[164] br[164] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_165 bl[165] br[165] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_166 bl[166] br[166] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_167 bl[167] br[167] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_168 bl[168] br[168] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_169 bl[169] br[169] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_170 bl[170] br[170] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_171 bl[171] br[171] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_172 bl[172] br[172] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_173 bl[173] br[173] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_174 bl[174] br[174] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_175 bl[175] br[175] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_176 bl[176] br[176] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_177 bl[177] br[177] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_178 bl[178] br[178] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_179 bl[179] br[179] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_180 bl[180] br[180] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_181 bl[181] br[181] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_182 bl[182] br[182] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_183 bl[183] br[183] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_184 bl[184] br[184] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_185 bl[185] br[185] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_186 bl[186] br[186] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_187 bl[187] br[187] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_188 bl[188] br[188] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_189 bl[189] br[189] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_190 bl[190] br[190] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_191 bl[191] br[191] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_192 bl[192] br[192] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_193 bl[193] br[193] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_194 bl[194] br[194] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_195 bl[195] br[195] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_196 bl[196] br[196] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_197 bl[197] br[197] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_198 bl[198] br[198] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_199 bl[199] br[199] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_200 bl[200] br[200] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_201 bl[201] br[201] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_202 bl[202] br[202] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_203 bl[203] br[203] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_204 bl[204] br[204] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_205 bl[205] br[205] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_206 bl[206] br[206] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_207 bl[207] br[207] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_208 bl[208] br[208] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_209 bl[209] br[209] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_210 bl[210] br[210] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_211 bl[211] br[211] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_212 bl[212] br[212] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_213 bl[213] br[213] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_214 bl[214] br[214] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_215 bl[215] br[215] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_216 bl[216] br[216] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_217 bl[217] br[217] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_218 bl[218] br[218] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_219 bl[219] br[219] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_220 bl[220] br[220] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_221 bl[221] br[221] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_222 bl[222] br[222] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_223 bl[223] br[223] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_224 bl[224] br[224] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_225 bl[225] br[225] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_226 bl[226] br[226] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_227 bl[227] br[227] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_228 bl[228] br[228] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_229 bl[229] br[229] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_230 bl[230] br[230] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_231 bl[231] br[231] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_232 bl[232] br[232] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_233 bl[233] br[233] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_234 bl[234] br[234] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_235 bl[235] br[235] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_236 bl[236] br[236] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_237 bl[237] br[237] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_238 bl[238] br[238] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_239 bl[239] br[239] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_240 bl[240] br[240] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_241 bl[241] br[241] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_242 bl[242] br[242] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_243 bl[243] br[243] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_244 bl[244] br[244] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_245 bl[245] br[245] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_246 bl[246] br[246] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_247 bl[247] br[247] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_248 bl[248] br[248] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_249 bl[249] br[249] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_250 bl[250] br[250] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_251 bl[251] br[251] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_252 bl[252] br[252] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_253 bl[253] br[253] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_254 bl[254] br[254] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_255 bl[255] br[255] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_119_0 bl[0] br[0] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_1 bl[1] br[1] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_2 bl[2] br[2] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_3 bl[3] br[3] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_4 bl[4] br[4] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_5 bl[5] br[5] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_6 bl[6] br[6] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_7 bl[7] br[7] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_8 bl[8] br[8] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_9 bl[9] br[9] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_10 bl[10] br[10] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_11 bl[11] br[11] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_12 bl[12] br[12] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_13 bl[13] br[13] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_14 bl[14] br[14] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_15 bl[15] br[15] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_16 bl[16] br[16] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_17 bl[17] br[17] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_18 bl[18] br[18] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_19 bl[19] br[19] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_20 bl[20] br[20] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_21 bl[21] br[21] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_22 bl[22] br[22] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_23 bl[23] br[23] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_24 bl[24] br[24] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_25 bl[25] br[25] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_26 bl[26] br[26] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_27 bl[27] br[27] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_28 bl[28] br[28] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_29 bl[29] br[29] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_30 bl[30] br[30] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_31 bl[31] br[31] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_32 bl[32] br[32] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_33 bl[33] br[33] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_34 bl[34] br[34] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_35 bl[35] br[35] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_36 bl[36] br[36] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_37 bl[37] br[37] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_38 bl[38] br[38] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_39 bl[39] br[39] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_40 bl[40] br[40] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_41 bl[41] br[41] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_42 bl[42] br[42] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_43 bl[43] br[43] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_44 bl[44] br[44] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_45 bl[45] br[45] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_46 bl[46] br[46] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_47 bl[47] br[47] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_48 bl[48] br[48] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_49 bl[49] br[49] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_50 bl[50] br[50] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_51 bl[51] br[51] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_52 bl[52] br[52] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_53 bl[53] br[53] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_54 bl[54] br[54] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_55 bl[55] br[55] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_56 bl[56] br[56] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_57 bl[57] br[57] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_58 bl[58] br[58] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_59 bl[59] br[59] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_60 bl[60] br[60] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_61 bl[61] br[61] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_62 bl[62] br[62] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_63 bl[63] br[63] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_64 bl[64] br[64] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_65 bl[65] br[65] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_66 bl[66] br[66] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_67 bl[67] br[67] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_68 bl[68] br[68] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_69 bl[69] br[69] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_70 bl[70] br[70] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_71 bl[71] br[71] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_72 bl[72] br[72] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_73 bl[73] br[73] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_74 bl[74] br[74] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_75 bl[75] br[75] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_76 bl[76] br[76] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_77 bl[77] br[77] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_78 bl[78] br[78] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_79 bl[79] br[79] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_80 bl[80] br[80] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_81 bl[81] br[81] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_82 bl[82] br[82] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_83 bl[83] br[83] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_84 bl[84] br[84] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_85 bl[85] br[85] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_86 bl[86] br[86] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_87 bl[87] br[87] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_88 bl[88] br[88] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_89 bl[89] br[89] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_90 bl[90] br[90] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_91 bl[91] br[91] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_92 bl[92] br[92] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_93 bl[93] br[93] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_94 bl[94] br[94] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_95 bl[95] br[95] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_96 bl[96] br[96] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_97 bl[97] br[97] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_98 bl[98] br[98] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_99 bl[99] br[99] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_100 bl[100] br[100] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_101 bl[101] br[101] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_102 bl[102] br[102] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_103 bl[103] br[103] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_104 bl[104] br[104] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_105 bl[105] br[105] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_106 bl[106] br[106] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_107 bl[107] br[107] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_108 bl[108] br[108] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_109 bl[109] br[109] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_110 bl[110] br[110] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_111 bl[111] br[111] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_112 bl[112] br[112] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_113 bl[113] br[113] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_114 bl[114] br[114] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_115 bl[115] br[115] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_116 bl[116] br[116] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_117 bl[117] br[117] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_118 bl[118] br[118] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_119 bl[119] br[119] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_120 bl[120] br[120] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_121 bl[121] br[121] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_122 bl[122] br[122] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_123 bl[123] br[123] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_124 bl[124] br[124] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_125 bl[125] br[125] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_126 bl[126] br[126] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_127 bl[127] br[127] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_128 bl[128] br[128] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_129 bl[129] br[129] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_130 bl[130] br[130] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_131 bl[131] br[131] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_132 bl[132] br[132] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_133 bl[133] br[133] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_134 bl[134] br[134] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_135 bl[135] br[135] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_136 bl[136] br[136] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_137 bl[137] br[137] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_138 bl[138] br[138] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_139 bl[139] br[139] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_140 bl[140] br[140] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_141 bl[141] br[141] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_142 bl[142] br[142] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_143 bl[143] br[143] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_144 bl[144] br[144] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_145 bl[145] br[145] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_146 bl[146] br[146] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_147 bl[147] br[147] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_148 bl[148] br[148] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_149 bl[149] br[149] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_150 bl[150] br[150] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_151 bl[151] br[151] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_152 bl[152] br[152] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_153 bl[153] br[153] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_154 bl[154] br[154] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_155 bl[155] br[155] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_156 bl[156] br[156] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_157 bl[157] br[157] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_158 bl[158] br[158] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_159 bl[159] br[159] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_160 bl[160] br[160] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_161 bl[161] br[161] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_162 bl[162] br[162] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_163 bl[163] br[163] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_164 bl[164] br[164] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_165 bl[165] br[165] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_166 bl[166] br[166] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_167 bl[167] br[167] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_168 bl[168] br[168] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_169 bl[169] br[169] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_170 bl[170] br[170] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_171 bl[171] br[171] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_172 bl[172] br[172] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_173 bl[173] br[173] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_174 bl[174] br[174] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_175 bl[175] br[175] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_176 bl[176] br[176] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_177 bl[177] br[177] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_178 bl[178] br[178] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_179 bl[179] br[179] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_180 bl[180] br[180] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_181 bl[181] br[181] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_182 bl[182] br[182] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_183 bl[183] br[183] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_184 bl[184] br[184] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_185 bl[185] br[185] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_186 bl[186] br[186] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_187 bl[187] br[187] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_188 bl[188] br[188] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_189 bl[189] br[189] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_190 bl[190] br[190] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_191 bl[191] br[191] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_192 bl[192] br[192] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_193 bl[193] br[193] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_194 bl[194] br[194] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_195 bl[195] br[195] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_196 bl[196] br[196] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_197 bl[197] br[197] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_198 bl[198] br[198] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_199 bl[199] br[199] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_200 bl[200] br[200] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_201 bl[201] br[201] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_202 bl[202] br[202] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_203 bl[203] br[203] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_204 bl[204] br[204] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_205 bl[205] br[205] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_206 bl[206] br[206] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_207 bl[207] br[207] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_208 bl[208] br[208] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_209 bl[209] br[209] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_210 bl[210] br[210] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_211 bl[211] br[211] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_212 bl[212] br[212] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_213 bl[213] br[213] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_214 bl[214] br[214] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_215 bl[215] br[215] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_216 bl[216] br[216] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_217 bl[217] br[217] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_218 bl[218] br[218] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_219 bl[219] br[219] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_220 bl[220] br[220] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_221 bl[221] br[221] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_222 bl[222] br[222] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_223 bl[223] br[223] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_224 bl[224] br[224] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_225 bl[225] br[225] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_226 bl[226] br[226] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_227 bl[227] br[227] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_228 bl[228] br[228] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_229 bl[229] br[229] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_230 bl[230] br[230] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_231 bl[231] br[231] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_232 bl[232] br[232] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_233 bl[233] br[233] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_234 bl[234] br[234] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_235 bl[235] br[235] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_236 bl[236] br[236] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_237 bl[237] br[237] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_238 bl[238] br[238] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_239 bl[239] br[239] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_240 bl[240] br[240] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_241 bl[241] br[241] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_242 bl[242] br[242] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_243 bl[243] br[243] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_244 bl[244] br[244] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_245 bl[245] br[245] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_246 bl[246] br[246] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_247 bl[247] br[247] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_248 bl[248] br[248] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_249 bl[249] br[249] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_250 bl[250] br[250] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_251 bl[251] br[251] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_252 bl[252] br[252] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_253 bl[253] br[253] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_254 bl[254] br[254] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_255 bl[255] br[255] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_120_0 bl[0] br[0] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_1 bl[1] br[1] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_2 bl[2] br[2] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_3 bl[3] br[3] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_4 bl[4] br[4] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_5 bl[5] br[5] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_6 bl[6] br[6] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_7 bl[7] br[7] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_8 bl[8] br[8] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_9 bl[9] br[9] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_10 bl[10] br[10] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_11 bl[11] br[11] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_12 bl[12] br[12] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_13 bl[13] br[13] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_14 bl[14] br[14] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_15 bl[15] br[15] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_16 bl[16] br[16] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_17 bl[17] br[17] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_18 bl[18] br[18] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_19 bl[19] br[19] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_20 bl[20] br[20] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_21 bl[21] br[21] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_22 bl[22] br[22] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_23 bl[23] br[23] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_24 bl[24] br[24] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_25 bl[25] br[25] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_26 bl[26] br[26] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_27 bl[27] br[27] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_28 bl[28] br[28] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_29 bl[29] br[29] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_30 bl[30] br[30] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_31 bl[31] br[31] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_32 bl[32] br[32] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_33 bl[33] br[33] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_34 bl[34] br[34] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_35 bl[35] br[35] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_36 bl[36] br[36] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_37 bl[37] br[37] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_38 bl[38] br[38] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_39 bl[39] br[39] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_40 bl[40] br[40] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_41 bl[41] br[41] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_42 bl[42] br[42] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_43 bl[43] br[43] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_44 bl[44] br[44] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_45 bl[45] br[45] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_46 bl[46] br[46] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_47 bl[47] br[47] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_48 bl[48] br[48] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_49 bl[49] br[49] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_50 bl[50] br[50] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_51 bl[51] br[51] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_52 bl[52] br[52] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_53 bl[53] br[53] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_54 bl[54] br[54] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_55 bl[55] br[55] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_56 bl[56] br[56] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_57 bl[57] br[57] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_58 bl[58] br[58] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_59 bl[59] br[59] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_60 bl[60] br[60] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_61 bl[61] br[61] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_62 bl[62] br[62] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_63 bl[63] br[63] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_64 bl[64] br[64] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_65 bl[65] br[65] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_66 bl[66] br[66] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_67 bl[67] br[67] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_68 bl[68] br[68] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_69 bl[69] br[69] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_70 bl[70] br[70] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_71 bl[71] br[71] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_72 bl[72] br[72] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_73 bl[73] br[73] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_74 bl[74] br[74] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_75 bl[75] br[75] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_76 bl[76] br[76] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_77 bl[77] br[77] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_78 bl[78] br[78] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_79 bl[79] br[79] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_80 bl[80] br[80] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_81 bl[81] br[81] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_82 bl[82] br[82] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_83 bl[83] br[83] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_84 bl[84] br[84] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_85 bl[85] br[85] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_86 bl[86] br[86] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_87 bl[87] br[87] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_88 bl[88] br[88] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_89 bl[89] br[89] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_90 bl[90] br[90] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_91 bl[91] br[91] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_92 bl[92] br[92] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_93 bl[93] br[93] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_94 bl[94] br[94] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_95 bl[95] br[95] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_96 bl[96] br[96] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_97 bl[97] br[97] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_98 bl[98] br[98] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_99 bl[99] br[99] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_100 bl[100] br[100] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_101 bl[101] br[101] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_102 bl[102] br[102] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_103 bl[103] br[103] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_104 bl[104] br[104] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_105 bl[105] br[105] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_106 bl[106] br[106] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_107 bl[107] br[107] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_108 bl[108] br[108] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_109 bl[109] br[109] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_110 bl[110] br[110] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_111 bl[111] br[111] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_112 bl[112] br[112] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_113 bl[113] br[113] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_114 bl[114] br[114] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_115 bl[115] br[115] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_116 bl[116] br[116] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_117 bl[117] br[117] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_118 bl[118] br[118] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_119 bl[119] br[119] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_120 bl[120] br[120] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_121 bl[121] br[121] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_122 bl[122] br[122] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_123 bl[123] br[123] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_124 bl[124] br[124] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_125 bl[125] br[125] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_126 bl[126] br[126] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_127 bl[127] br[127] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_128 bl[128] br[128] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_129 bl[129] br[129] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_130 bl[130] br[130] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_131 bl[131] br[131] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_132 bl[132] br[132] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_133 bl[133] br[133] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_134 bl[134] br[134] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_135 bl[135] br[135] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_136 bl[136] br[136] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_137 bl[137] br[137] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_138 bl[138] br[138] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_139 bl[139] br[139] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_140 bl[140] br[140] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_141 bl[141] br[141] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_142 bl[142] br[142] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_143 bl[143] br[143] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_144 bl[144] br[144] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_145 bl[145] br[145] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_146 bl[146] br[146] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_147 bl[147] br[147] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_148 bl[148] br[148] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_149 bl[149] br[149] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_150 bl[150] br[150] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_151 bl[151] br[151] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_152 bl[152] br[152] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_153 bl[153] br[153] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_154 bl[154] br[154] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_155 bl[155] br[155] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_156 bl[156] br[156] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_157 bl[157] br[157] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_158 bl[158] br[158] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_159 bl[159] br[159] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_160 bl[160] br[160] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_161 bl[161] br[161] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_162 bl[162] br[162] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_163 bl[163] br[163] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_164 bl[164] br[164] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_165 bl[165] br[165] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_166 bl[166] br[166] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_167 bl[167] br[167] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_168 bl[168] br[168] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_169 bl[169] br[169] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_170 bl[170] br[170] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_171 bl[171] br[171] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_172 bl[172] br[172] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_173 bl[173] br[173] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_174 bl[174] br[174] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_175 bl[175] br[175] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_176 bl[176] br[176] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_177 bl[177] br[177] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_178 bl[178] br[178] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_179 bl[179] br[179] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_180 bl[180] br[180] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_181 bl[181] br[181] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_182 bl[182] br[182] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_183 bl[183] br[183] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_184 bl[184] br[184] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_185 bl[185] br[185] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_186 bl[186] br[186] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_187 bl[187] br[187] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_188 bl[188] br[188] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_189 bl[189] br[189] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_190 bl[190] br[190] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_191 bl[191] br[191] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_192 bl[192] br[192] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_193 bl[193] br[193] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_194 bl[194] br[194] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_195 bl[195] br[195] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_196 bl[196] br[196] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_197 bl[197] br[197] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_198 bl[198] br[198] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_199 bl[199] br[199] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_200 bl[200] br[200] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_201 bl[201] br[201] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_202 bl[202] br[202] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_203 bl[203] br[203] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_204 bl[204] br[204] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_205 bl[205] br[205] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_206 bl[206] br[206] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_207 bl[207] br[207] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_208 bl[208] br[208] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_209 bl[209] br[209] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_210 bl[210] br[210] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_211 bl[211] br[211] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_212 bl[212] br[212] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_213 bl[213] br[213] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_214 bl[214] br[214] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_215 bl[215] br[215] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_216 bl[216] br[216] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_217 bl[217] br[217] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_218 bl[218] br[218] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_219 bl[219] br[219] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_220 bl[220] br[220] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_221 bl[221] br[221] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_222 bl[222] br[222] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_223 bl[223] br[223] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_224 bl[224] br[224] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_225 bl[225] br[225] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_226 bl[226] br[226] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_227 bl[227] br[227] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_228 bl[228] br[228] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_229 bl[229] br[229] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_230 bl[230] br[230] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_231 bl[231] br[231] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_232 bl[232] br[232] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_233 bl[233] br[233] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_234 bl[234] br[234] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_235 bl[235] br[235] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_236 bl[236] br[236] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_237 bl[237] br[237] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_238 bl[238] br[238] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_239 bl[239] br[239] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_240 bl[240] br[240] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_241 bl[241] br[241] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_242 bl[242] br[242] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_243 bl[243] br[243] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_244 bl[244] br[244] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_245 bl[245] br[245] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_246 bl[246] br[246] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_247 bl[247] br[247] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_248 bl[248] br[248] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_249 bl[249] br[249] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_250 bl[250] br[250] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_251 bl[251] br[251] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_252 bl[252] br[252] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_253 bl[253] br[253] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_254 bl[254] br[254] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_255 bl[255] br[255] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_121_0 bl[0] br[0] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_1 bl[1] br[1] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_2 bl[2] br[2] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_3 bl[3] br[3] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_4 bl[4] br[4] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_5 bl[5] br[5] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_6 bl[6] br[6] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_7 bl[7] br[7] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_8 bl[8] br[8] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_9 bl[9] br[9] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_10 bl[10] br[10] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_11 bl[11] br[11] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_12 bl[12] br[12] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_13 bl[13] br[13] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_14 bl[14] br[14] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_15 bl[15] br[15] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_16 bl[16] br[16] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_17 bl[17] br[17] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_18 bl[18] br[18] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_19 bl[19] br[19] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_20 bl[20] br[20] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_21 bl[21] br[21] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_22 bl[22] br[22] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_23 bl[23] br[23] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_24 bl[24] br[24] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_25 bl[25] br[25] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_26 bl[26] br[26] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_27 bl[27] br[27] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_28 bl[28] br[28] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_29 bl[29] br[29] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_30 bl[30] br[30] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_31 bl[31] br[31] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_32 bl[32] br[32] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_33 bl[33] br[33] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_34 bl[34] br[34] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_35 bl[35] br[35] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_36 bl[36] br[36] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_37 bl[37] br[37] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_38 bl[38] br[38] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_39 bl[39] br[39] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_40 bl[40] br[40] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_41 bl[41] br[41] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_42 bl[42] br[42] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_43 bl[43] br[43] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_44 bl[44] br[44] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_45 bl[45] br[45] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_46 bl[46] br[46] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_47 bl[47] br[47] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_48 bl[48] br[48] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_49 bl[49] br[49] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_50 bl[50] br[50] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_51 bl[51] br[51] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_52 bl[52] br[52] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_53 bl[53] br[53] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_54 bl[54] br[54] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_55 bl[55] br[55] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_56 bl[56] br[56] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_57 bl[57] br[57] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_58 bl[58] br[58] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_59 bl[59] br[59] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_60 bl[60] br[60] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_61 bl[61] br[61] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_62 bl[62] br[62] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_63 bl[63] br[63] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_64 bl[64] br[64] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_65 bl[65] br[65] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_66 bl[66] br[66] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_67 bl[67] br[67] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_68 bl[68] br[68] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_69 bl[69] br[69] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_70 bl[70] br[70] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_71 bl[71] br[71] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_72 bl[72] br[72] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_73 bl[73] br[73] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_74 bl[74] br[74] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_75 bl[75] br[75] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_76 bl[76] br[76] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_77 bl[77] br[77] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_78 bl[78] br[78] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_79 bl[79] br[79] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_80 bl[80] br[80] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_81 bl[81] br[81] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_82 bl[82] br[82] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_83 bl[83] br[83] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_84 bl[84] br[84] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_85 bl[85] br[85] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_86 bl[86] br[86] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_87 bl[87] br[87] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_88 bl[88] br[88] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_89 bl[89] br[89] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_90 bl[90] br[90] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_91 bl[91] br[91] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_92 bl[92] br[92] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_93 bl[93] br[93] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_94 bl[94] br[94] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_95 bl[95] br[95] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_96 bl[96] br[96] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_97 bl[97] br[97] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_98 bl[98] br[98] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_99 bl[99] br[99] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_100 bl[100] br[100] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_101 bl[101] br[101] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_102 bl[102] br[102] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_103 bl[103] br[103] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_104 bl[104] br[104] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_105 bl[105] br[105] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_106 bl[106] br[106] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_107 bl[107] br[107] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_108 bl[108] br[108] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_109 bl[109] br[109] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_110 bl[110] br[110] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_111 bl[111] br[111] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_112 bl[112] br[112] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_113 bl[113] br[113] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_114 bl[114] br[114] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_115 bl[115] br[115] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_116 bl[116] br[116] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_117 bl[117] br[117] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_118 bl[118] br[118] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_119 bl[119] br[119] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_120 bl[120] br[120] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_121 bl[121] br[121] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_122 bl[122] br[122] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_123 bl[123] br[123] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_124 bl[124] br[124] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_125 bl[125] br[125] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_126 bl[126] br[126] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_127 bl[127] br[127] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_128 bl[128] br[128] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_129 bl[129] br[129] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_130 bl[130] br[130] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_131 bl[131] br[131] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_132 bl[132] br[132] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_133 bl[133] br[133] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_134 bl[134] br[134] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_135 bl[135] br[135] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_136 bl[136] br[136] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_137 bl[137] br[137] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_138 bl[138] br[138] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_139 bl[139] br[139] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_140 bl[140] br[140] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_141 bl[141] br[141] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_142 bl[142] br[142] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_143 bl[143] br[143] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_144 bl[144] br[144] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_145 bl[145] br[145] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_146 bl[146] br[146] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_147 bl[147] br[147] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_148 bl[148] br[148] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_149 bl[149] br[149] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_150 bl[150] br[150] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_151 bl[151] br[151] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_152 bl[152] br[152] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_153 bl[153] br[153] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_154 bl[154] br[154] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_155 bl[155] br[155] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_156 bl[156] br[156] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_157 bl[157] br[157] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_158 bl[158] br[158] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_159 bl[159] br[159] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_160 bl[160] br[160] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_161 bl[161] br[161] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_162 bl[162] br[162] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_163 bl[163] br[163] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_164 bl[164] br[164] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_165 bl[165] br[165] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_166 bl[166] br[166] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_167 bl[167] br[167] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_168 bl[168] br[168] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_169 bl[169] br[169] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_170 bl[170] br[170] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_171 bl[171] br[171] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_172 bl[172] br[172] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_173 bl[173] br[173] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_174 bl[174] br[174] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_175 bl[175] br[175] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_176 bl[176] br[176] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_177 bl[177] br[177] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_178 bl[178] br[178] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_179 bl[179] br[179] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_180 bl[180] br[180] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_181 bl[181] br[181] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_182 bl[182] br[182] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_183 bl[183] br[183] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_184 bl[184] br[184] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_185 bl[185] br[185] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_186 bl[186] br[186] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_187 bl[187] br[187] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_188 bl[188] br[188] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_189 bl[189] br[189] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_190 bl[190] br[190] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_191 bl[191] br[191] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_192 bl[192] br[192] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_193 bl[193] br[193] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_194 bl[194] br[194] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_195 bl[195] br[195] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_196 bl[196] br[196] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_197 bl[197] br[197] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_198 bl[198] br[198] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_199 bl[199] br[199] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_200 bl[200] br[200] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_201 bl[201] br[201] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_202 bl[202] br[202] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_203 bl[203] br[203] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_204 bl[204] br[204] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_205 bl[205] br[205] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_206 bl[206] br[206] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_207 bl[207] br[207] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_208 bl[208] br[208] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_209 bl[209] br[209] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_210 bl[210] br[210] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_211 bl[211] br[211] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_212 bl[212] br[212] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_213 bl[213] br[213] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_214 bl[214] br[214] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_215 bl[215] br[215] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_216 bl[216] br[216] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_217 bl[217] br[217] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_218 bl[218] br[218] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_219 bl[219] br[219] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_220 bl[220] br[220] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_221 bl[221] br[221] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_222 bl[222] br[222] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_223 bl[223] br[223] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_224 bl[224] br[224] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_225 bl[225] br[225] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_226 bl[226] br[226] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_227 bl[227] br[227] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_228 bl[228] br[228] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_229 bl[229] br[229] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_230 bl[230] br[230] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_231 bl[231] br[231] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_232 bl[232] br[232] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_233 bl[233] br[233] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_234 bl[234] br[234] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_235 bl[235] br[235] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_236 bl[236] br[236] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_237 bl[237] br[237] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_238 bl[238] br[238] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_239 bl[239] br[239] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_240 bl[240] br[240] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_241 bl[241] br[241] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_242 bl[242] br[242] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_243 bl[243] br[243] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_244 bl[244] br[244] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_245 bl[245] br[245] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_246 bl[246] br[246] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_247 bl[247] br[247] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_248 bl[248] br[248] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_249 bl[249] br[249] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_250 bl[250] br[250] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_251 bl[251] br[251] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_252 bl[252] br[252] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_253 bl[253] br[253] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_254 bl[254] br[254] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_255 bl[255] br[255] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_122_0 bl[0] br[0] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_1 bl[1] br[1] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_2 bl[2] br[2] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_3 bl[3] br[3] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_4 bl[4] br[4] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_5 bl[5] br[5] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_6 bl[6] br[6] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_7 bl[7] br[7] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_8 bl[8] br[8] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_9 bl[9] br[9] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_10 bl[10] br[10] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_11 bl[11] br[11] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_12 bl[12] br[12] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_13 bl[13] br[13] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_14 bl[14] br[14] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_15 bl[15] br[15] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_16 bl[16] br[16] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_17 bl[17] br[17] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_18 bl[18] br[18] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_19 bl[19] br[19] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_20 bl[20] br[20] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_21 bl[21] br[21] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_22 bl[22] br[22] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_23 bl[23] br[23] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_24 bl[24] br[24] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_25 bl[25] br[25] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_26 bl[26] br[26] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_27 bl[27] br[27] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_28 bl[28] br[28] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_29 bl[29] br[29] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_30 bl[30] br[30] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_31 bl[31] br[31] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_32 bl[32] br[32] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_33 bl[33] br[33] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_34 bl[34] br[34] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_35 bl[35] br[35] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_36 bl[36] br[36] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_37 bl[37] br[37] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_38 bl[38] br[38] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_39 bl[39] br[39] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_40 bl[40] br[40] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_41 bl[41] br[41] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_42 bl[42] br[42] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_43 bl[43] br[43] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_44 bl[44] br[44] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_45 bl[45] br[45] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_46 bl[46] br[46] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_47 bl[47] br[47] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_48 bl[48] br[48] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_49 bl[49] br[49] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_50 bl[50] br[50] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_51 bl[51] br[51] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_52 bl[52] br[52] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_53 bl[53] br[53] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_54 bl[54] br[54] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_55 bl[55] br[55] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_56 bl[56] br[56] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_57 bl[57] br[57] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_58 bl[58] br[58] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_59 bl[59] br[59] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_60 bl[60] br[60] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_61 bl[61] br[61] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_62 bl[62] br[62] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_63 bl[63] br[63] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_64 bl[64] br[64] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_65 bl[65] br[65] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_66 bl[66] br[66] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_67 bl[67] br[67] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_68 bl[68] br[68] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_69 bl[69] br[69] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_70 bl[70] br[70] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_71 bl[71] br[71] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_72 bl[72] br[72] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_73 bl[73] br[73] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_74 bl[74] br[74] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_75 bl[75] br[75] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_76 bl[76] br[76] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_77 bl[77] br[77] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_78 bl[78] br[78] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_79 bl[79] br[79] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_80 bl[80] br[80] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_81 bl[81] br[81] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_82 bl[82] br[82] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_83 bl[83] br[83] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_84 bl[84] br[84] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_85 bl[85] br[85] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_86 bl[86] br[86] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_87 bl[87] br[87] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_88 bl[88] br[88] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_89 bl[89] br[89] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_90 bl[90] br[90] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_91 bl[91] br[91] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_92 bl[92] br[92] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_93 bl[93] br[93] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_94 bl[94] br[94] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_95 bl[95] br[95] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_96 bl[96] br[96] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_97 bl[97] br[97] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_98 bl[98] br[98] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_99 bl[99] br[99] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_100 bl[100] br[100] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_101 bl[101] br[101] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_102 bl[102] br[102] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_103 bl[103] br[103] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_104 bl[104] br[104] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_105 bl[105] br[105] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_106 bl[106] br[106] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_107 bl[107] br[107] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_108 bl[108] br[108] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_109 bl[109] br[109] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_110 bl[110] br[110] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_111 bl[111] br[111] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_112 bl[112] br[112] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_113 bl[113] br[113] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_114 bl[114] br[114] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_115 bl[115] br[115] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_116 bl[116] br[116] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_117 bl[117] br[117] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_118 bl[118] br[118] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_119 bl[119] br[119] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_120 bl[120] br[120] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_121 bl[121] br[121] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_122 bl[122] br[122] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_123 bl[123] br[123] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_124 bl[124] br[124] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_125 bl[125] br[125] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_126 bl[126] br[126] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_127 bl[127] br[127] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_128 bl[128] br[128] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_129 bl[129] br[129] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_130 bl[130] br[130] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_131 bl[131] br[131] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_132 bl[132] br[132] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_133 bl[133] br[133] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_134 bl[134] br[134] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_135 bl[135] br[135] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_136 bl[136] br[136] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_137 bl[137] br[137] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_138 bl[138] br[138] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_139 bl[139] br[139] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_140 bl[140] br[140] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_141 bl[141] br[141] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_142 bl[142] br[142] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_143 bl[143] br[143] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_144 bl[144] br[144] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_145 bl[145] br[145] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_146 bl[146] br[146] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_147 bl[147] br[147] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_148 bl[148] br[148] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_149 bl[149] br[149] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_150 bl[150] br[150] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_151 bl[151] br[151] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_152 bl[152] br[152] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_153 bl[153] br[153] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_154 bl[154] br[154] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_155 bl[155] br[155] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_156 bl[156] br[156] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_157 bl[157] br[157] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_158 bl[158] br[158] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_159 bl[159] br[159] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_160 bl[160] br[160] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_161 bl[161] br[161] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_162 bl[162] br[162] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_163 bl[163] br[163] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_164 bl[164] br[164] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_165 bl[165] br[165] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_166 bl[166] br[166] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_167 bl[167] br[167] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_168 bl[168] br[168] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_169 bl[169] br[169] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_170 bl[170] br[170] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_171 bl[171] br[171] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_172 bl[172] br[172] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_173 bl[173] br[173] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_174 bl[174] br[174] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_175 bl[175] br[175] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_176 bl[176] br[176] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_177 bl[177] br[177] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_178 bl[178] br[178] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_179 bl[179] br[179] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_180 bl[180] br[180] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_181 bl[181] br[181] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_182 bl[182] br[182] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_183 bl[183] br[183] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_184 bl[184] br[184] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_185 bl[185] br[185] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_186 bl[186] br[186] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_187 bl[187] br[187] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_188 bl[188] br[188] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_189 bl[189] br[189] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_190 bl[190] br[190] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_191 bl[191] br[191] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_192 bl[192] br[192] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_193 bl[193] br[193] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_194 bl[194] br[194] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_195 bl[195] br[195] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_196 bl[196] br[196] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_197 bl[197] br[197] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_198 bl[198] br[198] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_199 bl[199] br[199] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_200 bl[200] br[200] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_201 bl[201] br[201] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_202 bl[202] br[202] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_203 bl[203] br[203] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_204 bl[204] br[204] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_205 bl[205] br[205] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_206 bl[206] br[206] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_207 bl[207] br[207] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_208 bl[208] br[208] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_209 bl[209] br[209] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_210 bl[210] br[210] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_211 bl[211] br[211] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_212 bl[212] br[212] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_213 bl[213] br[213] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_214 bl[214] br[214] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_215 bl[215] br[215] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_216 bl[216] br[216] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_217 bl[217] br[217] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_218 bl[218] br[218] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_219 bl[219] br[219] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_220 bl[220] br[220] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_221 bl[221] br[221] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_222 bl[222] br[222] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_223 bl[223] br[223] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_224 bl[224] br[224] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_225 bl[225] br[225] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_226 bl[226] br[226] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_227 bl[227] br[227] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_228 bl[228] br[228] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_229 bl[229] br[229] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_230 bl[230] br[230] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_231 bl[231] br[231] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_232 bl[232] br[232] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_233 bl[233] br[233] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_234 bl[234] br[234] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_235 bl[235] br[235] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_236 bl[236] br[236] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_237 bl[237] br[237] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_238 bl[238] br[238] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_239 bl[239] br[239] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_240 bl[240] br[240] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_241 bl[241] br[241] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_242 bl[242] br[242] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_243 bl[243] br[243] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_244 bl[244] br[244] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_245 bl[245] br[245] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_246 bl[246] br[246] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_247 bl[247] br[247] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_248 bl[248] br[248] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_249 bl[249] br[249] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_250 bl[250] br[250] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_251 bl[251] br[251] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_252 bl[252] br[252] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_253 bl[253] br[253] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_254 bl[254] br[254] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_255 bl[255] br[255] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_123_0 bl[0] br[0] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_1 bl[1] br[1] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_2 bl[2] br[2] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_3 bl[3] br[3] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_4 bl[4] br[4] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_5 bl[5] br[5] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_6 bl[6] br[6] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_7 bl[7] br[7] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_8 bl[8] br[8] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_9 bl[9] br[9] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_10 bl[10] br[10] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_11 bl[11] br[11] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_12 bl[12] br[12] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_13 bl[13] br[13] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_14 bl[14] br[14] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_15 bl[15] br[15] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_16 bl[16] br[16] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_17 bl[17] br[17] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_18 bl[18] br[18] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_19 bl[19] br[19] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_20 bl[20] br[20] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_21 bl[21] br[21] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_22 bl[22] br[22] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_23 bl[23] br[23] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_24 bl[24] br[24] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_25 bl[25] br[25] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_26 bl[26] br[26] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_27 bl[27] br[27] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_28 bl[28] br[28] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_29 bl[29] br[29] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_30 bl[30] br[30] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_31 bl[31] br[31] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_32 bl[32] br[32] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_33 bl[33] br[33] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_34 bl[34] br[34] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_35 bl[35] br[35] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_36 bl[36] br[36] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_37 bl[37] br[37] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_38 bl[38] br[38] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_39 bl[39] br[39] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_40 bl[40] br[40] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_41 bl[41] br[41] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_42 bl[42] br[42] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_43 bl[43] br[43] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_44 bl[44] br[44] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_45 bl[45] br[45] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_46 bl[46] br[46] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_47 bl[47] br[47] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_48 bl[48] br[48] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_49 bl[49] br[49] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_50 bl[50] br[50] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_51 bl[51] br[51] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_52 bl[52] br[52] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_53 bl[53] br[53] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_54 bl[54] br[54] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_55 bl[55] br[55] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_56 bl[56] br[56] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_57 bl[57] br[57] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_58 bl[58] br[58] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_59 bl[59] br[59] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_60 bl[60] br[60] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_61 bl[61] br[61] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_62 bl[62] br[62] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_63 bl[63] br[63] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_64 bl[64] br[64] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_65 bl[65] br[65] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_66 bl[66] br[66] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_67 bl[67] br[67] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_68 bl[68] br[68] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_69 bl[69] br[69] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_70 bl[70] br[70] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_71 bl[71] br[71] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_72 bl[72] br[72] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_73 bl[73] br[73] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_74 bl[74] br[74] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_75 bl[75] br[75] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_76 bl[76] br[76] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_77 bl[77] br[77] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_78 bl[78] br[78] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_79 bl[79] br[79] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_80 bl[80] br[80] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_81 bl[81] br[81] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_82 bl[82] br[82] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_83 bl[83] br[83] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_84 bl[84] br[84] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_85 bl[85] br[85] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_86 bl[86] br[86] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_87 bl[87] br[87] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_88 bl[88] br[88] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_89 bl[89] br[89] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_90 bl[90] br[90] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_91 bl[91] br[91] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_92 bl[92] br[92] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_93 bl[93] br[93] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_94 bl[94] br[94] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_95 bl[95] br[95] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_96 bl[96] br[96] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_97 bl[97] br[97] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_98 bl[98] br[98] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_99 bl[99] br[99] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_100 bl[100] br[100] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_101 bl[101] br[101] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_102 bl[102] br[102] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_103 bl[103] br[103] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_104 bl[104] br[104] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_105 bl[105] br[105] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_106 bl[106] br[106] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_107 bl[107] br[107] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_108 bl[108] br[108] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_109 bl[109] br[109] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_110 bl[110] br[110] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_111 bl[111] br[111] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_112 bl[112] br[112] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_113 bl[113] br[113] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_114 bl[114] br[114] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_115 bl[115] br[115] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_116 bl[116] br[116] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_117 bl[117] br[117] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_118 bl[118] br[118] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_119 bl[119] br[119] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_120 bl[120] br[120] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_121 bl[121] br[121] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_122 bl[122] br[122] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_123 bl[123] br[123] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_124 bl[124] br[124] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_125 bl[125] br[125] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_126 bl[126] br[126] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_127 bl[127] br[127] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_128 bl[128] br[128] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_129 bl[129] br[129] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_130 bl[130] br[130] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_131 bl[131] br[131] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_132 bl[132] br[132] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_133 bl[133] br[133] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_134 bl[134] br[134] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_135 bl[135] br[135] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_136 bl[136] br[136] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_137 bl[137] br[137] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_138 bl[138] br[138] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_139 bl[139] br[139] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_140 bl[140] br[140] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_141 bl[141] br[141] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_142 bl[142] br[142] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_143 bl[143] br[143] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_144 bl[144] br[144] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_145 bl[145] br[145] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_146 bl[146] br[146] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_147 bl[147] br[147] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_148 bl[148] br[148] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_149 bl[149] br[149] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_150 bl[150] br[150] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_151 bl[151] br[151] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_152 bl[152] br[152] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_153 bl[153] br[153] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_154 bl[154] br[154] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_155 bl[155] br[155] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_156 bl[156] br[156] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_157 bl[157] br[157] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_158 bl[158] br[158] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_159 bl[159] br[159] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_160 bl[160] br[160] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_161 bl[161] br[161] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_162 bl[162] br[162] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_163 bl[163] br[163] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_164 bl[164] br[164] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_165 bl[165] br[165] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_166 bl[166] br[166] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_167 bl[167] br[167] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_168 bl[168] br[168] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_169 bl[169] br[169] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_170 bl[170] br[170] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_171 bl[171] br[171] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_172 bl[172] br[172] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_173 bl[173] br[173] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_174 bl[174] br[174] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_175 bl[175] br[175] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_176 bl[176] br[176] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_177 bl[177] br[177] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_178 bl[178] br[178] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_179 bl[179] br[179] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_180 bl[180] br[180] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_181 bl[181] br[181] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_182 bl[182] br[182] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_183 bl[183] br[183] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_184 bl[184] br[184] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_185 bl[185] br[185] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_186 bl[186] br[186] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_187 bl[187] br[187] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_188 bl[188] br[188] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_189 bl[189] br[189] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_190 bl[190] br[190] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_191 bl[191] br[191] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_192 bl[192] br[192] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_193 bl[193] br[193] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_194 bl[194] br[194] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_195 bl[195] br[195] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_196 bl[196] br[196] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_197 bl[197] br[197] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_198 bl[198] br[198] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_199 bl[199] br[199] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_200 bl[200] br[200] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_201 bl[201] br[201] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_202 bl[202] br[202] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_203 bl[203] br[203] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_204 bl[204] br[204] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_205 bl[205] br[205] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_206 bl[206] br[206] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_207 bl[207] br[207] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_208 bl[208] br[208] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_209 bl[209] br[209] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_210 bl[210] br[210] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_211 bl[211] br[211] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_212 bl[212] br[212] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_213 bl[213] br[213] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_214 bl[214] br[214] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_215 bl[215] br[215] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_216 bl[216] br[216] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_217 bl[217] br[217] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_218 bl[218] br[218] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_219 bl[219] br[219] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_220 bl[220] br[220] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_221 bl[221] br[221] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_222 bl[222] br[222] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_223 bl[223] br[223] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_224 bl[224] br[224] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_225 bl[225] br[225] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_226 bl[226] br[226] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_227 bl[227] br[227] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_228 bl[228] br[228] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_229 bl[229] br[229] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_230 bl[230] br[230] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_231 bl[231] br[231] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_232 bl[232] br[232] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_233 bl[233] br[233] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_234 bl[234] br[234] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_235 bl[235] br[235] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_236 bl[236] br[236] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_237 bl[237] br[237] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_238 bl[238] br[238] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_239 bl[239] br[239] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_240 bl[240] br[240] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_241 bl[241] br[241] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_242 bl[242] br[242] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_243 bl[243] br[243] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_244 bl[244] br[244] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_245 bl[245] br[245] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_246 bl[246] br[246] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_247 bl[247] br[247] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_248 bl[248] br[248] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_249 bl[249] br[249] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_250 bl[250] br[250] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_251 bl[251] br[251] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_252 bl[252] br[252] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_253 bl[253] br[253] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_254 bl[254] br[254] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_255 bl[255] br[255] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_124_0 bl[0] br[0] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_1 bl[1] br[1] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_2 bl[2] br[2] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_3 bl[3] br[3] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_4 bl[4] br[4] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_5 bl[5] br[5] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_6 bl[6] br[6] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_7 bl[7] br[7] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_8 bl[8] br[8] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_9 bl[9] br[9] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_10 bl[10] br[10] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_11 bl[11] br[11] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_12 bl[12] br[12] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_13 bl[13] br[13] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_14 bl[14] br[14] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_15 bl[15] br[15] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_16 bl[16] br[16] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_17 bl[17] br[17] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_18 bl[18] br[18] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_19 bl[19] br[19] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_20 bl[20] br[20] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_21 bl[21] br[21] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_22 bl[22] br[22] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_23 bl[23] br[23] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_24 bl[24] br[24] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_25 bl[25] br[25] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_26 bl[26] br[26] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_27 bl[27] br[27] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_28 bl[28] br[28] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_29 bl[29] br[29] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_30 bl[30] br[30] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_31 bl[31] br[31] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_32 bl[32] br[32] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_33 bl[33] br[33] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_34 bl[34] br[34] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_35 bl[35] br[35] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_36 bl[36] br[36] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_37 bl[37] br[37] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_38 bl[38] br[38] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_39 bl[39] br[39] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_40 bl[40] br[40] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_41 bl[41] br[41] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_42 bl[42] br[42] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_43 bl[43] br[43] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_44 bl[44] br[44] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_45 bl[45] br[45] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_46 bl[46] br[46] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_47 bl[47] br[47] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_48 bl[48] br[48] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_49 bl[49] br[49] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_50 bl[50] br[50] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_51 bl[51] br[51] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_52 bl[52] br[52] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_53 bl[53] br[53] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_54 bl[54] br[54] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_55 bl[55] br[55] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_56 bl[56] br[56] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_57 bl[57] br[57] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_58 bl[58] br[58] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_59 bl[59] br[59] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_60 bl[60] br[60] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_61 bl[61] br[61] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_62 bl[62] br[62] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_63 bl[63] br[63] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_64 bl[64] br[64] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_65 bl[65] br[65] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_66 bl[66] br[66] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_67 bl[67] br[67] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_68 bl[68] br[68] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_69 bl[69] br[69] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_70 bl[70] br[70] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_71 bl[71] br[71] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_72 bl[72] br[72] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_73 bl[73] br[73] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_74 bl[74] br[74] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_75 bl[75] br[75] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_76 bl[76] br[76] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_77 bl[77] br[77] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_78 bl[78] br[78] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_79 bl[79] br[79] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_80 bl[80] br[80] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_81 bl[81] br[81] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_82 bl[82] br[82] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_83 bl[83] br[83] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_84 bl[84] br[84] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_85 bl[85] br[85] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_86 bl[86] br[86] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_87 bl[87] br[87] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_88 bl[88] br[88] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_89 bl[89] br[89] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_90 bl[90] br[90] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_91 bl[91] br[91] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_92 bl[92] br[92] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_93 bl[93] br[93] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_94 bl[94] br[94] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_95 bl[95] br[95] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_96 bl[96] br[96] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_97 bl[97] br[97] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_98 bl[98] br[98] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_99 bl[99] br[99] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_100 bl[100] br[100] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_101 bl[101] br[101] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_102 bl[102] br[102] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_103 bl[103] br[103] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_104 bl[104] br[104] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_105 bl[105] br[105] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_106 bl[106] br[106] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_107 bl[107] br[107] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_108 bl[108] br[108] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_109 bl[109] br[109] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_110 bl[110] br[110] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_111 bl[111] br[111] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_112 bl[112] br[112] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_113 bl[113] br[113] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_114 bl[114] br[114] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_115 bl[115] br[115] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_116 bl[116] br[116] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_117 bl[117] br[117] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_118 bl[118] br[118] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_119 bl[119] br[119] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_120 bl[120] br[120] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_121 bl[121] br[121] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_122 bl[122] br[122] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_123 bl[123] br[123] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_124 bl[124] br[124] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_125 bl[125] br[125] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_126 bl[126] br[126] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_127 bl[127] br[127] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_128 bl[128] br[128] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_129 bl[129] br[129] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_130 bl[130] br[130] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_131 bl[131] br[131] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_132 bl[132] br[132] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_133 bl[133] br[133] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_134 bl[134] br[134] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_135 bl[135] br[135] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_136 bl[136] br[136] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_137 bl[137] br[137] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_138 bl[138] br[138] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_139 bl[139] br[139] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_140 bl[140] br[140] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_141 bl[141] br[141] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_142 bl[142] br[142] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_143 bl[143] br[143] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_144 bl[144] br[144] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_145 bl[145] br[145] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_146 bl[146] br[146] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_147 bl[147] br[147] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_148 bl[148] br[148] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_149 bl[149] br[149] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_150 bl[150] br[150] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_151 bl[151] br[151] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_152 bl[152] br[152] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_153 bl[153] br[153] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_154 bl[154] br[154] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_155 bl[155] br[155] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_156 bl[156] br[156] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_157 bl[157] br[157] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_158 bl[158] br[158] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_159 bl[159] br[159] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_160 bl[160] br[160] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_161 bl[161] br[161] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_162 bl[162] br[162] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_163 bl[163] br[163] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_164 bl[164] br[164] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_165 bl[165] br[165] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_166 bl[166] br[166] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_167 bl[167] br[167] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_168 bl[168] br[168] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_169 bl[169] br[169] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_170 bl[170] br[170] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_171 bl[171] br[171] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_172 bl[172] br[172] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_173 bl[173] br[173] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_174 bl[174] br[174] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_175 bl[175] br[175] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_176 bl[176] br[176] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_177 bl[177] br[177] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_178 bl[178] br[178] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_179 bl[179] br[179] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_180 bl[180] br[180] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_181 bl[181] br[181] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_182 bl[182] br[182] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_183 bl[183] br[183] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_184 bl[184] br[184] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_185 bl[185] br[185] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_186 bl[186] br[186] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_187 bl[187] br[187] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_188 bl[188] br[188] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_189 bl[189] br[189] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_190 bl[190] br[190] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_191 bl[191] br[191] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_192 bl[192] br[192] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_193 bl[193] br[193] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_194 bl[194] br[194] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_195 bl[195] br[195] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_196 bl[196] br[196] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_197 bl[197] br[197] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_198 bl[198] br[198] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_199 bl[199] br[199] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_200 bl[200] br[200] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_201 bl[201] br[201] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_202 bl[202] br[202] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_203 bl[203] br[203] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_204 bl[204] br[204] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_205 bl[205] br[205] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_206 bl[206] br[206] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_207 bl[207] br[207] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_208 bl[208] br[208] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_209 bl[209] br[209] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_210 bl[210] br[210] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_211 bl[211] br[211] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_212 bl[212] br[212] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_213 bl[213] br[213] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_214 bl[214] br[214] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_215 bl[215] br[215] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_216 bl[216] br[216] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_217 bl[217] br[217] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_218 bl[218] br[218] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_219 bl[219] br[219] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_220 bl[220] br[220] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_221 bl[221] br[221] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_222 bl[222] br[222] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_223 bl[223] br[223] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_224 bl[224] br[224] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_225 bl[225] br[225] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_226 bl[226] br[226] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_227 bl[227] br[227] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_228 bl[228] br[228] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_229 bl[229] br[229] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_230 bl[230] br[230] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_231 bl[231] br[231] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_232 bl[232] br[232] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_233 bl[233] br[233] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_234 bl[234] br[234] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_235 bl[235] br[235] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_236 bl[236] br[236] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_237 bl[237] br[237] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_238 bl[238] br[238] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_239 bl[239] br[239] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_240 bl[240] br[240] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_241 bl[241] br[241] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_242 bl[242] br[242] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_243 bl[243] br[243] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_244 bl[244] br[244] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_245 bl[245] br[245] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_246 bl[246] br[246] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_247 bl[247] br[247] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_248 bl[248] br[248] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_249 bl[249] br[249] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_250 bl[250] br[250] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_251 bl[251] br[251] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_252 bl[252] br[252] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_253 bl[253] br[253] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_254 bl[254] br[254] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_255 bl[255] br[255] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_125_0 bl[0] br[0] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_1 bl[1] br[1] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_2 bl[2] br[2] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_3 bl[3] br[3] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_4 bl[4] br[4] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_5 bl[5] br[5] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_6 bl[6] br[6] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_7 bl[7] br[7] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_8 bl[8] br[8] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_9 bl[9] br[9] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_10 bl[10] br[10] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_11 bl[11] br[11] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_12 bl[12] br[12] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_13 bl[13] br[13] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_14 bl[14] br[14] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_15 bl[15] br[15] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_16 bl[16] br[16] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_17 bl[17] br[17] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_18 bl[18] br[18] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_19 bl[19] br[19] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_20 bl[20] br[20] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_21 bl[21] br[21] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_22 bl[22] br[22] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_23 bl[23] br[23] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_24 bl[24] br[24] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_25 bl[25] br[25] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_26 bl[26] br[26] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_27 bl[27] br[27] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_28 bl[28] br[28] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_29 bl[29] br[29] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_30 bl[30] br[30] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_31 bl[31] br[31] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_32 bl[32] br[32] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_33 bl[33] br[33] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_34 bl[34] br[34] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_35 bl[35] br[35] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_36 bl[36] br[36] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_37 bl[37] br[37] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_38 bl[38] br[38] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_39 bl[39] br[39] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_40 bl[40] br[40] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_41 bl[41] br[41] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_42 bl[42] br[42] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_43 bl[43] br[43] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_44 bl[44] br[44] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_45 bl[45] br[45] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_46 bl[46] br[46] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_47 bl[47] br[47] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_48 bl[48] br[48] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_49 bl[49] br[49] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_50 bl[50] br[50] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_51 bl[51] br[51] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_52 bl[52] br[52] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_53 bl[53] br[53] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_54 bl[54] br[54] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_55 bl[55] br[55] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_56 bl[56] br[56] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_57 bl[57] br[57] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_58 bl[58] br[58] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_59 bl[59] br[59] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_60 bl[60] br[60] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_61 bl[61] br[61] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_62 bl[62] br[62] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_63 bl[63] br[63] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_64 bl[64] br[64] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_65 bl[65] br[65] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_66 bl[66] br[66] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_67 bl[67] br[67] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_68 bl[68] br[68] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_69 bl[69] br[69] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_70 bl[70] br[70] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_71 bl[71] br[71] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_72 bl[72] br[72] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_73 bl[73] br[73] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_74 bl[74] br[74] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_75 bl[75] br[75] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_76 bl[76] br[76] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_77 bl[77] br[77] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_78 bl[78] br[78] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_79 bl[79] br[79] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_80 bl[80] br[80] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_81 bl[81] br[81] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_82 bl[82] br[82] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_83 bl[83] br[83] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_84 bl[84] br[84] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_85 bl[85] br[85] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_86 bl[86] br[86] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_87 bl[87] br[87] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_88 bl[88] br[88] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_89 bl[89] br[89] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_90 bl[90] br[90] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_91 bl[91] br[91] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_92 bl[92] br[92] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_93 bl[93] br[93] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_94 bl[94] br[94] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_95 bl[95] br[95] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_96 bl[96] br[96] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_97 bl[97] br[97] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_98 bl[98] br[98] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_99 bl[99] br[99] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_100 bl[100] br[100] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_101 bl[101] br[101] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_102 bl[102] br[102] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_103 bl[103] br[103] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_104 bl[104] br[104] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_105 bl[105] br[105] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_106 bl[106] br[106] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_107 bl[107] br[107] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_108 bl[108] br[108] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_109 bl[109] br[109] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_110 bl[110] br[110] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_111 bl[111] br[111] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_112 bl[112] br[112] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_113 bl[113] br[113] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_114 bl[114] br[114] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_115 bl[115] br[115] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_116 bl[116] br[116] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_117 bl[117] br[117] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_118 bl[118] br[118] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_119 bl[119] br[119] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_120 bl[120] br[120] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_121 bl[121] br[121] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_122 bl[122] br[122] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_123 bl[123] br[123] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_124 bl[124] br[124] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_125 bl[125] br[125] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_126 bl[126] br[126] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_127 bl[127] br[127] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_128 bl[128] br[128] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_129 bl[129] br[129] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_130 bl[130] br[130] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_131 bl[131] br[131] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_132 bl[132] br[132] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_133 bl[133] br[133] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_134 bl[134] br[134] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_135 bl[135] br[135] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_136 bl[136] br[136] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_137 bl[137] br[137] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_138 bl[138] br[138] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_139 bl[139] br[139] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_140 bl[140] br[140] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_141 bl[141] br[141] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_142 bl[142] br[142] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_143 bl[143] br[143] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_144 bl[144] br[144] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_145 bl[145] br[145] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_146 bl[146] br[146] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_147 bl[147] br[147] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_148 bl[148] br[148] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_149 bl[149] br[149] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_150 bl[150] br[150] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_151 bl[151] br[151] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_152 bl[152] br[152] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_153 bl[153] br[153] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_154 bl[154] br[154] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_155 bl[155] br[155] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_156 bl[156] br[156] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_157 bl[157] br[157] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_158 bl[158] br[158] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_159 bl[159] br[159] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_160 bl[160] br[160] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_161 bl[161] br[161] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_162 bl[162] br[162] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_163 bl[163] br[163] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_164 bl[164] br[164] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_165 bl[165] br[165] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_166 bl[166] br[166] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_167 bl[167] br[167] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_168 bl[168] br[168] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_169 bl[169] br[169] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_170 bl[170] br[170] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_171 bl[171] br[171] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_172 bl[172] br[172] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_173 bl[173] br[173] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_174 bl[174] br[174] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_175 bl[175] br[175] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_176 bl[176] br[176] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_177 bl[177] br[177] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_178 bl[178] br[178] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_179 bl[179] br[179] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_180 bl[180] br[180] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_181 bl[181] br[181] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_182 bl[182] br[182] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_183 bl[183] br[183] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_184 bl[184] br[184] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_185 bl[185] br[185] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_186 bl[186] br[186] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_187 bl[187] br[187] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_188 bl[188] br[188] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_189 bl[189] br[189] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_190 bl[190] br[190] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_191 bl[191] br[191] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_192 bl[192] br[192] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_193 bl[193] br[193] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_194 bl[194] br[194] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_195 bl[195] br[195] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_196 bl[196] br[196] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_197 bl[197] br[197] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_198 bl[198] br[198] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_199 bl[199] br[199] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_200 bl[200] br[200] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_201 bl[201] br[201] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_202 bl[202] br[202] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_203 bl[203] br[203] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_204 bl[204] br[204] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_205 bl[205] br[205] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_206 bl[206] br[206] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_207 bl[207] br[207] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_208 bl[208] br[208] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_209 bl[209] br[209] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_210 bl[210] br[210] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_211 bl[211] br[211] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_212 bl[212] br[212] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_213 bl[213] br[213] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_214 bl[214] br[214] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_215 bl[215] br[215] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_216 bl[216] br[216] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_217 bl[217] br[217] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_218 bl[218] br[218] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_219 bl[219] br[219] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_220 bl[220] br[220] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_221 bl[221] br[221] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_222 bl[222] br[222] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_223 bl[223] br[223] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_224 bl[224] br[224] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_225 bl[225] br[225] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_226 bl[226] br[226] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_227 bl[227] br[227] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_228 bl[228] br[228] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_229 bl[229] br[229] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_230 bl[230] br[230] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_231 bl[231] br[231] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_232 bl[232] br[232] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_233 bl[233] br[233] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_234 bl[234] br[234] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_235 bl[235] br[235] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_236 bl[236] br[236] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_237 bl[237] br[237] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_238 bl[238] br[238] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_239 bl[239] br[239] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_240 bl[240] br[240] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_241 bl[241] br[241] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_242 bl[242] br[242] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_243 bl[243] br[243] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_244 bl[244] br[244] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_245 bl[245] br[245] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_246 bl[246] br[246] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_247 bl[247] br[247] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_248 bl[248] br[248] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_249 bl[249] br[249] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_250 bl[250] br[250] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_251 bl[251] br[251] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_252 bl[252] br[252] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_253 bl[253] br[253] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_254 bl[254] br[254] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_255 bl[255] br[255] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_126_0 bl[0] br[0] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_1 bl[1] br[1] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_2 bl[2] br[2] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_3 bl[3] br[3] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_4 bl[4] br[4] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_5 bl[5] br[5] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_6 bl[6] br[6] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_7 bl[7] br[7] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_8 bl[8] br[8] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_9 bl[9] br[9] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_10 bl[10] br[10] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_11 bl[11] br[11] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_12 bl[12] br[12] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_13 bl[13] br[13] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_14 bl[14] br[14] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_15 bl[15] br[15] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_16 bl[16] br[16] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_17 bl[17] br[17] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_18 bl[18] br[18] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_19 bl[19] br[19] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_20 bl[20] br[20] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_21 bl[21] br[21] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_22 bl[22] br[22] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_23 bl[23] br[23] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_24 bl[24] br[24] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_25 bl[25] br[25] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_26 bl[26] br[26] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_27 bl[27] br[27] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_28 bl[28] br[28] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_29 bl[29] br[29] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_30 bl[30] br[30] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_31 bl[31] br[31] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_32 bl[32] br[32] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_33 bl[33] br[33] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_34 bl[34] br[34] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_35 bl[35] br[35] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_36 bl[36] br[36] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_37 bl[37] br[37] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_38 bl[38] br[38] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_39 bl[39] br[39] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_40 bl[40] br[40] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_41 bl[41] br[41] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_42 bl[42] br[42] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_43 bl[43] br[43] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_44 bl[44] br[44] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_45 bl[45] br[45] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_46 bl[46] br[46] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_47 bl[47] br[47] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_48 bl[48] br[48] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_49 bl[49] br[49] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_50 bl[50] br[50] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_51 bl[51] br[51] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_52 bl[52] br[52] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_53 bl[53] br[53] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_54 bl[54] br[54] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_55 bl[55] br[55] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_56 bl[56] br[56] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_57 bl[57] br[57] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_58 bl[58] br[58] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_59 bl[59] br[59] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_60 bl[60] br[60] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_61 bl[61] br[61] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_62 bl[62] br[62] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_63 bl[63] br[63] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_64 bl[64] br[64] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_65 bl[65] br[65] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_66 bl[66] br[66] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_67 bl[67] br[67] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_68 bl[68] br[68] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_69 bl[69] br[69] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_70 bl[70] br[70] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_71 bl[71] br[71] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_72 bl[72] br[72] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_73 bl[73] br[73] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_74 bl[74] br[74] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_75 bl[75] br[75] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_76 bl[76] br[76] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_77 bl[77] br[77] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_78 bl[78] br[78] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_79 bl[79] br[79] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_80 bl[80] br[80] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_81 bl[81] br[81] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_82 bl[82] br[82] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_83 bl[83] br[83] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_84 bl[84] br[84] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_85 bl[85] br[85] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_86 bl[86] br[86] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_87 bl[87] br[87] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_88 bl[88] br[88] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_89 bl[89] br[89] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_90 bl[90] br[90] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_91 bl[91] br[91] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_92 bl[92] br[92] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_93 bl[93] br[93] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_94 bl[94] br[94] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_95 bl[95] br[95] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_96 bl[96] br[96] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_97 bl[97] br[97] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_98 bl[98] br[98] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_99 bl[99] br[99] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_100 bl[100] br[100] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_101 bl[101] br[101] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_102 bl[102] br[102] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_103 bl[103] br[103] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_104 bl[104] br[104] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_105 bl[105] br[105] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_106 bl[106] br[106] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_107 bl[107] br[107] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_108 bl[108] br[108] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_109 bl[109] br[109] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_110 bl[110] br[110] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_111 bl[111] br[111] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_112 bl[112] br[112] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_113 bl[113] br[113] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_114 bl[114] br[114] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_115 bl[115] br[115] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_116 bl[116] br[116] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_117 bl[117] br[117] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_118 bl[118] br[118] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_119 bl[119] br[119] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_120 bl[120] br[120] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_121 bl[121] br[121] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_122 bl[122] br[122] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_123 bl[123] br[123] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_124 bl[124] br[124] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_125 bl[125] br[125] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_126 bl[126] br[126] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_127 bl[127] br[127] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_128 bl[128] br[128] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_129 bl[129] br[129] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_130 bl[130] br[130] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_131 bl[131] br[131] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_132 bl[132] br[132] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_133 bl[133] br[133] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_134 bl[134] br[134] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_135 bl[135] br[135] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_136 bl[136] br[136] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_137 bl[137] br[137] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_138 bl[138] br[138] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_139 bl[139] br[139] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_140 bl[140] br[140] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_141 bl[141] br[141] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_142 bl[142] br[142] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_143 bl[143] br[143] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_144 bl[144] br[144] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_145 bl[145] br[145] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_146 bl[146] br[146] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_147 bl[147] br[147] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_148 bl[148] br[148] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_149 bl[149] br[149] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_150 bl[150] br[150] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_151 bl[151] br[151] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_152 bl[152] br[152] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_153 bl[153] br[153] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_154 bl[154] br[154] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_155 bl[155] br[155] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_156 bl[156] br[156] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_157 bl[157] br[157] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_158 bl[158] br[158] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_159 bl[159] br[159] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_160 bl[160] br[160] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_161 bl[161] br[161] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_162 bl[162] br[162] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_163 bl[163] br[163] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_164 bl[164] br[164] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_165 bl[165] br[165] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_166 bl[166] br[166] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_167 bl[167] br[167] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_168 bl[168] br[168] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_169 bl[169] br[169] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_170 bl[170] br[170] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_171 bl[171] br[171] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_172 bl[172] br[172] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_173 bl[173] br[173] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_174 bl[174] br[174] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_175 bl[175] br[175] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_176 bl[176] br[176] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_177 bl[177] br[177] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_178 bl[178] br[178] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_179 bl[179] br[179] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_180 bl[180] br[180] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_181 bl[181] br[181] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_182 bl[182] br[182] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_183 bl[183] br[183] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_184 bl[184] br[184] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_185 bl[185] br[185] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_186 bl[186] br[186] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_187 bl[187] br[187] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_188 bl[188] br[188] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_189 bl[189] br[189] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_190 bl[190] br[190] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_191 bl[191] br[191] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_192 bl[192] br[192] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_193 bl[193] br[193] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_194 bl[194] br[194] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_195 bl[195] br[195] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_196 bl[196] br[196] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_197 bl[197] br[197] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_198 bl[198] br[198] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_199 bl[199] br[199] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_200 bl[200] br[200] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_201 bl[201] br[201] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_202 bl[202] br[202] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_203 bl[203] br[203] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_204 bl[204] br[204] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_205 bl[205] br[205] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_206 bl[206] br[206] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_207 bl[207] br[207] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_208 bl[208] br[208] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_209 bl[209] br[209] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_210 bl[210] br[210] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_211 bl[211] br[211] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_212 bl[212] br[212] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_213 bl[213] br[213] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_214 bl[214] br[214] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_215 bl[215] br[215] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_216 bl[216] br[216] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_217 bl[217] br[217] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_218 bl[218] br[218] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_219 bl[219] br[219] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_220 bl[220] br[220] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_221 bl[221] br[221] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_222 bl[222] br[222] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_223 bl[223] br[223] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_224 bl[224] br[224] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_225 bl[225] br[225] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_226 bl[226] br[226] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_227 bl[227] br[227] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_228 bl[228] br[228] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_229 bl[229] br[229] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_230 bl[230] br[230] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_231 bl[231] br[231] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_232 bl[232] br[232] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_233 bl[233] br[233] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_234 bl[234] br[234] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_235 bl[235] br[235] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_236 bl[236] br[236] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_237 bl[237] br[237] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_238 bl[238] br[238] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_239 bl[239] br[239] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_240 bl[240] br[240] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_241 bl[241] br[241] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_242 bl[242] br[242] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_243 bl[243] br[243] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_244 bl[244] br[244] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_245 bl[245] br[245] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_246 bl[246] br[246] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_247 bl[247] br[247] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_248 bl[248] br[248] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_249 bl[249] br[249] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_250 bl[250] br[250] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_251 bl[251] br[251] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_252 bl[252] br[252] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_253 bl[253] br[253] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_254 bl[254] br[254] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_255 bl[255] br[255] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_127_0 bl[0] br[0] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_1 bl[1] br[1] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_2 bl[2] br[2] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_3 bl[3] br[3] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_4 bl[4] br[4] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_5 bl[5] br[5] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_6 bl[6] br[6] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_7 bl[7] br[7] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_8 bl[8] br[8] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_9 bl[9] br[9] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_10 bl[10] br[10] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_11 bl[11] br[11] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_12 bl[12] br[12] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_13 bl[13] br[13] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_14 bl[14] br[14] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_15 bl[15] br[15] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_16 bl[16] br[16] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_17 bl[17] br[17] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_18 bl[18] br[18] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_19 bl[19] br[19] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_20 bl[20] br[20] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_21 bl[21] br[21] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_22 bl[22] br[22] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_23 bl[23] br[23] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_24 bl[24] br[24] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_25 bl[25] br[25] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_26 bl[26] br[26] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_27 bl[27] br[27] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_28 bl[28] br[28] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_29 bl[29] br[29] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_30 bl[30] br[30] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_31 bl[31] br[31] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_32 bl[32] br[32] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_33 bl[33] br[33] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_34 bl[34] br[34] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_35 bl[35] br[35] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_36 bl[36] br[36] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_37 bl[37] br[37] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_38 bl[38] br[38] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_39 bl[39] br[39] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_40 bl[40] br[40] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_41 bl[41] br[41] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_42 bl[42] br[42] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_43 bl[43] br[43] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_44 bl[44] br[44] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_45 bl[45] br[45] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_46 bl[46] br[46] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_47 bl[47] br[47] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_48 bl[48] br[48] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_49 bl[49] br[49] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_50 bl[50] br[50] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_51 bl[51] br[51] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_52 bl[52] br[52] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_53 bl[53] br[53] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_54 bl[54] br[54] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_55 bl[55] br[55] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_56 bl[56] br[56] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_57 bl[57] br[57] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_58 bl[58] br[58] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_59 bl[59] br[59] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_60 bl[60] br[60] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_61 bl[61] br[61] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_62 bl[62] br[62] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_63 bl[63] br[63] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_64 bl[64] br[64] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_65 bl[65] br[65] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_66 bl[66] br[66] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_67 bl[67] br[67] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_68 bl[68] br[68] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_69 bl[69] br[69] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_70 bl[70] br[70] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_71 bl[71] br[71] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_72 bl[72] br[72] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_73 bl[73] br[73] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_74 bl[74] br[74] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_75 bl[75] br[75] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_76 bl[76] br[76] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_77 bl[77] br[77] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_78 bl[78] br[78] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_79 bl[79] br[79] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_80 bl[80] br[80] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_81 bl[81] br[81] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_82 bl[82] br[82] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_83 bl[83] br[83] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_84 bl[84] br[84] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_85 bl[85] br[85] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_86 bl[86] br[86] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_87 bl[87] br[87] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_88 bl[88] br[88] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_89 bl[89] br[89] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_90 bl[90] br[90] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_91 bl[91] br[91] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_92 bl[92] br[92] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_93 bl[93] br[93] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_94 bl[94] br[94] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_95 bl[95] br[95] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_96 bl[96] br[96] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_97 bl[97] br[97] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_98 bl[98] br[98] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_99 bl[99] br[99] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_100 bl[100] br[100] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_101 bl[101] br[101] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_102 bl[102] br[102] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_103 bl[103] br[103] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_104 bl[104] br[104] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_105 bl[105] br[105] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_106 bl[106] br[106] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_107 bl[107] br[107] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_108 bl[108] br[108] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_109 bl[109] br[109] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_110 bl[110] br[110] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_111 bl[111] br[111] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_112 bl[112] br[112] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_113 bl[113] br[113] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_114 bl[114] br[114] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_115 bl[115] br[115] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_116 bl[116] br[116] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_117 bl[117] br[117] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_118 bl[118] br[118] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_119 bl[119] br[119] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_120 bl[120] br[120] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_121 bl[121] br[121] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_122 bl[122] br[122] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_123 bl[123] br[123] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_124 bl[124] br[124] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_125 bl[125] br[125] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_126 bl[126] br[126] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_127 bl[127] br[127] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_128 bl[128] br[128] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_129 bl[129] br[129] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_130 bl[130] br[130] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_131 bl[131] br[131] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_132 bl[132] br[132] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_133 bl[133] br[133] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_134 bl[134] br[134] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_135 bl[135] br[135] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_136 bl[136] br[136] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_137 bl[137] br[137] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_138 bl[138] br[138] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_139 bl[139] br[139] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_140 bl[140] br[140] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_141 bl[141] br[141] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_142 bl[142] br[142] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_143 bl[143] br[143] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_144 bl[144] br[144] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_145 bl[145] br[145] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_146 bl[146] br[146] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_147 bl[147] br[147] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_148 bl[148] br[148] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_149 bl[149] br[149] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_150 bl[150] br[150] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_151 bl[151] br[151] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_152 bl[152] br[152] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_153 bl[153] br[153] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_154 bl[154] br[154] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_155 bl[155] br[155] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_156 bl[156] br[156] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_157 bl[157] br[157] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_158 bl[158] br[158] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_159 bl[159] br[159] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_160 bl[160] br[160] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_161 bl[161] br[161] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_162 bl[162] br[162] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_163 bl[163] br[163] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_164 bl[164] br[164] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_165 bl[165] br[165] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_166 bl[166] br[166] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_167 bl[167] br[167] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_168 bl[168] br[168] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_169 bl[169] br[169] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_170 bl[170] br[170] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_171 bl[171] br[171] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_172 bl[172] br[172] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_173 bl[173] br[173] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_174 bl[174] br[174] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_175 bl[175] br[175] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_176 bl[176] br[176] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_177 bl[177] br[177] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_178 bl[178] br[178] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_179 bl[179] br[179] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_180 bl[180] br[180] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_181 bl[181] br[181] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_182 bl[182] br[182] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_183 bl[183] br[183] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_184 bl[184] br[184] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_185 bl[185] br[185] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_186 bl[186] br[186] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_187 bl[187] br[187] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_188 bl[188] br[188] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_189 bl[189] br[189] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_190 bl[190] br[190] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_191 bl[191] br[191] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_192 bl[192] br[192] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_193 bl[193] br[193] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_194 bl[194] br[194] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_195 bl[195] br[195] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_196 bl[196] br[196] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_197 bl[197] br[197] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_198 bl[198] br[198] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_199 bl[199] br[199] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_200 bl[200] br[200] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_201 bl[201] br[201] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_202 bl[202] br[202] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_203 bl[203] br[203] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_204 bl[204] br[204] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_205 bl[205] br[205] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_206 bl[206] br[206] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_207 bl[207] br[207] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_208 bl[208] br[208] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_209 bl[209] br[209] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_210 bl[210] br[210] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_211 bl[211] br[211] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_212 bl[212] br[212] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_213 bl[213] br[213] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_214 bl[214] br[214] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_215 bl[215] br[215] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_216 bl[216] br[216] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_217 bl[217] br[217] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_218 bl[218] br[218] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_219 bl[219] br[219] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_220 bl[220] br[220] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_221 bl[221] br[221] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_222 bl[222] br[222] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_223 bl[223] br[223] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_224 bl[224] br[224] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_225 bl[225] br[225] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_226 bl[226] br[226] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_227 bl[227] br[227] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_228 bl[228] br[228] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_229 bl[229] br[229] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_230 bl[230] br[230] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_231 bl[231] br[231] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_232 bl[232] br[232] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_233 bl[233] br[233] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_234 bl[234] br[234] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_235 bl[235] br[235] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_236 bl[236] br[236] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_237 bl[237] br[237] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_238 bl[238] br[238] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_239 bl[239] br[239] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_240 bl[240] br[240] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_241 bl[241] br[241] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_242 bl[242] br[242] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_243 bl[243] br[243] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_244 bl[244] br[244] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_245 bl[245] br[245] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_246 bl[246] br[246] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_247 bl[247] br[247] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_248 bl[248] br[248] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_249 bl[249] br[249] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_250 bl[250] br[250] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_251 bl[251] br[251] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_252 bl[252] br[252] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_253 bl[253] br[253] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_254 bl[254] br[254] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_255 bl[255] br[255] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_0 dummy_bl dummy_br vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_0 vdd vdd vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_1 dummy_bl dummy_br vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_1 vdd vdd vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_2 dummy_bl dummy_br vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_2 vdd vdd vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_3 dummy_bl dummy_br vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_3 vdd vdd vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_4 dummy_bl dummy_br vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_4 vdd vdd vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_5 dummy_bl dummy_br vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_5 vdd vdd vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_6 dummy_bl dummy_br vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_6 vdd vdd vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_7 dummy_bl dummy_br vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_7 vdd vdd vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_8 dummy_bl dummy_br vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_8 vdd vdd vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_9 dummy_bl dummy_br vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_9 vdd vdd vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_10 dummy_bl dummy_br vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_10 vdd vdd vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_11 dummy_bl dummy_br vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_11 vdd vdd vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_12 dummy_bl dummy_br vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_12 vdd vdd vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_13 dummy_bl dummy_br vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_13 vdd vdd vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_14 dummy_bl dummy_br vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_14 vdd vdd vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_15 dummy_bl dummy_br vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_15 vdd vdd vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_16 dummy_bl dummy_br vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_16 vdd vdd vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_17 dummy_bl dummy_br vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_17 vdd vdd vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_18 dummy_bl dummy_br vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_18 vdd vdd vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_19 dummy_bl dummy_br vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_19 vdd vdd vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_20 dummy_bl dummy_br vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_20 vdd vdd vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_21 dummy_bl dummy_br vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_21 vdd vdd vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_22 dummy_bl dummy_br vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_22 vdd vdd vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_23 dummy_bl dummy_br vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_23 vdd vdd vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_24 dummy_bl dummy_br vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_24 vdd vdd vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_25 dummy_bl dummy_br vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_25 vdd vdd vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_26 dummy_bl dummy_br vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_26 vdd vdd vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_27 dummy_bl dummy_br vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_27 vdd vdd vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_28 dummy_bl dummy_br vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_28 vdd vdd vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_29 dummy_bl dummy_br vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_29 vdd vdd vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_30 dummy_bl dummy_br vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_30 vdd vdd vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_31 dummy_bl dummy_br vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_31 vdd vdd vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_32 dummy_bl dummy_br vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_32 vdd vdd vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_33 dummy_bl dummy_br vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_33 vdd vdd vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_34 dummy_bl dummy_br vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_34 vdd vdd vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_35 dummy_bl dummy_br vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_35 vdd vdd vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_36 dummy_bl dummy_br vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_36 vdd vdd vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_37 dummy_bl dummy_br vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_37 vdd vdd vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_38 dummy_bl dummy_br vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_38 vdd vdd vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_39 dummy_bl dummy_br vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_39 vdd vdd vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_40 dummy_bl dummy_br vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_40 vdd vdd vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_41 dummy_bl dummy_br vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_41 vdd vdd vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_42 dummy_bl dummy_br vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_42 vdd vdd vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_43 dummy_bl dummy_br vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_43 vdd vdd vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_44 dummy_bl dummy_br vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_44 vdd vdd vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_45 dummy_bl dummy_br vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_45 vdd vdd vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_46 dummy_bl dummy_br vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_46 vdd vdd vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_47 dummy_bl dummy_br vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_47 vdd vdd vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_48 dummy_bl dummy_br vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_48 vdd vdd vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_49 dummy_bl dummy_br vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_49 vdd vdd vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_50 dummy_bl dummy_br vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_50 vdd vdd vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_51 dummy_bl dummy_br vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_51 vdd vdd vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_52 dummy_bl dummy_br vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_52 vdd vdd vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_53 dummy_bl dummy_br vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_53 vdd vdd vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_54 dummy_bl dummy_br vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_54 vdd vdd vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_55 dummy_bl dummy_br vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_55 vdd vdd vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_56 dummy_bl dummy_br vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_56 vdd vdd vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_57 dummy_bl dummy_br vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_57 vdd vdd vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_58 dummy_bl dummy_br vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_58 vdd vdd vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_59 dummy_bl dummy_br vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_59 vdd vdd vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_60 dummy_bl dummy_br vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_60 vdd vdd vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_61 dummy_bl dummy_br vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_61 vdd vdd vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_62 dummy_bl dummy_br vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_62 vdd vdd vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_63 dummy_bl dummy_br vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_63 vdd vdd vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_64 dummy_bl dummy_br vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_64 vdd vdd vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_65 dummy_bl dummy_br vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_65 vdd vdd vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_66 dummy_bl dummy_br vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_66 vdd vdd vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_67 dummy_bl dummy_br vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_67 vdd vdd vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_68 dummy_bl dummy_br vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_68 vdd vdd vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_69 dummy_bl dummy_br vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_69 vdd vdd vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_70 dummy_bl dummy_br vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_70 vdd vdd vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_71 dummy_bl dummy_br vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_71 vdd vdd vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_72 dummy_bl dummy_br vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_72 vdd vdd vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_73 dummy_bl dummy_br vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_73 vdd vdd vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_74 dummy_bl dummy_br vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_74 vdd vdd vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_75 dummy_bl dummy_br vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_75 vdd vdd vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_76 dummy_bl dummy_br vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_76 vdd vdd vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_77 dummy_bl dummy_br vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_77 vdd vdd vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_78 dummy_bl dummy_br vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_78 vdd vdd vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_79 dummy_bl dummy_br vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_79 vdd vdd vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_80 dummy_bl dummy_br vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_80 vdd vdd vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_81 dummy_bl dummy_br vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_81 vdd vdd vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_82 dummy_bl dummy_br vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_82 vdd vdd vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_83 dummy_bl dummy_br vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_83 vdd vdd vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_84 dummy_bl dummy_br vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_84 vdd vdd vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_85 dummy_bl dummy_br vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_85 vdd vdd vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_86 dummy_bl dummy_br vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_86 vdd vdd vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_87 dummy_bl dummy_br vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_87 vdd vdd vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_88 dummy_bl dummy_br vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_88 vdd vdd vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_89 dummy_bl dummy_br vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_89 vdd vdd vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_90 dummy_bl dummy_br vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_90 vdd vdd vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_91 dummy_bl dummy_br vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_91 vdd vdd vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_92 dummy_bl dummy_br vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_92 vdd vdd vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_93 dummy_bl dummy_br vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_93 vdd vdd vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_94 dummy_bl dummy_br vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_94 vdd vdd vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_95 dummy_bl dummy_br vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_95 vdd vdd vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_96 dummy_bl dummy_br vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_96 vdd vdd vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_97 dummy_bl dummy_br vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_97 vdd vdd vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_98 dummy_bl dummy_br vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_98 vdd vdd vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_99 dummy_bl dummy_br vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_99 vdd vdd vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_100 dummy_bl dummy_br vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_100 vdd vdd vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_101 dummy_bl dummy_br vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_101 vdd vdd vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_102 dummy_bl dummy_br vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_102 vdd vdd vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_103 dummy_bl dummy_br vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_103 vdd vdd vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_104 dummy_bl dummy_br vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_104 vdd vdd vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_105 dummy_bl dummy_br vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_105 vdd vdd vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_106 dummy_bl dummy_br vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_106 vdd vdd vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_107 dummy_bl dummy_br vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_107 vdd vdd vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_108 dummy_bl dummy_br vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_108 vdd vdd vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_109 dummy_bl dummy_br vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_109 vdd vdd vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_110 dummy_bl dummy_br vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_110 vdd vdd vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_111 dummy_bl dummy_br vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_111 vdd vdd vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_112 dummy_bl dummy_br vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_112 vdd vdd vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_113 dummy_bl dummy_br vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_113 vdd vdd vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_114 dummy_bl dummy_br vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_114 vdd vdd vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_115 dummy_bl dummy_br vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_115 vdd vdd vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_116 dummy_bl dummy_br vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_116 vdd vdd vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_117 dummy_bl dummy_br vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_117 vdd vdd vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_118 dummy_bl dummy_br vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_118 vdd vdd vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_119 dummy_bl dummy_br vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_119 vdd vdd vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_120 dummy_bl dummy_br vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_120 vdd vdd vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_121 dummy_bl dummy_br vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_121 vdd vdd vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_122 dummy_bl dummy_br vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_122 vdd vdd vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_123 dummy_bl dummy_br vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_123 vdd vdd vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_124 dummy_bl dummy_br vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_124 vdd vdd vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_125 dummy_bl dummy_br vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_125 vdd vdd vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_126 dummy_bl dummy_br vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_126 vdd vdd vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_127 dummy_bl dummy_br vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_127 vdd vdd vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_128 dummy_bl dummy_br vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_128 vdd vdd vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_129 dummy_bl dummy_br vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_129 vdd vdd vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_0 bl[0] br[0] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_0 bl[0] br[0] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_1 bl[1] br[1] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_1 bl[1] br[1] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_2 bl[2] br[2] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_2 bl[2] br[2] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_3 bl[3] br[3] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_3 bl[3] br[3] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_4 bl[4] br[4] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_4 bl[4] br[4] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_5 bl[5] br[5] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_5 bl[5] br[5] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_6 bl[6] br[6] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_6 bl[6] br[6] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_7 bl[7] br[7] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_7 bl[7] br[7] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_8 bl[8] br[8] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_8 bl[8] br[8] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_9 bl[9] br[9] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_9 bl[9] br[9] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_10 bl[10] br[10] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_10 bl[10] br[10] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_11 bl[11] br[11] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_11 bl[11] br[11] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_12 bl[12] br[12] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_12 bl[12] br[12] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_13 bl[13] br[13] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_13 bl[13] br[13] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_14 bl[14] br[14] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_14 bl[14] br[14] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_15 bl[15] br[15] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_15 bl[15] br[15] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_16 bl[16] br[16] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_16 bl[16] br[16] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_17 bl[17] br[17] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_17 bl[17] br[17] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_18 bl[18] br[18] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_18 bl[18] br[18] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_19 bl[19] br[19] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_19 bl[19] br[19] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_20 bl[20] br[20] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_20 bl[20] br[20] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_21 bl[21] br[21] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_21 bl[21] br[21] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_22 bl[22] br[22] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_22 bl[22] br[22] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_23 bl[23] br[23] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_23 bl[23] br[23] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_24 bl[24] br[24] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_24 bl[24] br[24] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_25 bl[25] br[25] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_25 bl[25] br[25] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_26 bl[26] br[26] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_26 bl[26] br[26] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_27 bl[27] br[27] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_27 bl[27] br[27] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_28 bl[28] br[28] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_28 bl[28] br[28] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_29 bl[29] br[29] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_29 bl[29] br[29] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_30 bl[30] br[30] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_30 bl[30] br[30] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_31 bl[31] br[31] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_31 bl[31] br[31] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_32 bl[32] br[32] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_32 bl[32] br[32] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_33 bl[33] br[33] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_33 bl[33] br[33] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_34 bl[34] br[34] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_34 bl[34] br[34] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_35 bl[35] br[35] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_35 bl[35] br[35] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_36 bl[36] br[36] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_36 bl[36] br[36] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_37 bl[37] br[37] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_37 bl[37] br[37] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_38 bl[38] br[38] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_38 bl[38] br[38] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_39 bl[39] br[39] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_39 bl[39] br[39] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_40 bl[40] br[40] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_40 bl[40] br[40] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_41 bl[41] br[41] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_41 bl[41] br[41] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_42 bl[42] br[42] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_42 bl[42] br[42] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_43 bl[43] br[43] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_43 bl[43] br[43] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_44 bl[44] br[44] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_44 bl[44] br[44] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_45 bl[45] br[45] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_45 bl[45] br[45] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_46 bl[46] br[46] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_46 bl[46] br[46] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_47 bl[47] br[47] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_47 bl[47] br[47] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_48 bl[48] br[48] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_48 bl[48] br[48] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_49 bl[49] br[49] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_49 bl[49] br[49] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_50 bl[50] br[50] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_50 bl[50] br[50] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_51 bl[51] br[51] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_51 bl[51] br[51] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_52 bl[52] br[52] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_52 bl[52] br[52] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_53 bl[53] br[53] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_53 bl[53] br[53] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_54 bl[54] br[54] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_54 bl[54] br[54] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_55 bl[55] br[55] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_55 bl[55] br[55] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_56 bl[56] br[56] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_56 bl[56] br[56] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_57 bl[57] br[57] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_57 bl[57] br[57] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_58 bl[58] br[58] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_58 bl[58] br[58] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_59 bl[59] br[59] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_59 bl[59] br[59] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_60 bl[60] br[60] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_60 bl[60] br[60] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_61 bl[61] br[61] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_61 bl[61] br[61] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_62 bl[62] br[62] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_62 bl[62] br[62] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_63 bl[63] br[63] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_63 bl[63] br[63] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_64 bl[64] br[64] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_64 bl[64] br[64] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_65 bl[65] br[65] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_65 bl[65] br[65] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_66 bl[66] br[66] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_66 bl[66] br[66] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_67 bl[67] br[67] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_67 bl[67] br[67] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_68 bl[68] br[68] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_68 bl[68] br[68] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_69 bl[69] br[69] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_69 bl[69] br[69] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_70 bl[70] br[70] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_70 bl[70] br[70] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_71 bl[71] br[71] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_71 bl[71] br[71] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_72 bl[72] br[72] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_72 bl[72] br[72] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_73 bl[73] br[73] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_73 bl[73] br[73] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_74 bl[74] br[74] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_74 bl[74] br[74] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_75 bl[75] br[75] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_75 bl[75] br[75] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_76 bl[76] br[76] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_76 bl[76] br[76] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_77 bl[77] br[77] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_77 bl[77] br[77] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_78 bl[78] br[78] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_78 bl[78] br[78] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_79 bl[79] br[79] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_79 bl[79] br[79] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_80 bl[80] br[80] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_80 bl[80] br[80] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_81 bl[81] br[81] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_81 bl[81] br[81] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_82 bl[82] br[82] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_82 bl[82] br[82] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_83 bl[83] br[83] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_83 bl[83] br[83] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_84 bl[84] br[84] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_84 bl[84] br[84] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_85 bl[85] br[85] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_85 bl[85] br[85] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_86 bl[86] br[86] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_86 bl[86] br[86] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_87 bl[87] br[87] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_87 bl[87] br[87] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_88 bl[88] br[88] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_88 bl[88] br[88] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_89 bl[89] br[89] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_89 bl[89] br[89] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_90 bl[90] br[90] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_90 bl[90] br[90] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_91 bl[91] br[91] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_91 bl[91] br[91] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_92 bl[92] br[92] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_92 bl[92] br[92] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_93 bl[93] br[93] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_93 bl[93] br[93] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_94 bl[94] br[94] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_94 bl[94] br[94] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_95 bl[95] br[95] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_95 bl[95] br[95] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_96 bl[96] br[96] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_96 bl[96] br[96] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_97 bl[97] br[97] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_97 bl[97] br[97] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_98 bl[98] br[98] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_98 bl[98] br[98] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_99 bl[99] br[99] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_99 bl[99] br[99] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_100 bl[100] br[100] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_100 bl[100] br[100] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_101 bl[101] br[101] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_101 bl[101] br[101] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_102 bl[102] br[102] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_102 bl[102] br[102] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_103 bl[103] br[103] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_103 bl[103] br[103] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_104 bl[104] br[104] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_104 bl[104] br[104] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_105 bl[105] br[105] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_105 bl[105] br[105] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_106 bl[106] br[106] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_106 bl[106] br[106] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_107 bl[107] br[107] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_107 bl[107] br[107] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_108 bl[108] br[108] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_108 bl[108] br[108] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_109 bl[109] br[109] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_109 bl[109] br[109] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_110 bl[110] br[110] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_110 bl[110] br[110] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_111 bl[111] br[111] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_111 bl[111] br[111] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_112 bl[112] br[112] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_112 bl[112] br[112] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_113 bl[113] br[113] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_113 bl[113] br[113] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_114 bl[114] br[114] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_114 bl[114] br[114] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_115 bl[115] br[115] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_115 bl[115] br[115] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_116 bl[116] br[116] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_116 bl[116] br[116] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_117 bl[117] br[117] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_117 bl[117] br[117] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_118 bl[118] br[118] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_118 bl[118] br[118] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_119 bl[119] br[119] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_119 bl[119] br[119] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_120 bl[120] br[120] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_120 bl[120] br[120] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_121 bl[121] br[121] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_121 bl[121] br[121] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_122 bl[122] br[122] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_122 bl[122] br[122] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_123 bl[123] br[123] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_123 bl[123] br[123] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_124 bl[124] br[124] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_124 bl[124] br[124] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_125 bl[125] br[125] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_125 bl[125] br[125] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_126 bl[126] br[126] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_126 bl[126] br[126] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_127 bl[127] br[127] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_127 bl[127] br[127] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_128 bl[128] br[128] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_128 bl[128] br[128] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_129 bl[129] br[129] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_129 bl[129] br[129] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_130 bl[130] br[130] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_130 bl[130] br[130] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_131 bl[131] br[131] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_131 bl[131] br[131] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_132 bl[132] br[132] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_132 bl[132] br[132] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_133 bl[133] br[133] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_133 bl[133] br[133] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_134 bl[134] br[134] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_134 bl[134] br[134] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_135 bl[135] br[135] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_135 bl[135] br[135] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_136 bl[136] br[136] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_136 bl[136] br[136] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_137 bl[137] br[137] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_137 bl[137] br[137] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_138 bl[138] br[138] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_138 bl[138] br[138] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_139 bl[139] br[139] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_139 bl[139] br[139] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_140 bl[140] br[140] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_140 bl[140] br[140] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_141 bl[141] br[141] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_141 bl[141] br[141] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_142 bl[142] br[142] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_142 bl[142] br[142] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_143 bl[143] br[143] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_143 bl[143] br[143] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_144 bl[144] br[144] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_144 bl[144] br[144] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_145 bl[145] br[145] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_145 bl[145] br[145] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_146 bl[146] br[146] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_146 bl[146] br[146] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_147 bl[147] br[147] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_147 bl[147] br[147] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_148 bl[148] br[148] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_148 bl[148] br[148] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_149 bl[149] br[149] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_149 bl[149] br[149] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_150 bl[150] br[150] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_150 bl[150] br[150] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_151 bl[151] br[151] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_151 bl[151] br[151] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_152 bl[152] br[152] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_152 bl[152] br[152] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_153 bl[153] br[153] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_153 bl[153] br[153] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_154 bl[154] br[154] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_154 bl[154] br[154] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_155 bl[155] br[155] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_155 bl[155] br[155] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_156 bl[156] br[156] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_156 bl[156] br[156] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_157 bl[157] br[157] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_157 bl[157] br[157] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_158 bl[158] br[158] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_158 bl[158] br[158] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_159 bl[159] br[159] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_159 bl[159] br[159] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_160 bl[160] br[160] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_160 bl[160] br[160] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_161 bl[161] br[161] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_161 bl[161] br[161] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_162 bl[162] br[162] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_162 bl[162] br[162] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_163 bl[163] br[163] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_163 bl[163] br[163] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_164 bl[164] br[164] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_164 bl[164] br[164] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_165 bl[165] br[165] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_165 bl[165] br[165] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_166 bl[166] br[166] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_166 bl[166] br[166] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_167 bl[167] br[167] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_167 bl[167] br[167] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_168 bl[168] br[168] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_168 bl[168] br[168] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_169 bl[169] br[169] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_169 bl[169] br[169] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_170 bl[170] br[170] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_170 bl[170] br[170] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_171 bl[171] br[171] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_171 bl[171] br[171] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_172 bl[172] br[172] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_172 bl[172] br[172] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_173 bl[173] br[173] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_173 bl[173] br[173] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_174 bl[174] br[174] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_174 bl[174] br[174] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_175 bl[175] br[175] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_175 bl[175] br[175] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_176 bl[176] br[176] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_176 bl[176] br[176] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_177 bl[177] br[177] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_177 bl[177] br[177] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_178 bl[178] br[178] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_178 bl[178] br[178] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_179 bl[179] br[179] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_179 bl[179] br[179] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_180 bl[180] br[180] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_180 bl[180] br[180] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_181 bl[181] br[181] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_181 bl[181] br[181] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_182 bl[182] br[182] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_182 bl[182] br[182] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_183 bl[183] br[183] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_183 bl[183] br[183] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_184 bl[184] br[184] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_184 bl[184] br[184] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_185 bl[185] br[185] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_185 bl[185] br[185] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_186 bl[186] br[186] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_186 bl[186] br[186] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_187 bl[187] br[187] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_187 bl[187] br[187] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_188 bl[188] br[188] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_188 bl[188] br[188] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_189 bl[189] br[189] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_189 bl[189] br[189] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_190 bl[190] br[190] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_190 bl[190] br[190] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_191 bl[191] br[191] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_191 bl[191] br[191] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_192 bl[192] br[192] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_192 bl[192] br[192] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_193 bl[193] br[193] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_193 bl[193] br[193] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_194 bl[194] br[194] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_194 bl[194] br[194] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_195 bl[195] br[195] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_195 bl[195] br[195] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_196 bl[196] br[196] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_196 bl[196] br[196] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_197 bl[197] br[197] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_197 bl[197] br[197] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_198 bl[198] br[198] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_198 bl[198] br[198] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_199 bl[199] br[199] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_199 bl[199] br[199] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_200 bl[200] br[200] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_200 bl[200] br[200] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_201 bl[201] br[201] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_201 bl[201] br[201] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_202 bl[202] br[202] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_202 bl[202] br[202] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_203 bl[203] br[203] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_203 bl[203] br[203] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_204 bl[204] br[204] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_204 bl[204] br[204] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_205 bl[205] br[205] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_205 bl[205] br[205] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_206 bl[206] br[206] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_206 bl[206] br[206] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_207 bl[207] br[207] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_207 bl[207] br[207] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_208 bl[208] br[208] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_208 bl[208] br[208] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_209 bl[209] br[209] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_209 bl[209] br[209] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_210 bl[210] br[210] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_210 bl[210] br[210] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_211 bl[211] br[211] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_211 bl[211] br[211] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_212 bl[212] br[212] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_212 bl[212] br[212] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_213 bl[213] br[213] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_213 bl[213] br[213] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_214 bl[214] br[214] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_214 bl[214] br[214] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_215 bl[215] br[215] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_215 bl[215] br[215] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_216 bl[216] br[216] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_216 bl[216] br[216] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_217 bl[217] br[217] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_217 bl[217] br[217] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_218 bl[218] br[218] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_218 bl[218] br[218] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_219 bl[219] br[219] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_219 bl[219] br[219] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_220 bl[220] br[220] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_220 bl[220] br[220] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_221 bl[221] br[221] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_221 bl[221] br[221] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_222 bl[222] br[222] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_222 bl[222] br[222] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_223 bl[223] br[223] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_223 bl[223] br[223] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_224 bl[224] br[224] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_224 bl[224] br[224] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_225 bl[225] br[225] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_225 bl[225] br[225] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_226 bl[226] br[226] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_226 bl[226] br[226] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_227 bl[227] br[227] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_227 bl[227] br[227] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_228 bl[228] br[228] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_228 bl[228] br[228] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_229 bl[229] br[229] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_229 bl[229] br[229] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_230 bl[230] br[230] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_230 bl[230] br[230] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_231 bl[231] br[231] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_231 bl[231] br[231] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_232 bl[232] br[232] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_232 bl[232] br[232] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_233 bl[233] br[233] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_233 bl[233] br[233] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_234 bl[234] br[234] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_234 bl[234] br[234] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_235 bl[235] br[235] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_235 bl[235] br[235] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_236 bl[236] br[236] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_236 bl[236] br[236] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_237 bl[237] br[237] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_237 bl[237] br[237] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_238 bl[238] br[238] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_238 bl[238] br[238] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_239 bl[239] br[239] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_239 bl[239] br[239] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_240 bl[240] br[240] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_240 bl[240] br[240] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_241 bl[241] br[241] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_241 bl[241] br[241] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_242 bl[242] br[242] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_242 bl[242] br[242] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_243 bl[243] br[243] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_243 bl[243] br[243] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_244 bl[244] br[244] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_244 bl[244] br[244] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_245 bl[245] br[245] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_245 bl[245] br[245] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_246 bl[246] br[246] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_246 bl[246] br[246] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_247 bl[247] br[247] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_247 bl[247] br[247] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_248 bl[248] br[248] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_248 bl[248] br[248] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_249 bl[249] br[249] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_249 bl[249] br[249] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_250 bl[250] br[250] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_250 bl[250] br[250] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_251 bl[251] br[251] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_251 bl[251] br[251] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_252 bl[252] br[252] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_252 bl[252] br[252] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_253 bl[253] br[253] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_253 bl[253] br[253] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_254 bl[254] br[254] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_254 bl[254] br[254] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_255 bl[255] br[255] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_255 bl[255] br[255] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xcolend_top_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_colend_wrapper
  Xcolend_bot_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_colend_wrapper
  Xhstrap_0_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_1 br[0] vdd vss bl[0] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_1 br[0] vdd vss bl[0] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_2 br[1] vdd vss bl[1] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_2 br[1] vdd vss bl[1] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_3 br[2] vdd vss bl[2] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_3 br[2] vdd vss bl[2] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_4 br[3] vdd vss bl[3] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_4 br[3] vdd vss bl[3] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_5 br[4] vdd vss bl[4] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_5 br[4] vdd vss bl[4] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_6 br[5] vdd vss bl[5] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_6 br[5] vdd vss bl[5] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_7 br[6] vdd vss bl[6] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_7 br[6] vdd vss bl[6] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_8 br[7] vdd vss bl[7] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_8 br[7] vdd vss bl[7] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_9 br[8] vdd vss bl[8] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_9 br[8] vdd vss bl[8] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_10 br[9] vdd vss bl[9] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_10 br[9] vdd vss bl[9] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_11 br[10] vdd vss bl[10] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_11 br[10] vdd vss bl[10] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_12 br[11] vdd vss bl[11] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_12 br[11] vdd vss bl[11] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_13 br[12] vdd vss bl[12] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_13 br[12] vdd vss bl[12] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_14 br[13] vdd vss bl[13] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_14 br[13] vdd vss bl[13] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_15 br[14] vdd vss bl[14] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_15 br[14] vdd vss bl[14] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_16 br[15] vdd vss bl[15] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_16 br[15] vdd vss bl[15] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_17 br[16] vdd vss bl[16] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_17 br[16] vdd vss bl[16] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_18 br[17] vdd vss bl[17] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_18 br[17] vdd vss bl[17] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_19 br[18] vdd vss bl[18] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_19 br[18] vdd vss bl[18] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_20 br[19] vdd vss bl[19] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_20 br[19] vdd vss bl[19] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_21 br[20] vdd vss bl[20] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_21 br[20] vdd vss bl[20] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_22 br[21] vdd vss bl[21] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_22 br[21] vdd vss bl[21] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_23 br[22] vdd vss bl[22] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_23 br[22] vdd vss bl[22] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_24 br[23] vdd vss bl[23] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_24 br[23] vdd vss bl[23] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_25 br[24] vdd vss bl[24] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_25 br[24] vdd vss bl[24] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_26 br[25] vdd vss bl[25] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_26 br[25] vdd vss bl[25] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_27 br[26] vdd vss bl[26] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_27 br[26] vdd vss bl[26] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_28 br[27] vdd vss bl[27] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_28 br[27] vdd vss bl[27] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_29 br[28] vdd vss bl[28] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_29 br[28] vdd vss bl[28] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_30 br[29] vdd vss bl[29] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_30 br[29] vdd vss bl[29] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_31 br[30] vdd vss bl[30] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_31 br[30] vdd vss bl[30] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_32 br[31] vdd vss bl[31] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_32 br[31] vdd vss bl[31] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_33 br[32] vdd vss bl[32] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_33 br[32] vdd vss bl[32] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_34 br[33] vdd vss bl[33] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_34 br[33] vdd vss bl[33] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_35 br[34] vdd vss bl[34] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_35 br[34] vdd vss bl[34] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_36 br[35] vdd vss bl[35] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_36 br[35] vdd vss bl[35] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_37 br[36] vdd vss bl[36] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_37 br[36] vdd vss bl[36] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_38 br[37] vdd vss bl[37] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_38 br[37] vdd vss bl[37] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_39 br[38] vdd vss bl[38] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_39 br[38] vdd vss bl[38] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_40 br[39] vdd vss bl[39] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_40 br[39] vdd vss bl[39] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_41 br[40] vdd vss bl[40] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_41 br[40] vdd vss bl[40] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_42 br[41] vdd vss bl[41] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_42 br[41] vdd vss bl[41] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_43 br[42] vdd vss bl[42] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_43 br[42] vdd vss bl[42] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_44 br[43] vdd vss bl[43] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_44 br[43] vdd vss bl[43] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_45 br[44] vdd vss bl[44] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_45 br[44] vdd vss bl[44] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_46 br[45] vdd vss bl[45] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_46 br[45] vdd vss bl[45] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_47 br[46] vdd vss bl[46] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_47 br[46] vdd vss bl[46] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_48 br[47] vdd vss bl[47] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_48 br[47] vdd vss bl[47] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_49 br[48] vdd vss bl[48] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_49 br[48] vdd vss bl[48] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_50 br[49] vdd vss bl[49] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_50 br[49] vdd vss bl[49] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_51 br[50] vdd vss bl[50] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_51 br[50] vdd vss bl[50] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_52 br[51] vdd vss bl[51] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_52 br[51] vdd vss bl[51] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_53 br[52] vdd vss bl[52] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_53 br[52] vdd vss bl[52] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_54 br[53] vdd vss bl[53] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_54 br[53] vdd vss bl[53] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_55 br[54] vdd vss bl[54] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_55 br[54] vdd vss bl[54] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_56 br[55] vdd vss bl[55] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_56 br[55] vdd vss bl[55] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_57 br[56] vdd vss bl[56] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_57 br[56] vdd vss bl[56] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_58 br[57] vdd vss bl[57] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_58 br[57] vdd vss bl[57] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_59 br[58] vdd vss bl[58] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_59 br[58] vdd vss bl[58] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_60 br[59] vdd vss bl[59] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_60 br[59] vdd vss bl[59] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_61 br[60] vdd vss bl[60] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_61 br[60] vdd vss bl[60] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_62 br[61] vdd vss bl[61] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_62 br[61] vdd vss bl[61] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_63 br[62] vdd vss bl[62] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_63 br[62] vdd vss bl[62] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_64 br[63] vdd vss bl[63] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_64 br[63] vdd vss bl[63] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_65 br[64] vdd vss bl[64] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_65 br[64] vdd vss bl[64] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_66 br[65] vdd vss bl[65] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_66 br[65] vdd vss bl[65] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_67 br[66] vdd vss bl[66] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_67 br[66] vdd vss bl[66] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_68 br[67] vdd vss bl[67] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_68 br[67] vdd vss bl[67] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_69 br[68] vdd vss bl[68] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_69 br[68] vdd vss bl[68] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_70 br[69] vdd vss bl[69] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_70 br[69] vdd vss bl[69] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_71 br[70] vdd vss bl[70] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_71 br[70] vdd vss bl[70] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_72 br[71] vdd vss bl[71] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_72 br[71] vdd vss bl[71] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_73 br[72] vdd vss bl[72] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_73 br[72] vdd vss bl[72] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_74 br[73] vdd vss bl[73] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_74 br[73] vdd vss bl[73] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_75 br[74] vdd vss bl[74] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_75 br[74] vdd vss bl[74] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_76 br[75] vdd vss bl[75] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_76 br[75] vdd vss bl[75] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_77 br[76] vdd vss bl[76] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_77 br[76] vdd vss bl[76] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_78 br[77] vdd vss bl[77] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_78 br[77] vdd vss bl[77] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_79 br[78] vdd vss bl[78] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_79 br[78] vdd vss bl[78] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_80 br[79] vdd vss bl[79] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_80 br[79] vdd vss bl[79] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_81 br[80] vdd vss bl[80] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_81 br[80] vdd vss bl[80] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_82 br[81] vdd vss bl[81] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_82 br[81] vdd vss bl[81] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_83 br[82] vdd vss bl[82] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_83 br[82] vdd vss bl[82] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_84 br[83] vdd vss bl[83] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_84 br[83] vdd vss bl[83] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_85 br[84] vdd vss bl[84] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_85 br[84] vdd vss bl[84] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_86 br[85] vdd vss bl[85] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_86 br[85] vdd vss bl[85] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_87 br[86] vdd vss bl[86] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_87 br[86] vdd vss bl[86] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_88 br[87] vdd vss bl[87] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_88 br[87] vdd vss bl[87] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_89 br[88] vdd vss bl[88] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_89 br[88] vdd vss bl[88] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_90 br[89] vdd vss bl[89] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_90 br[89] vdd vss bl[89] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_91 br[90] vdd vss bl[90] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_91 br[90] vdd vss bl[90] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_92 br[91] vdd vss bl[91] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_92 br[91] vdd vss bl[91] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_93 br[92] vdd vss bl[92] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_93 br[92] vdd vss bl[92] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_94 br[93] vdd vss bl[93] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_94 br[93] vdd vss bl[93] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_95 br[94] vdd vss bl[94] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_95 br[94] vdd vss bl[94] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_96 br[95] vdd vss bl[95] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_96 br[95] vdd vss bl[95] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_97 br[96] vdd vss bl[96] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_97 br[96] vdd vss bl[96] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_98 br[97] vdd vss bl[97] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_98 br[97] vdd vss bl[97] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_99 br[98] vdd vss bl[98] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_99 br[98] vdd vss bl[98] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_100 br[99] vdd vss bl[99] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_100 br[99] vdd vss bl[99] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_101 br[100] vdd vss bl[100] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_101 br[100] vdd vss bl[100] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_102 br[101] vdd vss bl[101] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_102 br[101] vdd vss bl[101] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_103 br[102] vdd vss bl[102] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_103 br[102] vdd vss bl[102] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_104 br[103] vdd vss bl[103] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_104 br[103] vdd vss bl[103] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_105 br[104] vdd vss bl[104] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_105 br[104] vdd vss bl[104] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_106 br[105] vdd vss bl[105] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_106 br[105] vdd vss bl[105] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_107 br[106] vdd vss bl[106] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_107 br[106] vdd vss bl[106] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_108 br[107] vdd vss bl[107] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_108 br[107] vdd vss bl[107] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_109 br[108] vdd vss bl[108] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_109 br[108] vdd vss bl[108] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_110 br[109] vdd vss bl[109] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_110 br[109] vdd vss bl[109] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_111 br[110] vdd vss bl[110] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_111 br[110] vdd vss bl[110] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_112 br[111] vdd vss bl[111] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_112 br[111] vdd vss bl[111] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_113 br[112] vdd vss bl[112] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_113 br[112] vdd vss bl[112] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_114 br[113] vdd vss bl[113] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_114 br[113] vdd vss bl[113] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_115 br[114] vdd vss bl[114] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_115 br[114] vdd vss bl[114] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_116 br[115] vdd vss bl[115] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_116 br[115] vdd vss bl[115] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_117 br[116] vdd vss bl[116] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_117 br[116] vdd vss bl[116] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_118 br[117] vdd vss bl[117] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_118 br[117] vdd vss bl[117] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_119 br[118] vdd vss bl[118] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_119 br[118] vdd vss bl[118] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_120 br[119] vdd vss bl[119] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_120 br[119] vdd vss bl[119] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_121 br[120] vdd vss bl[120] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_121 br[120] vdd vss bl[120] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_122 br[121] vdd vss bl[121] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_122 br[121] vdd vss bl[121] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_123 br[122] vdd vss bl[122] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_123 br[122] vdd vss bl[122] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_124 br[123] vdd vss bl[123] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_124 br[123] vdd vss bl[123] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_125 br[124] vdd vss bl[124] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_125 br[124] vdd vss bl[124] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_126 br[125] vdd vss bl[125] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_126 br[125] vdd vss bl[125] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_127 br[126] vdd vss bl[126] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_127 br[126] vdd vss bl[126] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_128 br[127] vdd vss bl[127] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_128 br[127] vdd vss bl[127] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_129 br[128] vdd vss bl[128] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_129 br[128] vdd vss bl[128] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_130 br[129] vdd vss bl[129] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_130 br[129] vdd vss bl[129] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_131 br[130] vdd vss bl[130] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_131 br[130] vdd vss bl[130] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_132 br[131] vdd vss bl[131] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_132 br[131] vdd vss bl[131] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_133 br[132] vdd vss bl[132] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_133 br[132] vdd vss bl[132] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_134 br[133] vdd vss bl[133] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_134 br[133] vdd vss bl[133] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_135 br[134] vdd vss bl[134] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_135 br[134] vdd vss bl[134] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_136 br[135] vdd vss bl[135] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_136 br[135] vdd vss bl[135] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_137 br[136] vdd vss bl[136] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_137 br[136] vdd vss bl[136] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_138 br[137] vdd vss bl[137] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_138 br[137] vdd vss bl[137] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_139 br[138] vdd vss bl[138] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_139 br[138] vdd vss bl[138] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_140 br[139] vdd vss bl[139] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_140 br[139] vdd vss bl[139] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_141 br[140] vdd vss bl[140] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_141 br[140] vdd vss bl[140] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_142 br[141] vdd vss bl[141] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_142 br[141] vdd vss bl[141] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_143 br[142] vdd vss bl[142] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_143 br[142] vdd vss bl[142] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_144 br[143] vdd vss bl[143] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_144 br[143] vdd vss bl[143] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_145 br[144] vdd vss bl[144] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_145 br[144] vdd vss bl[144] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_146 br[145] vdd vss bl[145] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_146 br[145] vdd vss bl[145] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_147 br[146] vdd vss bl[146] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_147 br[146] vdd vss bl[146] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_148 br[147] vdd vss bl[147] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_148 br[147] vdd vss bl[147] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_149 br[148] vdd vss bl[148] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_149 br[148] vdd vss bl[148] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_150 br[149] vdd vss bl[149] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_150 br[149] vdd vss bl[149] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_151 br[150] vdd vss bl[150] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_151 br[150] vdd vss bl[150] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_152 br[151] vdd vss bl[151] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_152 br[151] vdd vss bl[151] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_153 br[152] vdd vss bl[152] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_153 br[152] vdd vss bl[152] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_154 br[153] vdd vss bl[153] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_154 br[153] vdd vss bl[153] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_155 br[154] vdd vss bl[154] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_155 br[154] vdd vss bl[154] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_156 br[155] vdd vss bl[155] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_156 br[155] vdd vss bl[155] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_157 br[156] vdd vss bl[156] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_157 br[156] vdd vss bl[156] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_158 br[157] vdd vss bl[157] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_158 br[157] vdd vss bl[157] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_159 br[158] vdd vss bl[158] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_159 br[158] vdd vss bl[158] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_160 br[159] vdd vss bl[159] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_160 br[159] vdd vss bl[159] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_161 br[160] vdd vss bl[160] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_161 br[160] vdd vss bl[160] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_162 br[161] vdd vss bl[161] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_162 br[161] vdd vss bl[161] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_163 br[162] vdd vss bl[162] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_163 br[162] vdd vss bl[162] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_164 br[163] vdd vss bl[163] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_164 br[163] vdd vss bl[163] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_165 br[164] vdd vss bl[164] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_165 br[164] vdd vss bl[164] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_166 br[165] vdd vss bl[165] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_166 br[165] vdd vss bl[165] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_167 br[166] vdd vss bl[166] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_167 br[166] vdd vss bl[166] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_168 br[167] vdd vss bl[167] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_168 br[167] vdd vss bl[167] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_169 br[168] vdd vss bl[168] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_169 br[168] vdd vss bl[168] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_170 br[169] vdd vss bl[169] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_170 br[169] vdd vss bl[169] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_171 br[170] vdd vss bl[170] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_171 br[170] vdd vss bl[170] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_172 br[171] vdd vss bl[171] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_172 br[171] vdd vss bl[171] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_173 br[172] vdd vss bl[172] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_173 br[172] vdd vss bl[172] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_174 br[173] vdd vss bl[173] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_174 br[173] vdd vss bl[173] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_175 br[174] vdd vss bl[174] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_175 br[174] vdd vss bl[174] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_176 br[175] vdd vss bl[175] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_176 br[175] vdd vss bl[175] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_177 br[176] vdd vss bl[176] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_177 br[176] vdd vss bl[176] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_178 br[177] vdd vss bl[177] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_178 br[177] vdd vss bl[177] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_179 br[178] vdd vss bl[178] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_179 br[178] vdd vss bl[178] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_180 br[179] vdd vss bl[179] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_180 br[179] vdd vss bl[179] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_181 br[180] vdd vss bl[180] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_181 br[180] vdd vss bl[180] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_182 br[181] vdd vss bl[181] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_182 br[181] vdd vss bl[181] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_183 br[182] vdd vss bl[182] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_183 br[182] vdd vss bl[182] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_184 br[183] vdd vss bl[183] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_184 br[183] vdd vss bl[183] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_185 br[184] vdd vss bl[184] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_185 br[184] vdd vss bl[184] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_186 br[185] vdd vss bl[185] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_186 br[185] vdd vss bl[185] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_187 br[186] vdd vss bl[186] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_187 br[186] vdd vss bl[186] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_188 br[187] vdd vss bl[187] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_188 br[187] vdd vss bl[187] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_189 br[188] vdd vss bl[188] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_189 br[188] vdd vss bl[188] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_190 br[189] vdd vss bl[189] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_190 br[189] vdd vss bl[189] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_191 br[190] vdd vss bl[190] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_191 br[190] vdd vss bl[190] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_192 br[191] vdd vss bl[191] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_192 br[191] vdd vss bl[191] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_193 br[192] vdd vss bl[192] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_193 br[192] vdd vss bl[192] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_194 br[193] vdd vss bl[193] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_194 br[193] vdd vss bl[193] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_195 br[194] vdd vss bl[194] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_195 br[194] vdd vss bl[194] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_196 br[195] vdd vss bl[195] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_196 br[195] vdd vss bl[195] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_197 br[196] vdd vss bl[196] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_197 br[196] vdd vss bl[196] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_198 br[197] vdd vss bl[197] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_198 br[197] vdd vss bl[197] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_199 br[198] vdd vss bl[198] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_199 br[198] vdd vss bl[198] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_200 br[199] vdd vss bl[199] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_200 br[199] vdd vss bl[199] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_201 br[200] vdd vss bl[200] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_201 br[200] vdd vss bl[200] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_202 br[201] vdd vss bl[201] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_202 br[201] vdd vss bl[201] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_203 br[202] vdd vss bl[202] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_203 br[202] vdd vss bl[202] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_204 br[203] vdd vss bl[203] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_204 br[203] vdd vss bl[203] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_205 br[204] vdd vss bl[204] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_205 br[204] vdd vss bl[204] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_206 br[205] vdd vss bl[205] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_206 br[205] vdd vss bl[205] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_207 br[206] vdd vss bl[206] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_207 br[206] vdd vss bl[206] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_208 br[207] vdd vss bl[207] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_208 br[207] vdd vss bl[207] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_209 br[208] vdd vss bl[208] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_209 br[208] vdd vss bl[208] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_210 br[209] vdd vss bl[209] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_210 br[209] vdd vss bl[209] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_211 br[210] vdd vss bl[210] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_211 br[210] vdd vss bl[210] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_212 br[211] vdd vss bl[211] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_212 br[211] vdd vss bl[211] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_213 br[212] vdd vss bl[212] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_213 br[212] vdd vss bl[212] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_214 br[213] vdd vss bl[213] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_214 br[213] vdd vss bl[213] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_215 br[214] vdd vss bl[214] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_215 br[214] vdd vss bl[214] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_216 br[215] vdd vss bl[215] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_216 br[215] vdd vss bl[215] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_217 br[216] vdd vss bl[216] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_217 br[216] vdd vss bl[216] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_218 br[217] vdd vss bl[217] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_218 br[217] vdd vss bl[217] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_219 br[218] vdd vss bl[218] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_219 br[218] vdd vss bl[218] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_220 br[219] vdd vss bl[219] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_220 br[219] vdd vss bl[219] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_221 br[220] vdd vss bl[220] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_221 br[220] vdd vss bl[220] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_222 br[221] vdd vss bl[221] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_222 br[221] vdd vss bl[221] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_223 br[222] vdd vss bl[222] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_223 br[222] vdd vss bl[222] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_224 br[223] vdd vss bl[223] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_224 br[223] vdd vss bl[223] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_225 br[224] vdd vss bl[224] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_225 br[224] vdd vss bl[224] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_226 br[225] vdd vss bl[225] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_226 br[225] vdd vss bl[225] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_227 br[226] vdd vss bl[226] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_227 br[226] vdd vss bl[226] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_228 br[227] vdd vss bl[227] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_228 br[227] vdd vss bl[227] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_229 br[228] vdd vss bl[228] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_229 br[228] vdd vss bl[228] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_230 br[229] vdd vss bl[229] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_230 br[229] vdd vss bl[229] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_231 br[230] vdd vss bl[230] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_231 br[230] vdd vss bl[230] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_232 br[231] vdd vss bl[231] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_232 br[231] vdd vss bl[231] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_233 br[232] vdd vss bl[232] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_233 br[232] vdd vss bl[232] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_234 br[233] vdd vss bl[233] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_234 br[233] vdd vss bl[233] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_235 br[234] vdd vss bl[234] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_235 br[234] vdd vss bl[234] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_236 br[235] vdd vss bl[235] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_236 br[235] vdd vss bl[235] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_237 br[236] vdd vss bl[236] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_237 br[236] vdd vss bl[236] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_238 br[237] vdd vss bl[237] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_238 br[237] vdd vss bl[237] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_239 br[238] vdd vss bl[238] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_239 br[238] vdd vss bl[238] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_240 br[239] vdd vss bl[239] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_240 br[239] vdd vss bl[239] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_241 br[240] vdd vss bl[240] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_241 br[240] vdd vss bl[240] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_242 br[241] vdd vss bl[241] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_242 br[241] vdd vss bl[241] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_243 br[242] vdd vss bl[242] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_243 br[242] vdd vss bl[242] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_244 br[243] vdd vss bl[243] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_244 br[243] vdd vss bl[243] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_245 br[244] vdd vss bl[244] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_245 br[244] vdd vss bl[244] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_246 br[245] vdd vss bl[245] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_246 br[245] vdd vss bl[245] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_247 br[246] vdd vss bl[246] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_247 br[246] vdd vss bl[246] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_248 br[247] vdd vss bl[247] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_248 br[247] vdd vss bl[247] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_249 br[248] vdd vss bl[248] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_249 br[248] vdd vss bl[248] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_250 br[249] vdd vss bl[249] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_250 br[249] vdd vss bl[249] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_251 br[250] vdd vss bl[250] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_251 br[250] vdd vss bl[250] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_252 br[251] vdd vss bl[251] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_252 br[251] vdd vss bl[251] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_253 br[252] vdd vss bl[252] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_253 br[252] vdd vss bl[252] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_254 br[253] vdd vss bl[253] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_254 br[253] vdd vss bl[253] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_255 br[254] vdd vss bl[254] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_255 br[254] vdd vss bl[254] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_256 br[255] vdd vss bl[255] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_256 br[255] vdd vss bl[255] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_257 vdd vdd vss vdd vss vdd sram_sp_colend_wrapper
  Xcolend_bot_257 vdd vdd vss vdd vss vdd sram_sp_colend_wrapper
  Xhstrap_0_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_257 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhoriz_wlstrap_0_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper

.ENDS sp_cell_array

.SUBCKT sky130_fd_sc_hs__inv_4 A VGND VNB VPB VPWR Y

  X0 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X4 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X7 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__inv_4

.SUBCKT sky130_fd_sc_hs__inv_4_wrapper A VGND VNB VPB VPWR Y

  X0 A VGND VNB VPB VPWR Y sky130_fd_sc_hs__inv_4

.ENDS sky130_fd_sc_hs__inv_4_wrapper

.SUBCKT mos_w3550_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=3.550


.ENDS mos_w3550_l150_m1_nf1_id1

.SUBCKT mos_w3200_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=3.200


.ENDS mos_w3200_l150_m1_nf1_id1

.SUBCKT mos_w1280_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.280


.ENDS mos_w1280_l150_m1_nf1_id0

.SUBCKT folded_inv_10 vdd vss a y

  XMP0 y a vdd vdd mos_w3200_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w1280_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w3200_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w1280_l150_m1_nf1_id0

.ENDS folded_inv_10

.SUBCKT decoder_stage_10 vdd vss y[0] y[1] y[2] y[3] y_b[0] y_b[1] y_b[2] y_b[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1

  Xgate_0_0_0 vdd vss predecode_0_0 predecode_1_0 y_b[0] nand2_1
  Xgate_0_1_0 vdd vss predecode_0_1 predecode_1_0 y_b[1] nand2_1
  Xgate_0_2_0 vdd vss predecode_0_0 predecode_1_1 y_b[2] nand2_1
  Xgate_0_3_0 vdd vss predecode_0_1 predecode_1_1 y_b[3] nand2_1
  Xgate_1_0_0 vdd vss y_b[0] y[0] folded_inv_10
  Xgate_1_1_0 vdd vss y_b[1] y[1] folded_inv_10
  Xgate_1_2_0 vdd vss y_b[2] y[2] folded_inv_10
  Xgate_1_3_0 vdd vss y_b[3] y[3] folded_inv_10

.ENDS decoder_stage_10

.SUBCKT decoder_4 vdd vss y[0] y[1] y[2] y[3] y_b[0] y_b[1] y_b[2] y_b[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1

  X0 vdd vss y[0] y[1] y[2] y[3] y_b[0] y_b[1] y_b[2] y_b[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 decoder_stage_10

.ENDS decoder_4

.SUBCKT mos_w2850_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=2.850


.ENDS mos_w2850_l150_m1_nf1_id0

.SUBCKT nand2_2 vdd vss a b y

  Xn1 x a vss vss mos_w2850_l150_m1_nf1_id0
  Xn2 y b x vss mos_w2850_l150_m1_nf1_id0
  Xp1 y a vdd vdd mos_w3550_l150_m1_nf1_id1
  Xp2 y b vdd vdd mos_w3550_l150_m1_nf1_id1

.ENDS nand2_2

.SUBCKT mos_w2270_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.270


.ENDS mos_w2270_l150_m1_nf1_id1

.SUBCKT mos_w900_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.900


.ENDS mos_w900_l150_m1_nf1_id0

.SUBCKT folded_inv_6 vdd vss a y

  XMP0 y a vdd vdd mos_w2270_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w900_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w2270_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w900_l150_m1_nf1_id0

.ENDS folded_inv_6

.SUBCKT decoder_stage_8 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y[12] y[13] y[14] y[15] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] y_b[12] y_b[13] y_b[14] y_b[15] predecode_0_0 predecode_0_1 predecode_0_2 predecode_0_3 predecode_1_0 predecode_1_1 predecode_1_2 predecode_1_3

  Xgate_0_0_0 vdd vss predecode_0_0 predecode_1_0 y_b[0] nand2_2
  Xgate_0_1_0 vdd vss predecode_0_1 predecode_1_0 y_b[1] nand2_2
  Xgate_0_2_0 vdd vss predecode_0_2 predecode_1_0 y_b[2] nand2_2
  Xgate_0_3_0 vdd vss predecode_0_3 predecode_1_0 y_b[3] nand2_2
  Xgate_0_4_0 vdd vss predecode_0_0 predecode_1_1 y_b[4] nand2_2
  Xgate_0_5_0 vdd vss predecode_0_1 predecode_1_1 y_b[5] nand2_2
  Xgate_0_6_0 vdd vss predecode_0_2 predecode_1_1 y_b[6] nand2_2
  Xgate_0_7_0 vdd vss predecode_0_3 predecode_1_1 y_b[7] nand2_2
  Xgate_0_8_0 vdd vss predecode_0_0 predecode_1_2 y_b[8] nand2_2
  Xgate_0_9_0 vdd vss predecode_0_1 predecode_1_2 y_b[9] nand2_2
  Xgate_0_10_0 vdd vss predecode_0_2 predecode_1_2 y_b[10] nand2_2
  Xgate_0_11_0 vdd vss predecode_0_3 predecode_1_2 y_b[11] nand2_2
  Xgate_0_12_0 vdd vss predecode_0_0 predecode_1_3 y_b[12] nand2_2
  Xgate_0_13_0 vdd vss predecode_0_1 predecode_1_3 y_b[13] nand2_2
  Xgate_0_14_0 vdd vss predecode_0_2 predecode_1_3 y_b[14] nand2_2
  Xgate_0_15_0 vdd vss predecode_0_3 predecode_1_3 y_b[15] nand2_2
  Xgate_1_0_0 vdd vss y_b[0] y[0] folded_inv_6
  Xgate_1_0_1 vdd vss y_b[0] y[0] folded_inv_6
  Xgate_1_1_0 vdd vss y_b[1] y[1] folded_inv_6
  Xgate_1_1_1 vdd vss y_b[1] y[1] folded_inv_6
  Xgate_1_2_0 vdd vss y_b[2] y[2] folded_inv_6
  Xgate_1_2_1 vdd vss y_b[2] y[2] folded_inv_6
  Xgate_1_3_0 vdd vss y_b[3] y[3] folded_inv_6
  Xgate_1_3_1 vdd vss y_b[3] y[3] folded_inv_6
  Xgate_1_4_0 vdd vss y_b[4] y[4] folded_inv_6
  Xgate_1_4_1 vdd vss y_b[4] y[4] folded_inv_6
  Xgate_1_5_0 vdd vss y_b[5] y[5] folded_inv_6
  Xgate_1_5_1 vdd vss y_b[5] y[5] folded_inv_6
  Xgate_1_6_0 vdd vss y_b[6] y[6] folded_inv_6
  Xgate_1_6_1 vdd vss y_b[6] y[6] folded_inv_6
  Xgate_1_7_0 vdd vss y_b[7] y[7] folded_inv_6
  Xgate_1_7_1 vdd vss y_b[7] y[7] folded_inv_6
  Xgate_1_8_0 vdd vss y_b[8] y[8] folded_inv_6
  Xgate_1_8_1 vdd vss y_b[8] y[8] folded_inv_6
  Xgate_1_9_0 vdd vss y_b[9] y[9] folded_inv_6
  Xgate_1_9_1 vdd vss y_b[9] y[9] folded_inv_6
  Xgate_1_10_0 vdd vss y_b[10] y[10] folded_inv_6
  Xgate_1_10_1 vdd vss y_b[10] y[10] folded_inv_6
  Xgate_1_11_0 vdd vss y_b[11] y[11] folded_inv_6
  Xgate_1_11_1 vdd vss y_b[11] y[11] folded_inv_6
  Xgate_1_12_0 vdd vss y_b[12] y[12] folded_inv_6
  Xgate_1_12_1 vdd vss y_b[12] y[12] folded_inv_6
  Xgate_1_13_0 vdd vss y_b[13] y[13] folded_inv_6
  Xgate_1_13_1 vdd vss y_b[13] y[13] folded_inv_6
  Xgate_1_14_0 vdd vss y_b[14] y[14] folded_inv_6
  Xgate_1_14_1 vdd vss y_b[14] y[14] folded_inv_6
  Xgate_1_15_0 vdd vss y_b[15] y[15] folded_inv_6
  Xgate_1_15_1 vdd vss y_b[15] y[15] folded_inv_6

.ENDS decoder_stage_8

.SUBCKT decoder_2 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y[12] y[13] y[14] y[15] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] y_b[12] y_b[13] y_b[14] y_b[15] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 predecode_2_0 predecode_2_1 predecode_3_0 predecode_3_1

  X0 vdd vss child_conn_0[0] child_conn_0[1] child_conn_0[2] child_conn_0[3] child_noconn_0[0] child_noconn_0[1] child_noconn_0[2] child_noconn_0[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 decoder_4
  X0_1 vdd vss child_conn_1[0] child_conn_1[1] child_conn_1[2] child_conn_1[3] child_noconn_1[0] child_noconn_1[1] child_noconn_1[2] child_noconn_1[3] predecode_2_0 predecode_2_1 predecode_3_0 predecode_3_1 decoder_4
  X0_2 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y[12] y[13] y[14] y[15] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] y_b[12] y_b[13] y_b[14] y_b[15] child_conn_0[0] child_conn_0[1] child_conn_0[2] child_conn_0[3] child_conn_1[0] child_conn_1[1] child_conn_1[2] child_conn_1[3] decoder_stage_8

.ENDS decoder_2

.SUBCKT mos_w3000_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=3.000


.ENDS mos_w3000_l150_m1_nf1_id0

.SUBCKT nand3 vdd vss a b c y

  Xn1 x1 a vss vss mos_w3000_l150_m1_nf1_id0
  Xn2 x2 b x1 vss mos_w3000_l150_m1_nf1_id0
  Xn3 y c x2 vss mos_w3000_l150_m1_nf1_id0
  Xp1 y a vdd vdd mos_w2500_l150_m1_nf1_id1
  Xp2 y b vdd vdd mos_w2500_l150_m1_nf1_id1
  Xp3 y c vdd vdd mos_w2500_l150_m1_nf1_id1

.ENDS nand3

.SUBCKT mos_w2690_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.690


.ENDS mos_w2690_l150_m1_nf1_id1

.SUBCKT mos_w1080_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.080


.ENDS mos_w1080_l150_m1_nf1_id0

.SUBCKT folded_inv_7 vdd vss a y

  XMP0 y a vdd vdd mos_w2690_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w1080_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w2690_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w1080_l150_m1_nf1_id0

.ENDS folded_inv_7

.SUBCKT decoder_stage_9 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 predecode_2_0 predecode_2_1

  Xgate_0_0_0 vdd vss predecode_0_0 predecode_1_0 predecode_2_0 y_b[0] nand3
  Xgate_0_1_0 vdd vss predecode_0_1 predecode_1_0 predecode_2_0 y_b[1] nand3
  Xgate_0_2_0 vdd vss predecode_0_0 predecode_1_1 predecode_2_0 y_b[2] nand3
  Xgate_0_3_0 vdd vss predecode_0_1 predecode_1_1 predecode_2_0 y_b[3] nand3
  Xgate_0_4_0 vdd vss predecode_0_0 predecode_1_0 predecode_2_1 y_b[4] nand3
  Xgate_0_5_0 vdd vss predecode_0_1 predecode_1_0 predecode_2_1 y_b[5] nand3
  Xgate_0_6_0 vdd vss predecode_0_0 predecode_1_1 predecode_2_1 y_b[6] nand3
  Xgate_0_7_0 vdd vss predecode_0_1 predecode_1_1 predecode_2_1 y_b[7] nand3
  Xgate_1_0_0 vdd vss y_b[0] y[0] folded_inv_7
  Xgate_1_0_1 vdd vss y_b[0] y[0] folded_inv_7
  Xgate_1_1_0 vdd vss y_b[1] y[1] folded_inv_7
  Xgate_1_1_1 vdd vss y_b[1] y[1] folded_inv_7
  Xgate_1_2_0 vdd vss y_b[2] y[2] folded_inv_7
  Xgate_1_2_1 vdd vss y_b[2] y[2] folded_inv_7
  Xgate_1_3_0 vdd vss y_b[3] y[3] folded_inv_7
  Xgate_1_3_1 vdd vss y_b[3] y[3] folded_inv_7
  Xgate_1_4_0 vdd vss y_b[4] y[4] folded_inv_7
  Xgate_1_4_1 vdd vss y_b[4] y[4] folded_inv_7
  Xgate_1_5_0 vdd vss y_b[5] y[5] folded_inv_7
  Xgate_1_5_1 vdd vss y_b[5] y[5] folded_inv_7
  Xgate_1_6_0 vdd vss y_b[6] y[6] folded_inv_7
  Xgate_1_6_1 vdd vss y_b[6] y[6] folded_inv_7
  Xgate_1_7_0 vdd vss y_b[7] y[7] folded_inv_7
  Xgate_1_7_1 vdd vss y_b[7] y[7] folded_inv_7

.ENDS decoder_stage_9

.SUBCKT decoder_3 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 predecode_2_0 predecode_2_1

  X0 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 predecode_2_0 predecode_2_1 decoder_stage_9

.ENDS decoder_3

.SUBCKT decoder vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y[12] y[13] y[14] y[15] y[16] y[17] y[18] y[19] y[20] y[21] y[22] y[23] y[24] y[25] y[26] y[27] y[28] y[29] y[30] y[31] y[32] y[33] y[34] y[35] y[36] y[37] y[38] y[39] y[40] y[41] y[42] y[43] y[44] y[45] y[46] y[47] y[48] y[49] y[50] y[51] y[52] y[53] y[54] y[55] y[56] y[57] y[58] y[59] y[60] y[61] y[62] y[63] y[64] y[65] y[66] y[67] y[68] y[69] y[70] y[71] y[72] y[73] y[74] y[75] y[76] y[77] y[78] y[79] y[80] y[81] y[82] y[83] y[84] y[85] y[86] y[87] y[88] y[89] y[90] y[91] y[92] y[93] y[94] y[95] y[96] y[97] y[98] y[99] y[100] y[101] y[102] y[103] y[104] y[105] y[106] y[107] y[108] y[109] y[110] y[111] y[112] y[113] y[114] y[115] y[116] y[117] y[118] y[119] y[120] y[121] y[122] y[123] y[124] y[125] y[126] y[127] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] y_b[12] y_b[13] y_b[14] y_b[15] y_b[16] y_b[17] y_b[18] y_b[19] y_b[20] y_b[21] y_b[22] y_b[23] y_b[24] y_b[25] y_b[26] y_b[27] y_b[28] y_b[29] y_b[30] y_b[31] y_b[32] y_b[33] y_b[34] y_b[35] y_b[36] y_b[37] y_b[38] y_b[39] y_b[40] y_b[41] y_b[42] y_b[43] y_b[44] y_b[45] y_b[46] y_b[47] y_b[48] y_b[49] y_b[50] y_b[51] y_b[52] y_b[53] y_b[54] y_b[55] y_b[56] y_b[57] y_b[58] y_b[59] y_b[60] y_b[61] y_b[62] y_b[63] y_b[64] y_b[65] y_b[66] y_b[67] y_b[68] y_b[69] y_b[70] y_b[71] y_b[72] y_b[73] y_b[74] y_b[75] y_b[76] y_b[77] y_b[78] y_b[79] y_b[80] y_b[81] y_b[82] y_b[83] y_b[84] y_b[85] y_b[86] y_b[87] y_b[88] y_b[89] y_b[90] y_b[91] y_b[92] y_b[93] y_b[94] y_b[95] y_b[96] y_b[97] y_b[98] y_b[99] y_b[100] y_b[101] y_b[102] y_b[103] y_b[104] y_b[105] y_b[106] y_b[107] y_b[108] y_b[109] y_b[110] y_b[111] y_b[112] y_b[113] y_b[114] y_b[115] y_b[116] y_b[117] y_b[118] y_b[119] y_b[120] y_b[121] y_b[122] y_b[123] y_b[124] y_b[125] y_b[126] y_b[127] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 predecode_2_0 predecode_2_1 predecode_3_0 predecode_3_1 predecode_4_0 predecode_4_1 predecode_5_0 predecode_5_1 predecode_6_0 predecode_6_1

  X0 vdd vss child_conn_0[0] child_conn_0[1] child_conn_0[2] child_conn_0[3] child_conn_0[4] child_conn_0[5] child_conn_0[6] child_conn_0[7] child_conn_0[8] child_conn_0[9] child_conn_0[10] child_conn_0[11] child_conn_0[12] child_conn_0[13] child_conn_0[14] child_conn_0[15] child_noconn_0[0] child_noconn_0[1] child_noconn_0[2] child_noconn_0[3] child_noconn_0[4] child_noconn_0[5] child_noconn_0[6] child_noconn_0[7] child_noconn_0[8] child_noconn_0[9] child_noconn_0[10] child_noconn_0[11] child_noconn_0[12] child_noconn_0[13] child_noconn_0[14] child_noconn_0[15] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 predecode_2_0 predecode_2_1 predecode_3_0 predecode_3_1 decoder_2
  X0_1 vdd vss child_conn_1[0] child_conn_1[1] child_conn_1[2] child_conn_1[3] child_conn_1[4] child_conn_1[5] child_conn_1[6] child_conn_1[7] child_noconn_1[0] child_noconn_1[1] child_noconn_1[2] child_noconn_1[3] child_noconn_1[4] child_noconn_1[5] child_noconn_1[6] child_noconn_1[7] predecode_4_0 predecode_4_1 predecode_5_0 predecode_5_1 predecode_6_0 predecode_6_1 decoder_3
  X0_2 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y[12] y[13] y[14] y[15] y[16] y[17] y[18] y[19] y[20] y[21] y[22] y[23] y[24] y[25] y[26] y[27] y[28] y[29] y[30] y[31] y[32] y[33] y[34] y[35] y[36] y[37] y[38] y[39] y[40] y[41] y[42] y[43] y[44] y[45] y[46] y[47] y[48] y[49] y[50] y[51] y[52] y[53] y[54] y[55] y[56] y[57] y[58] y[59] y[60] y[61] y[62] y[63] y[64] y[65] y[66] y[67] y[68] y[69] y[70] y[71] y[72] y[73] y[74] y[75] y[76] y[77] y[78] y[79] y[80] y[81] y[82] y[83] y[84] y[85] y[86] y[87] y[88] y[89] y[90] y[91] y[92] y[93] y[94] y[95] y[96] y[97] y[98] y[99] y[100] y[101] y[102] y[103] y[104] y[105] y[106] y[107] y[108] y[109] y[110] y[111] y[112] y[113] y[114] y[115] y[116] y[117] y[118] y[119] y[120] y[121] y[122] y[123] y[124] y[125] y[126] y[127] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] y_b[12] y_b[13] y_b[14] y_b[15] y_b[16] y_b[17] y_b[18] y_b[19] y_b[20] y_b[21] y_b[22] y_b[23] y_b[24] y_b[25] y_b[26] y_b[27] y_b[28] y_b[29] y_b[30] y_b[31] y_b[32] y_b[33] y_b[34] y_b[35] y_b[36] y_b[37] y_b[38] y_b[39] y_b[40] y_b[41] y_b[42] y_b[43] y_b[44] y_b[45] y_b[46] y_b[47] y_b[48] y_b[49] y_b[50] y_b[51] y_b[52] y_b[53] y_b[54] y_b[55] y_b[56] y_b[57] y_b[58] y_b[59] y_b[60] y_b[61] y_b[62] y_b[63] y_b[64] y_b[65] y_b[66] y_b[67] y_b[68] y_b[69] y_b[70] y_b[71] y_b[72] y_b[73] y_b[74] y_b[75] y_b[76] y_b[77] y_b[78] y_b[79] y_b[80] y_b[81] y_b[82] y_b[83] y_b[84] y_b[85] y_b[86] y_b[87] y_b[88] y_b[89] y_b[90] y_b[91] y_b[92] y_b[93] y_b[94] y_b[95] y_b[96] y_b[97] y_b[98] y_b[99] y_b[100] y_b[101] y_b[102] y_b[103] y_b[104] y_b[105] y_b[106] y_b[107] y_b[108] y_b[109] y_b[110] y_b[111] y_b[112] y_b[113] y_b[114] y_b[115] y_b[116] y_b[117] y_b[118] y_b[119] y_b[120] y_b[121] y_b[122] y_b[123] y_b[124] y_b[125] y_b[126] y_b[127] child_conn_0[0] child_conn_0[1] child_conn_0[2] child_conn_0[3] child_conn_0[4] child_conn_0[5] child_conn_0[6] child_conn_0[7] child_conn_0[8] child_conn_0[9] child_conn_0[10] child_conn_0[11] child_conn_0[12] child_conn_0[13] child_conn_0[14] child_conn_0[15] child_conn_1[0] child_conn_1[1] child_conn_1[2] child_conn_1[3] child_conn_1[4] child_conn_1[5] child_conn_1[6] child_conn_1[7] decoder_stage_5

.ENDS decoder

.SUBCKT sky130_fd_sc_hs__dfrbp_2 CLK D RESET_B VGND VNB VPB VPWR Q Q_N

  X0 a_1800_291# a_1586_149# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X1 VGND CLK a_728_331# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X2 Q a_2363_352# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X3 VPWR CLK a_728_331# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X4 a_1499_149# a_728_331# a_1586_149# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X5 a_536_81# a_331_392# a_614_81# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X6 a_156_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X7 a_298_294# a_818_418# a_614_81# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X8 a_70_74# a_728_331# a_298_294# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X9 a_331_392# a_728_331# a_1586_149# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X10 a_70_74# D a_156_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X11 a_818_418# a_728_331# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X12 a_818_418# a_728_331# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X13 a_1586_149# a_818_418# a_1755_389# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X14 Q_N a_1586_149# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X15 a_298_294# a_818_418# a_70_74# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X16 VGND RESET_B a_536_81# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X17 a_1755_389# a_1800_291# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X18 a_1586_149# a_818_418# a_331_392# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X19 Q a_2363_352# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X20 VGND a_1586_149# Q_N VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X21 VGND a_1586_149# a_2363_352# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X22 VPWR a_298_294# a_331_392# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X23 a_298_294# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X24 a_1499_149# a_1800_291# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X25 VPWR a_331_392# a_683_485# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X26 VPWR D a_70_74# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X27 VPWR RESET_B a_1800_291# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X28 a_1974_74# a_1586_149# a_1800_291# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X29 a_70_74# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X30 Q_N a_1586_149# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X31 VPWR a_1586_149# a_2363_352# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X32 VGND a_2363_352# Q VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X33 VPWR a_1586_149# Q_N VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X34 VGND RESET_B a_1974_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X35 a_683_485# a_728_331# a_298_294# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X36 VGND a_298_294# a_331_392# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X37 VPWR a_2363_352# Q VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120


.ENDS sky130_fd_sc_hs__dfrbp_2

.SUBCKT sky130_fd_sc_hs__dfrbp_2_wrapper CLK D RESET_B VGND VNB VPB VPWR Q Q_N

  X0 CLK D RESET_B VGND VNB VPB VPWR Q Q_N sky130_fd_sc_hs__dfrbp_2

.ENDS sky130_fd_sc_hs__dfrbp_2_wrapper

.SUBCKT dff_array_11 vdd vss clk rb d[0] d[1] d[2] d[3] d[4] d[5] d[6] d[7] d[8] d[9] d[10] q[0] q[1] q[2] q[3] q[4] q[5] q[6] q[7] q[8] q[9] q[10] qn[0] qn[1] qn[2] qn[3] qn[4] qn[5] qn[6] qn[7] qn[8] qn[9] qn[10]

  Xdff_0 clk d[0] rb vss vss vdd vdd q[0] qn[0] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_1 clk d[1] rb vss vss vdd vdd q[1] qn[1] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_2 clk d[2] rb vss vss vdd vdd q[2] qn[2] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_3 clk d[3] rb vss vss vdd vdd q[3] qn[3] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_4 clk d[4] rb vss vss vdd vdd q[4] qn[4] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_5 clk d[5] rb vss vss vdd vdd q[5] qn[5] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_6 clk d[6] rb vss vss vdd vdd q[6] qn[6] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_7 clk d[7] rb vss vss vdd vdd q[7] qn[7] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_8 clk d[8] rb vss vss vdd vdd q[8] qn[8] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_9 clk d[9] rb vss vss vdd vdd q[9] qn[9] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_10 clk d[10] rb vss vss vdd vdd q[10] qn[10] sky130_fd_sc_hs__dfrbp_2_wrapper

.ENDS dff_array_11

.SUBCKT mos_w2480_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.480


.ENDS mos_w2480_l150_m1_nf1_id1

.SUBCKT mos_w1000_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.000


.ENDS mos_w1000_l150_m1_nf1_id0

.SUBCKT folded_inv_2 vdd vss a y

  XMP0 y a vdd vdd mos_w2480_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w1000_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w2480_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w1000_l150_m1_nf1_id0

.ENDS folded_inv_2

.SUBCKT sky130_fd_sc_hs__inv_2 A VGND VNB VPB VPWR Y

  X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X3 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__inv_2

.SUBCKT sky130_fd_sc_hs__inv_2_wrapper A VGND VNB VPB VPWR Y

  X0 A VGND VNB VPB VPWR Y sky130_fd_sc_hs__inv_2

.ENDS sky130_fd_sc_hs__inv_2_wrapper

.SUBCKT mos_w3000_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=3.000


.ENDS mos_w3000_l150_m1_nf1_id1

.SUBCKT mos_w7050_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=7.050


.ENDS mos_w7050_l150_m1_nf1_id1

.SUBCKT mos_w600_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.600


.ENDS mos_w600_l150_m1_nf1_id0

.SUBCKT sky130_fd_sc_hs__nor2_4 A B VGND VNB VPB VPWR Y

  X0 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 a_27_368# B Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X3 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X4 Y B a_27_368# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X5 a_27_368# B Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X6 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X7 VPWR A a_27_368# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X8 VPWR A a_27_368# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X11 Y B a_27_368# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120


.ENDS sky130_fd_sc_hs__nor2_4

.SUBCKT sky130_fd_sc_hs__nor2_4_wrapper A B VGND VNB VPB VPWR Y

  X0 A B VGND VNB VPB VPWR Y sky130_fd_sc_hs__nor2_4

.ENDS sky130_fd_sc_hs__nor2_4_wrapper

.SUBCKT sky130_fd_sc_hs__inv_16 A VGND VNB VPB VPWR Y

  X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X5 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X7 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X11 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X13 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X14 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X15 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X16 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X17 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X18 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X19 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X20 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X21 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X22 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X23 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X24 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X25 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X26 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X27 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X28 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X30 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X31 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120


.ENDS sky130_fd_sc_hs__inv_16

.SUBCKT sky130_fd_sc_hs__nand2_4 A B VGND VNB VPB VPWR Y

  X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X2 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X3 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X4 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X5 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X6 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X8 Y B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X11 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__nand2_4

.SUBCKT sky130_fd_sc_hs__nand2_4_wrapper A B VGND VNB VPB VPWR Y

  X0 A B VGND VNB VPB VPWR Y sky130_fd_sc_hs__nand2_4

.ENDS sky130_fd_sc_hs__nand2_4_wrapper

.SUBCKT mos_w5000_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=5.000


.ENDS mos_w5000_l150_m1_nf1_id1

.SUBCKT folded_inv_1 vdd vss a y

  XMP0 y a vdd vdd mos_w5000_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w2000_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w5000_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w2000_l150_m1_nf1_id0

.ENDS folded_inv_1

.SUBCKT sky130_fd_sc_hs__and2_2 A B VGND VNB VPB VPWR X

  X0 a_31_74# B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X1 X a_31_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X2 X a_31_74# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 a_118_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X4 a_31_74# A a_118_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X5 VPWR A a_31_74# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X6 VPWR a_31_74# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X7 VGND a_31_74# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__and2_2

.SUBCKT sky130_fd_sc_hs__and2_4 A B VGND VNB VPB VPWR X

  X0 VPWR a_83_269# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 VPWR B a_83_269# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.840

  X2 VPWR a_83_269# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 a_504_119# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X4 a_83_269# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.840

  X5 VGND B a_504_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X6 VGND a_83_269# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X7 a_83_269# B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.840

  X8 X a_83_269# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 VGND a_83_269# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 X a_83_269# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X11 X a_83_269# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X12 a_504_119# A a_83_269# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X13 a_83_269# A a_504_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X14 VPWR A a_83_269# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.840

  X15 X a_83_269# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__and2_4

.SUBCKT multi_finger_inv vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv

.SUBCKT and2 vdd a b y yb vss

  X0 vdd vss a b yb nand2
  X0_1 vdd vss yb y folded_inv_1

.ENDS and2

.SUBCKT decoder_stage vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y[12] y[13] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] y_b[12] y_b[13] wl_en in[0] in[1] in[2] in[3] in[4] in[5] in[6] in[7] in[8] in[9] in[10] in[11] in[12] in[13]

  Xgate_0_0_0 vdd wl_en in[0] y[0] y_b[0] vss and2
  Xgate_0_1_0 vdd wl_en in[1] y[1] y_b[1] vss and2
  Xgate_0_2_0 vdd wl_en in[2] y[2] y_b[2] vss and2
  Xgate_0_3_0 vdd wl_en in[3] y[3] y_b[3] vss and2
  Xgate_0_4_0 vdd wl_en in[4] y[4] y_b[4] vss and2
  Xgate_0_5_0 vdd wl_en in[5] y[5] y_b[5] vss and2
  Xgate_0_6_0 vdd wl_en in[6] y[6] y_b[6] vss and2
  Xgate_0_7_0 vdd wl_en in[7] y[7] y_b[7] vss and2
  Xgate_0_8_0 vdd wl_en in[8] y[8] y_b[8] vss and2
  Xgate_0_9_0 vdd wl_en in[9] y[9] y_b[9] vss and2
  Xgate_0_10_0 vdd wl_en in[10] y[10] y_b[10] vss and2
  Xgate_0_11_0 vdd wl_en in[11] y[11] y_b[11] vss and2
  Xgate_0_12_0 vdd wl_en in[12] y[12] y_b[12] vss and2
  Xgate_0_13_0 vdd wl_en in[13] y[13] y_b[13] vss and2

.ENDS decoder_stage

.SUBCKT sky130_fd_sc_hs__inv_16_wrapper A VGND VNB VPB VPWR Y

  X0 A VGND VNB VPB VPWR Y sky130_fd_sc_hs__inv_16

.ENDS sky130_fd_sc_hs__inv_16_wrapper

.SUBCKT inv_chain_12 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sky130_fd_sc_hs__inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd x[2] sky130_fd_sc_hs__inv_2_wrapper
  Xinv3 x[2] vss vss vdd vdd x[3] sky130_fd_sc_hs__inv_2_wrapper
  Xinv4 x[3] vss vss vdd vdd x[4] sky130_fd_sc_hs__inv_2_wrapper
  Xinv5 x[4] vss vss vdd vdd x[5] sky130_fd_sc_hs__inv_2_wrapper
  Xinv6 x[5] vss vss vdd vdd x[6] sky130_fd_sc_hs__inv_2_wrapper
  Xinv7 x[6] vss vss vdd vdd x[7] sky130_fd_sc_hs__inv_2_wrapper
  Xinv8 x[7] vss vss vdd vdd x[8] sky130_fd_sc_hs__inv_2_wrapper
  Xinv9 x[8] vss vss vdd vdd x[9] sky130_fd_sc_hs__inv_2_wrapper
  Xinv10 x[9] vss vss vdd vdd x[10] sky130_fd_sc_hs__inv_2_wrapper
  Xinv11 x[10] vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_12

.SUBCKT sky130_fd_sc_hs__and2_2_wrapper A B VGND VNB VPB VPWR X

  X0 A B VGND VNB VPB VPWR X sky130_fd_sc_hs__and2_2

.ENDS sky130_fd_sc_hs__and2_2_wrapper

.SUBCKT inv_chain_9 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sky130_fd_sc_hs__inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd x[2] sky130_fd_sc_hs__inv_2_wrapper
  Xinv3 x[2] vss vss vdd vdd x[3] sky130_fd_sc_hs__inv_2_wrapper
  Xinv4 x[3] vss vss vdd vdd x[4] sky130_fd_sc_hs__inv_2_wrapper
  Xinv5 x[4] vss vss vdd vdd x[5] sky130_fd_sc_hs__inv_2_wrapper
  Xinv6 x[5] vss vss vdd vdd x[6] sky130_fd_sc_hs__inv_2_wrapper
  Xinv7 x[6] vss vss vdd vdd x[7] sky130_fd_sc_hs__inv_2_wrapper
  Xinv8 x[7] vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_9

.SUBCKT sky130_fd_sc_hs__and2_4_wrapper A B VGND VNB VPB VPWR X

  X0 A B VGND VNB VPB VPWR X sky130_fd_sc_hs__and2_4

.ENDS sky130_fd_sc_hs__and2_4_wrapper

.SUBCKT edge_detector din dout vdd vss

  Xdelay_chain din delayed vdd vss inv_chain_9
  Xand din delayed vss vss vdd vdd dout sky130_fd_sc_hs__and2_4_wrapper

.ENDS edge_detector

.SUBCKT sky130_fd_sc_hs__buf_16 A VGND VNB VPB VPWR X

  X0 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X3 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X4 VPWR A a_83_260# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X5 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X6 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X7 VPWR A a_83_260# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X8 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X9 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 VPWR A a_83_260# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X11 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X12 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X13 a_83_260# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X14 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X15 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X16 VGND A a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X17 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X18 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X19 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X20 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X21 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X22 VGND A a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X23 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X24 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X25 a_83_260# A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X26 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X27 a_83_260# A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X28 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X29 a_83_260# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X30 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X31 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X32 a_83_260# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X33 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X34 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X35 a_83_260# A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X36 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X37 VGND A a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X38 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X39 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X40 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X41 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X42 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X43 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__buf_16

.SUBCKT sky130_fd_sc_hs__buf_16_wrapper A VGND VNB VPB VPWR X

  X0 A VGND VNB VPB VPWR X sky130_fd_sc_hs__buf_16

.ENDS sky130_fd_sc_hs__buf_16_wrapper

.SUBCKT inv_chain_3 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sky130_fd_sc_hs__inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_3

.SUBCKT inv_chain_15 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sky130_fd_sc_hs__inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd x[2] sky130_fd_sc_hs__inv_2_wrapper
  Xinv3 x[2] vss vss vdd vdd x[3] sky130_fd_sc_hs__inv_2_wrapper
  Xinv4 x[3] vss vss vdd vdd x[4] sky130_fd_sc_hs__inv_2_wrapper
  Xinv5 x[4] vss vss vdd vdd x[5] sky130_fd_sc_hs__inv_2_wrapper
  Xinv6 x[5] vss vss vdd vdd x[6] sky130_fd_sc_hs__inv_2_wrapper
  Xinv7 x[6] vss vss vdd vdd x[7] sky130_fd_sc_hs__inv_2_wrapper
  Xinv8 x[7] vss vss vdd vdd x[8] sky130_fd_sc_hs__inv_2_wrapper
  Xinv9 x[8] vss vss vdd vdd x[9] sky130_fd_sc_hs__inv_2_wrapper
  Xinv10 x[9] vss vss vdd vdd x[10] sky130_fd_sc_hs__inv_2_wrapper
  Xinv11 x[10] vss vss vdd vdd x[11] sky130_fd_sc_hs__inv_2_wrapper
  Xinv12 x[11] vss vss vdd vdd x[12] sky130_fd_sc_hs__inv_2_wrapper
  Xinv13 x[12] vss vss vdd vdd x[13] sky130_fd_sc_hs__inv_2_wrapper
  Xinv14 x[13] vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_15

.SUBCKT sramgen_svt_inv_2 A VGND VNB VPB VPWR Y

  X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740

  X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740


.ENDS sramgen_svt_inv_2

.SUBCKT sramgen_svt_inv_2_wrapper A VGND VNB VPB VPWR Y

  X0 A VGND VNB VPB VPWR Y sramgen_svt_inv_2

.ENDS sramgen_svt_inv_2_wrapper

.SUBCKT sramgen_svt_inv_4 A VGND VNB VPB VPWR Y

  X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740

  X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740

  X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740

  X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740


.ENDS sramgen_svt_inv_4

.SUBCKT sramgen_svt_inv_4_wrapper A VGND VNB VPB VPWR Y

  X0 A VGND VNB VPB VPWR Y sramgen_svt_inv_4

.ENDS sramgen_svt_inv_4_wrapper

.SUBCKT svt_inv_chain_28 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sramgen_svt_inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sramgen_svt_inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd x[2] sramgen_svt_inv_2_wrapper
  Xinv3 x[2] vss vss vdd vdd x[3] sramgen_svt_inv_2_wrapper
  Xinv4 x[3] vss vss vdd vdd x[4] sramgen_svt_inv_2_wrapper
  Xinv5 x[4] vss vss vdd vdd x[5] sramgen_svt_inv_2_wrapper
  Xinv6 x[5] vss vss vdd vdd x[6] sramgen_svt_inv_2_wrapper
  Xinv7 x[6] vss vss vdd vdd x[7] sramgen_svt_inv_2_wrapper
  Xinv8 x[7] vss vss vdd vdd x[8] sramgen_svt_inv_2_wrapper
  Xinv9 x[8] vss vss vdd vdd x[9] sramgen_svt_inv_2_wrapper
  Xinv10 x[9] vss vss vdd vdd x[10] sramgen_svt_inv_2_wrapper
  Xinv11 x[10] vss vss vdd vdd x[11] sramgen_svt_inv_2_wrapper
  Xinv12 x[11] vss vss vdd vdd x[12] sramgen_svt_inv_2_wrapper
  Xinv13 x[12] vss vss vdd vdd x[13] sramgen_svt_inv_2_wrapper
  Xinv14 x[13] vss vss vdd vdd x[14] sramgen_svt_inv_2_wrapper
  Xinv15 x[14] vss vss vdd vdd x[15] sramgen_svt_inv_2_wrapper
  Xinv16 x[15] vss vss vdd vdd x[16] sramgen_svt_inv_2_wrapper
  Xinv17 x[16] vss vss vdd vdd x[17] sramgen_svt_inv_2_wrapper
  Xinv18 x[17] vss vss vdd vdd x[18] sramgen_svt_inv_2_wrapper
  Xinv19 x[18] vss vss vdd vdd x[19] sramgen_svt_inv_2_wrapper
  Xinv20 x[19] vss vss vdd vdd x[20] sramgen_svt_inv_2_wrapper
  Xinv21 x[20] vss vss vdd vdd x[21] sramgen_svt_inv_2_wrapper
  Xinv22 x[21] vss vss vdd vdd x[22] sramgen_svt_inv_2_wrapper
  Xinv23 x[22] vss vss vdd vdd x[23] sramgen_svt_inv_2_wrapper
  Xinv24 x[23] vss vss vdd vdd x[24] sramgen_svt_inv_2_wrapper
  Xinv25 x[24] vss vss vdd vdd x[25] sramgen_svt_inv_2_wrapper
  Xinv26 x[25] vss vss vdd vdd x[26] sramgen_svt_inv_2_wrapper
  Xinv27 x[26] vss vss vdd vdd dout sramgen_svt_inv_4_wrapper

.ENDS svt_inv_chain_28

.SUBCKT inv_chain_20 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sky130_fd_sc_hs__inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd x[2] sky130_fd_sc_hs__inv_2_wrapper
  Xinv3 x[2] vss vss vdd vdd x[3] sky130_fd_sc_hs__inv_2_wrapper
  Xinv4 x[3] vss vss vdd vdd x[4] sky130_fd_sc_hs__inv_2_wrapper
  Xinv5 x[4] vss vss vdd vdd x[5] sky130_fd_sc_hs__inv_2_wrapper
  Xinv6 x[5] vss vss vdd vdd x[6] sky130_fd_sc_hs__inv_2_wrapper
  Xinv7 x[6] vss vss vdd vdd x[7] sky130_fd_sc_hs__inv_2_wrapper
  Xinv8 x[7] vss vss vdd vdd x[8] sky130_fd_sc_hs__inv_2_wrapper
  Xinv9 x[8] vss vss vdd vdd x[9] sky130_fd_sc_hs__inv_2_wrapper
  Xinv10 x[9] vss vss vdd vdd x[10] sky130_fd_sc_hs__inv_2_wrapper
  Xinv11 x[10] vss vss vdd vdd x[11] sky130_fd_sc_hs__inv_2_wrapper
  Xinv12 x[11] vss vss vdd vdd x[12] sky130_fd_sc_hs__inv_2_wrapper
  Xinv13 x[12] vss vss vdd vdd x[13] sky130_fd_sc_hs__inv_2_wrapper
  Xinv14 x[13] vss vss vdd vdd x[14] sky130_fd_sc_hs__inv_2_wrapper
  Xinv15 x[14] vss vss vdd vdd x[15] sky130_fd_sc_hs__inv_2_wrapper
  Xinv16 x[15] vss vss vdd vdd x[16] sky130_fd_sc_hs__inv_2_wrapper
  Xinv17 x[16] vss vss vdd vdd x[17] sky130_fd_sc_hs__inv_2_wrapper
  Xinv18 x[17] vss vss vdd vdd x[18] sky130_fd_sc_hs__inv_2_wrapper
  Xinv19 x[18] vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_20

.SUBCKT sky130_fd_sc_hs__nand2_8 A B VGND VNB VPB VPWR Y

  X0 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X1 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X2 Y B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X4 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X5 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X6 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X7 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X11 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X12 VPWR B Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X13 VPWR B Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X14 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X16 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X17 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X18 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X19 Y B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X20 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X21 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X22 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X23 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120


.ENDS sky130_fd_sc_hs__nand2_8

.SUBCKT sky130_fd_sc_hs__nand2_8_wrapper A B VGND VNB VPB VPWR Y

  X0 A B VGND VNB VPB VPWR Y sky130_fd_sc_hs__nand2_8

.ENDS sky130_fd_sc_hs__nand2_8_wrapper

.SUBCKT sr_latch sb rb q qb vdd vss

  Xnand_set q0b sb vss vss vdd vdd q0 sky130_fd_sc_hs__nand2_8_wrapper
  Xnand_reset q0 rb vss vss vdd vdd q0b sky130_fd_sc_hs__nand2_8_wrapper
  Xqb_inv q0 vss vss vdd vdd qb sky130_fd_sc_hs__inv_2_wrapper
  Xq_inv q0b vss vss vdd vdd q sky130_fd_sc_hs__inv_2_wrapper

.ENDS sr_latch

.SUBCKT inv_chain_2 din dout vdd vss

  Xinv0 din vss vss vdd vdd x sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_2

.SUBCKT control_logic_replica_v2 clk ce we rstb rbl saen pc_b rwl wlen wrdrven vdd vss

  Xreset_inv rstb vss vss vdd vdd reset sky130_fd_sc_hs__inv_16_wrapper
  Xclk_delay clk clkd vdd vss inv_chain_12
  Xclk_gate clkd ce vss vss vdd vdd clk_buf sky130_fd_sc_hs__and2_2_wrapper
  Xclk_pulse clk_buf clkp0 vdd vss edge_detector
  Xclk_pulse_buf clkp0 vss vss vdd vdd clkp sky130_fd_sc_hs__buf_16_wrapper
  Xclk_pulse_inv clkp vss vss vdd vdd clkp_b sky130_fd_sc_hs__inv_16_wrapper
  Xclkp_delay clkp_b clkpd vdd vss inv_chain_3
  Xclkpd_inv clkpd vss vss vdd vdd clkpd_b sky130_fd_sc_hs__inv_2_wrapper
  Xclkpd_delay clkpd_b clkpdd vdd vss inv_chain_15
  Xmux_wlen_rst rbl_b clkpdd we vss vss vdd vdd decrepstart sky130_fd_sc_hs__mux2_4_wrapper
  Xdecoder_replica decrepstart decrepend vdd vss svt_inv_chain_28
  Xdecoder_replica_delay decrepend wlen_rst_decoderd vdd vss inv_chain_20
  Xinv_we we vss vss vdd vdd we_b sky130_fd_sc_hs__inv_2_wrapper
  Xinv_rbl rbl vss vss vdd vdd rbl_b sky130_fd_sc_hs__inv_2_wrapper
  Xwlen_grst decrepstart reset vss vss vdd vdd wlen_grst_b sky130_fd_sc_hs__nor2_4_wrapper
  Xpc_set wlen_rst_decoderd reset vss vss vdd vdd pc_set_b sky130_fd_sc_hs__nor2_4_wrapper
  Xwrdrven_grst decrepend reset vss vss vdd vdd wrdrven_grst_b sky130_fd_sc_hs__nor2_4_wrapper
  Xclkp_grst clkp reset vss vss vdd vdd clkp_grst_b sky130_fd_sc_hs__nor2_4_wrapper
  Xnand_sense_en we_b decrepend vss vss vdd vdd saen_set_b sky130_fd_sc_hs__nand2_4_wrapper
  Xnand_wlendb_web rbl_b we_b vss vss vdd vdd wlend sky130_fd_sc_hs__nand2_4_wrapper
  Xand_wlen wlen_q wlend vss vss vdd vdd wlen sky130_fd_sc_hs__and2_4_wrapper
  Xrwl_buf wlen_q vss vss vdd vdd rwl sky130_fd_sc_hs__buf_16_wrapper
  Xwl_ctl clkpd_b wlen_grst_b wlen_q wlen_b vdd vss sr_latch
  Xsaen_ctl saen_set_b clkp_grst_b saen saen_b vdd vss sr_latch
  Xpc_ctl pc_set_b clkp_b pc pc_b0 vdd vss sr_latch
  Xpc_b_buf pc_b0 vss vss vdd vdd pc_b sky130_fd_sc_hs__buf_16_wrapper
  Xwrdrven_set clkpd we vss vss vdd vdd wrdrven_set_b0 sky130_fd_sc_hs__nand2_4_wrapper
  Xwrdrven_set_delay wrdrven_set_b0 wrdrven_set_b vdd vss inv_chain_2
  Xwrdrven_ctl wrdrven_set_b wrdrven_grst_b wrdrven wrdrven_b vdd vss sr_latch

.ENDS control_logic_replica_v2

.SUBCKT mos_w1250_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.250


.ENDS mos_w1250_l150_m1_nf1_id1

.SUBCKT mos_w500_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.500


.ENDS mos_w500_l150_m1_nf1_id0

.SUBCKT folded_inv vdd vss a y

  XMP0 y a vdd vdd mos_w1250_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w500_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w1250_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w500_l150_m1_nf1_id0

.ENDS folded_inv

.SUBCKT multi_finger_inv_1 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_1

.SUBCKT multi_finger_inv_2 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_2

.SUBCKT multi_finger_inv_3 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_3

.SUBCKT multi_finger_inv_4 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP19 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP20 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP21 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP22 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP23 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP24 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP25 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP26 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP27 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP28 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP29 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP30 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP31 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP32 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP33 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP34 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP35 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP36 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP37 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP38 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP39 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP40 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP41 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP42 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP43 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP44 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP45 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP46 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN7 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN8 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN9 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN10 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN11 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN12 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN13 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN14 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN15 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN16 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN17 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN18 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_4

.SUBCKT decoder_stage_1 vdd vss y y_b predecode_0_0

  Xgate_0_0_0 vdd vss predecode_0_0 x_0 folded_inv
  Xgate_1_0_0 vdd vss x_0 x_1 multi_finger_inv
  Xgate_2_0_0 vdd vss x_1 x_2 multi_finger_inv_1
  Xgate_2_0_1 vdd vss x_1 x_2 multi_finger_inv_1
  Xgate_2_0_2 vdd vss x_1 x_2 multi_finger_inv_1
  Xgate_2_0_3 vdd vss x_1 x_2 multi_finger_inv_1
  Xgate_3_0_0 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_1 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_2 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_3 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_4 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_5 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_6 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_7 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_8 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_9 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_10 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_11 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_12 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_13 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_4_0_0 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_1 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_2 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_3 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_4 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_5 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_6 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_7 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_8 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_9 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_10 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_11 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_12 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_13 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_14 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_15 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_16 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_5_0_0 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_1 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_2 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_3 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_4 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_5 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_6 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_7 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_8 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_9 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_10 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_11 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_12 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_13 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_14 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_15 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_16 vdd vss y_b y multi_finger_inv_4

.ENDS decoder_stage_1

.SUBCKT multi_finger_inv_5 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_5

.SUBCKT decoder_stage_2 vdd vss y y_b predecode_0_0

  Xgate_0_0_0 vdd vss predecode_0_0 y_b folded_inv
  Xgate_1_0_0 vdd vss y_b y multi_finger_inv_5
  Xgate_1_0_1 vdd vss y_b y multi_finger_inv_5

.ENDS decoder_stage_2

.SUBCKT multi_finger_inv_6 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_6

.SUBCKT decoder_stage_3 vdd vss y y_b predecode_0_0

  Xgate_0_0_0 vdd vss predecode_0_0 y_b folded_inv
  Xgate_1_0_0 vdd vss y_b y multi_finger_inv_6
  Xgate_1_0_1 vdd vss y_b y multi_finger_inv_6

.ENDS decoder_stage_3

.SUBCKT multi_finger_inv_7 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_7

.SUBCKT multi_finger_inv_8 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_8

.SUBCKT multi_finger_inv_9 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP19 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP20 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP21 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP22 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP23 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP24 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP25 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP26 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP27 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP28 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP29 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP30 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP31 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP32 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP33 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP34 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP35 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP36 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP37 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP38 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP39 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP40 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP41 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP42 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP43 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP44 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP45 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP46 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP47 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP48 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP49 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP50 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP51 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP52 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP53 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP54 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP55 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP56 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN7 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN8 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN9 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN10 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN11 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN12 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN13 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN14 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN15 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN16 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN17 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN18 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN19 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN20 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN21 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN22 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_9

.SUBCKT decoder_stage_4 vdd vss y y_b predecode_0_0

  Xgate_0_0_0 vdd vss predecode_0_0 x_0 folded_inv
  Xgate_1_0_0 vdd vss x_0 x_1 multi_finger_inv_7
  Xgate_1_0_1 vdd vss x_0 x_1 multi_finger_inv_7
  Xgate_2_0_0 vdd vss x_1 y_b multi_finger_inv_8
  Xgate_2_0_1 vdd vss x_1 y_b multi_finger_inv_8
  Xgate_2_0_2 vdd vss x_1 y_b multi_finger_inv_8
  Xgate_3_0_0 vdd vss y_b y multi_finger_inv_9
  Xgate_3_0_1 vdd vss y_b y multi_finger_inv_9
  Xgate_3_0_2 vdd vss y_b y multi_finger_inv_9

.ENDS decoder_stage_4

.SUBCKT sram_sp_cell_replica BL BR VSS VDD VPB VNB WL

  X0 VDD WL BR VNB sky130_fd_pr__special_nfet_pass l=0.150 nf=1 w=0.140

  X1 Q VDD VSS VNB sky130_fd_pr__special_nfet_latch l=0.150 nf=1 w=0.210

  X2 BL WL Q VNB sky130_fd_pr__special_nfet_pass l=0.150 nf=1 w=0.140

  X3 Q WL Q VPB sky130_fd_pr__special_pfet_pass l=0.025 nf=1 w=0.140

  X4 VDD WL VDD VPB sky130_fd_pr__special_pfet_pass l=0.025 nf=1 w=0.140

  X5 VDD Q VDD VPB sky130_fd_pr__special_pfet_pass l=0.150 nf=1 w=0.140

  X6 Q VDD VDD VPB sky130_fd_pr__special_pfet_pass l=0.150 nf=1 w=0.140

  X7 VSS Q VDD VNB sky130_fd_pr__special_nfet_latch l=0.150 nf=1 w=0.210


.ENDS sram_sp_cell_replica

.SUBCKT sram_sp_cell_replica_wrapper BL BR VSS VDD VPB VNB WL

  X0 BL BR VSS VDD VPB VNB WL sram_sp_cell_replica

.ENDS sram_sp_cell_replica_wrapper

.SUBCKT sram_sp_rowtapend_replica VSS VNB

  X0 VSS VSS VSS VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.420


.ENDS sram_sp_rowtapend_replica

.SUBCKT sram_sp_rowtapend_replica_wrapper VSS VNB

  X0 VSS VNB sram_sp_rowtapend_replica

.ENDS sram_sp_rowtapend_replica_wrapper

.SUBCKT replica_cell_array vdd vss rbl rbr rwl

  Xcell_0_0 rbl rbr vss vdd vdd vss rwl sram_sp_cell_replica_wrapper
  Xcell_0_1 rbl rbr vss vdd vdd vss rwl sram_sp_cell_replica_wrapper
  Xcell_1_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_1_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_2_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_2_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_3_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_3_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_4_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_4_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_5_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_5_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_6_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_6_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_7_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_7_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_8_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_8_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_9_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_9_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_10_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_10_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_11_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_11_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_12_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_12_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_13_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_13_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_14_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_14_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_15_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_15_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_16_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_16_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_17_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_17_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_18_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_18_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_19_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_19_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_20_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_20_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_21_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_21_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_22_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_22_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_23_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_23_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_24_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_24_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_25_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_25_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcolend_0_0 rbr vdd vss rbl vss vdd sram_sp_colend_wrapper
  Xcolend_1_0 rbr vdd vss rbl vss vdd sram_sp_colend_wrapper
  Xcolend_0_1 rbr vdd vss rbl vss vdd sram_sp_colend_wrapper
  Xcolend_1_1 rbr vdd vss rbl vss vdd sram_sp_colend_wrapper
  Xrowtapend_0_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_0_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_0_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_0_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xrowtapend_1_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_1_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_1_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xrowtapend_2_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_2_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_2_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xrowtapend_3_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_3_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_3_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xrowtapend_4_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_4_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_4_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xrowtapend_5_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_5_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_5_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xrowtapend_6_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_6_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_6_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper

.ENDS replica_cell_array

.SUBCKT dff_array_8 vdd vss clk rb d[0] d[1] d[2] d[3] d[4] d[5] d[6] d[7] q[0] q[1] q[2] q[3] q[4] q[5] q[6] q[7] qn[0] qn[1] qn[2] qn[3] qn[4] qn[5] qn[6] qn[7]

  Xdff_0 clk d[0] rb vss vss vdd vdd q[0] qn[0] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_1 clk d[1] rb vss vss vdd vdd q[1] qn[1] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_2 clk d[2] rb vss vss vdd vdd q[2] qn[2] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_3 clk d[3] rb vss vss vdd vdd q[3] qn[3] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_4 clk d[4] rb vss vss vdd vdd q[4] qn[4] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_5 clk d[5] rb vss vss vdd vdd q[5] qn[5] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_6 clk d[6] rb vss vss vdd vdd q[6] qn[6] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_7 clk d[7] rb vss vss vdd vdd q[7] qn[7] sky130_fd_sc_hs__dfrbp_2_wrapper

.ENDS dff_array_8

.SUBCKT mos_w2550_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.550


.ENDS mos_w2550_l150_m1_nf1_id1

.SUBCKT mos_w1030_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.030


.ENDS mos_w1030_l150_m1_nf1_id0

.SUBCKT folded_inv_3 vdd vss a y

  XMP0 y a vdd vdd mos_w2550_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w1030_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w2550_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w1030_l150_m1_nf1_id0

.ENDS folded_inv_3

.SUBCKT mos_w2640_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.640


.ENDS mos_w2640_l150_m1_nf1_id1

.SUBCKT mos_w1060_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.060


.ENDS mos_w1060_l150_m1_nf1_id0

.SUBCKT folded_inv_4 vdd vss a y

  XMP0 y a vdd vdd mos_w2640_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w1060_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w2640_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w1060_l150_m1_nf1_id0

.ENDS folded_inv_4

.SUBCKT mos_w2420_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.420


.ENDS mos_w2420_l150_m1_nf1_id1

.SUBCKT mos_w970_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.970


.ENDS mos_w970_l150_m1_nf1_id0

.SUBCKT folded_inv_5 vdd vss a y

  XMP0 y a vdd vdd mos_w2420_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w970_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w2420_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w970_l150_m1_nf1_id0

.ENDS folded_inv_5

.SUBCKT decoder_stage_7 vdd vss y y_b predecode_0_0 predecode_1_0

  Xgate_0_0_0 vdd vss predecode_0_0 predecode_1_0 x_0 nand2_1
  Xgate_1_0_0 vdd vss x_0 x_1 folded_inv_2
  Xgate_2_0_0 vdd vss x_1 x_2 folded_inv_3
  Xgate_2_0_1 vdd vss x_1 x_2 folded_inv_3
  Xgate_3_0_0 vdd vss x_2 x_3 folded_inv_4
  Xgate_3_0_1 vdd vss x_2 x_3 folded_inv_4
  Xgate_3_0_2 vdd vss x_2 x_3 folded_inv_4
  Xgate_3_0_3 vdd vss x_2 x_3 folded_inv_4
  Xgate_4_0_0 vdd vss x_3 y_b folded_inv_5
  Xgate_4_0_1 vdd vss x_3 y_b folded_inv_5
  Xgate_4_0_2 vdd vss x_3 y_b folded_inv_5
  Xgate_4_0_3 vdd vss x_3 y_b folded_inv_5
  Xgate_4_0_4 vdd vss x_3 y_b folded_inv_5
  Xgate_4_0_5 vdd vss x_3 y_b folded_inv_5
  Xgate_4_0_6 vdd vss x_3 y_b folded_inv_5
  Xgate_4_0_7 vdd vss x_3 y_b folded_inv_5
  Xgate_4_0_8 vdd vss x_3 y_b folded_inv_5
  Xgate_5_0_0 vdd vss y_b y folded_inv_5
  Xgate_5_0_1 vdd vss y_b y folded_inv_5
  Xgate_5_0_2 vdd vss y_b y folded_inv_5
  Xgate_5_0_3 vdd vss y_b y folded_inv_5
  Xgate_5_0_4 vdd vss y_b y folded_inv_5
  Xgate_5_0_5 vdd vss y_b y folded_inv_5
  Xgate_5_0_6 vdd vss y_b y folded_inv_5
  Xgate_5_0_7 vdd vss y_b y folded_inv_5
  Xgate_5_0_8 vdd vss y_b y folded_inv_5

.ENDS decoder_stage_7

.SUBCKT precharge_1 vdd bl br en_b

  Xbl_pull_up bl en_b vdd vdd mos_w5000_l150_m1_nf1_id1
  Xbr_pull_up br en_b vdd vdd mos_w5000_l150_m1_nf1_id1
  Xequalizer bl en_b br vdd mos_w3000_l150_m1_nf1_id1

.ENDS precharge_1

.SUBCKT mos_w4700_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=4.700


.ENDS mos_w4700_l150_m1_nf1_id0

.SUBCKT tgate_mux sel_b sel bl br bl_out br_out vdd vss

  XMPBL bl_out sel_b bl vdd mos_w7050_l150_m1_nf1_id1
  XMPBR br_out sel_b br vdd mos_w7050_l150_m1_nf1_id1
  XMNBL bl_out sel bl vss mos_w4700_l150_m1_nf1_id0
  XMNBR br_out sel br vss mos_w4700_l150_m1_nf1_id0

.ENDS tgate_mux

.SUBCKT mos_w5000_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=5.000


.ENDS mos_w5000_l150_m1_nf1_id0

.SUBCKT tristate_inv din en en_b din_b vdd vss

  Xmn_en din_b en nint vss mos_w5000_l150_m1_nf1_id0
  Xmn_pd nint din vss vss mos_w5000_l150_m1_nf1_id0
  Xmp_en din_b en_b pint vdd mos_w5000_l150_m1_nf1_id1
  Xmp_pu pint din vdd vdd mos_w5000_l150_m1_nf1_id1

.ENDS tristate_inv

.SUBCKT write_driver en en_b data data_b bl br vdd vss

  Xbldriver data_b en en_b bl vdd vss tristate_inv
  Xbrdriver data en en_b br vdd vss tristate_inv

.ENDS write_driver

.SUBCKT sramgen_sp_sense_amp clk inn inp outn outp VDD VSS

  XSWOP outp clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=1.000

  XSWON outn clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=1.000

  XSWMP midp clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=1.000

  XSWMN midn clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=1.000

  XPFBP outp outn VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=2.000

  XPFBN outn outp VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=2.000

  XTAIL tail clk VSS VSS sky130_fd_pr__nfet_01v8 l=0.150 nf=4 w=1.680

  XNFBP outp outn midp VSS sky130_fd_pr__nfet_01v8 l=0.150 nf=2 w=1.680

  XNFBN outn outp midn VSS sky130_fd_pr__nfet_01v8 l=0.150 nf=2 w=1.680

  XINP midn inp tail VSS sky130_fd_pr__nfet_01v8 l=0.150 nf=2 w=1.680

  XINN midp inn tail VSS sky130_fd_pr__nfet_01v8 l=0.150 nf=2 w=1.680


.ENDS sramgen_sp_sense_amp

.SUBCKT sramgen_sp_sense_amp_wrapper clk inn inp outn outp VDD VSS

  X0 clk inn inp outn outp VDD VSS sramgen_sp_sense_amp

.ENDS sramgen_sp_sense_amp_wrapper

.SUBCKT mos_w1000_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000


.ENDS mos_w1000_l150_m1_nf1_id1

.SUBCKT folded_inv_9 vdd vss a y

  XMP0 y a vdd vdd mos_w1000_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w600_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w1000_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w600_l150_m1_nf1_id0

.ENDS folded_inv_9

.SUBCKT diff_latch vdd vss din1 din2 dout1 dout2

  Xinbuf_1 vdd vss din1 rst folded_inv_9
  Xinbuf_2 vdd vss din2 set folded_inv_9
  Xoutbuf_1 vdd vss q dout2 folded_inv_9
  Xoutbuf_2 vdd vss qb dout1 folded_inv_9
  Xinvq_1 vdd vss q qb folded_inv_9
  Xinvq_2 vdd vss qb q folded_inv_9
  XMN10 q rst vss vss mos_w1000_l150_m1_nf1_id0
  XMN11 q rst vss vss mos_w1000_l150_m1_nf1_id0
  XMN20 qb set vss vss mos_w1000_l150_m1_nf1_id0
  XMN21 qb set vss vss mos_w1000_l150_m1_nf1_id0

.ENDS diff_latch

.SUBCKT column clk rstb vdd vss bl[0] bl[1] bl[2] bl[3] br[0] br[1] br[2] br[3] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we we_b din dout sense_en

  Xprecharge_0 vdd bl[0] br[0] pc_b precharge_1
  Xmux_0 sel_b[0] sel[0] bl[0] br[0] bl_out br_out vdd vss tgate_mux
  Xprecharge_1 vdd bl[1] br[1] pc_b precharge_1
  Xmux_1 sel_b[1] sel[1] bl[1] br[1] bl_out br_out vdd vss tgate_mux
  Xprecharge_2 vdd bl[2] br[2] pc_b precharge_1
  Xmux_2 sel_b[2] sel[2] bl[2] br[2] bl_out br_out vdd vss tgate_mux
  Xprecharge_3 vdd bl[3] br[3] pc_b precharge_1
  Xmux_3 sel_b[3] sel[3] bl[3] br[3] bl_out br_out vdd vss tgate_mux
  Xwrite_driver we we_b q q_b bl_out br_out vdd vss write_driver
  Xsense_amp sense_en br_out bl_out sa_outn sa_outp vdd vss sramgen_sp_sense_amp_wrapper
  Xlatch vdd vss sa_outp sa_outn dout diff_latch_outn diff_latch
  Xdff clk din rstb vss vss vdd vdd q q_b sky130_fd_sc_hs__dfrbp_2_wrapper

.ENDS column

.SUBCKT col_peripherals clk rstb vdd vss sense_en bl[0] bl[1] bl[2] bl[3] bl[4] bl[5] bl[6] bl[7] bl[8] bl[9] bl[10] bl[11] bl[12] bl[13] bl[14] bl[15] bl[16] bl[17] bl[18] bl[19] bl[20] bl[21] bl[22] bl[23] bl[24] bl[25] bl[26] bl[27] bl[28] bl[29] bl[30] bl[31] bl[32] bl[33] bl[34] bl[35] bl[36] bl[37] bl[38] bl[39] bl[40] bl[41] bl[42] bl[43] bl[44] bl[45] bl[46] bl[47] bl[48] bl[49] bl[50] bl[51] bl[52] bl[53] bl[54] bl[55] bl[56] bl[57] bl[58] bl[59] bl[60] bl[61] bl[62] bl[63] bl[64] bl[65] bl[66] bl[67] bl[68] bl[69] bl[70] bl[71] bl[72] bl[73] bl[74] bl[75] bl[76] bl[77] bl[78] bl[79] bl[80] bl[81] bl[82] bl[83] bl[84] bl[85] bl[86] bl[87] bl[88] bl[89] bl[90] bl[91] bl[92] bl[93] bl[94] bl[95] bl[96] bl[97] bl[98] bl[99] bl[100] bl[101] bl[102] bl[103] bl[104] bl[105] bl[106] bl[107] bl[108] bl[109] bl[110] bl[111] bl[112] bl[113] bl[114] bl[115] bl[116] bl[117] bl[118] bl[119] bl[120] bl[121] bl[122] bl[123] bl[124] bl[125] bl[126] bl[127] bl[128] bl[129] bl[130] bl[131] bl[132] bl[133] bl[134] bl[135] bl[136] bl[137] bl[138] bl[139] bl[140] bl[141] bl[142] bl[143] bl[144] bl[145] bl[146] bl[147] bl[148] bl[149] bl[150] bl[151] bl[152] bl[153] bl[154] bl[155] bl[156] bl[157] bl[158] bl[159] bl[160] bl[161] bl[162] bl[163] bl[164] bl[165] bl[166] bl[167] bl[168] bl[169] bl[170] bl[171] bl[172] bl[173] bl[174] bl[175] bl[176] bl[177] bl[178] bl[179] bl[180] bl[181] bl[182] bl[183] bl[184] bl[185] bl[186] bl[187] bl[188] bl[189] bl[190] bl[191] bl[192] bl[193] bl[194] bl[195] bl[196] bl[197] bl[198] bl[199] bl[200] bl[201] bl[202] bl[203] bl[204] bl[205] bl[206] bl[207] bl[208] bl[209] bl[210] bl[211] bl[212] bl[213] bl[214] bl[215] bl[216] bl[217] bl[218] bl[219] bl[220] bl[221] bl[222] bl[223] bl[224] bl[225] bl[226] bl[227] bl[228] bl[229] bl[230] bl[231] bl[232] bl[233] bl[234] bl[235] bl[236] bl[237] bl[238] bl[239] bl[240] bl[241] bl[242] bl[243] bl[244] bl[245] bl[246] bl[247] bl[248] bl[249] bl[250] bl[251] bl[252] bl[253] bl[254] bl[255] br[0] br[1] br[2] br[3] br[4] br[5] br[6] br[7] br[8] br[9] br[10] br[11] br[12] br[13] br[14] br[15] br[16] br[17] br[18] br[19] br[20] br[21] br[22] br[23] br[24] br[25] br[26] br[27] br[28] br[29] br[30] br[31] br[32] br[33] br[34] br[35] br[36] br[37] br[38] br[39] br[40] br[41] br[42] br[43] br[44] br[45] br[46] br[47] br[48] br[49] br[50] br[51] br[52] br[53] br[54] br[55] br[56] br[57] br[58] br[59] br[60] br[61] br[62] br[63] br[64] br[65] br[66] br[67] br[68] br[69] br[70] br[71] br[72] br[73] br[74] br[75] br[76] br[77] br[78] br[79] br[80] br[81] br[82] br[83] br[84] br[85] br[86] br[87] br[88] br[89] br[90] br[91] br[92] br[93] br[94] br[95] br[96] br[97] br[98] br[99] br[100] br[101] br[102] br[103] br[104] br[105] br[106] br[107] br[108] br[109] br[110] br[111] br[112] br[113] br[114] br[115] br[116] br[117] br[118] br[119] br[120] br[121] br[122] br[123] br[124] br[125] br[126] br[127] br[128] br[129] br[130] br[131] br[132] br[133] br[134] br[135] br[136] br[137] br[138] br[139] br[140] br[141] br[142] br[143] br[144] br[145] br[146] br[147] br[148] br[149] br[150] br[151] br[152] br[153] br[154] br[155] br[156] br[157] br[158] br[159] br[160] br[161] br[162] br[163] br[164] br[165] br[166] br[167] br[168] br[169] br[170] br[171] br[172] br[173] br[174] br[175] br[176] br[177] br[178] br[179] br[180] br[181] br[182] br[183] br[184] br[185] br[186] br[187] br[188] br[189] br[190] br[191] br[192] br[193] br[194] br[195] br[196] br[197] br[198] br[199] br[200] br[201] br[202] br[203] br[204] br[205] br[206] br[207] br[208] br[209] br[210] br[211] br[212] br[213] br[214] br[215] br[216] br[217] br[218] br[219] br[220] br[221] br[222] br[223] br[224] br[225] br[226] br[227] br[228] br[229] br[230] br[231] br[232] br[233] br[234] br[235] br[236] br[237] br[238] br[239] br[240] br[241] br[242] br[243] br[244] br[245] br[246] br[247] br[248] br[249] br[250] br[251] br[252] br[253] br[254] br[255] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we wmask[0] wmask[1] wmask[2] wmask[3] wmask[4] wmask[5] wmask[6] wmask[7] din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] din[8] din[9] din[10] din[11] din[12] din[13] din[14] din[15] din[16] din[17] din[18] din[19] din[20] din[21] din[22] din[23] din[24] din[25] din[26] din[27] din[28] din[29] din[30] din[31] din[32] din[33] din[34] din[35] din[36] din[37] din[38] din[39] din[40] din[41] din[42] din[43] din[44] din[45] din[46] din[47] din[48] din[49] din[50] din[51] din[52] din[53] din[54] din[55] din[56] din[57] din[58] din[59] din[60] din[61] din[62] din[63] dout[0] dout[1] dout[2] dout[3] dout[4] dout[5] dout[6] dout[7] dout[8] dout[9] dout[10] dout[11] dout[12] dout[13] dout[14] dout[15] dout[16] dout[17] dout[18] dout[19] dout[20] dout[21] dout[22] dout[23] dout[24] dout[25] dout[26] dout[27] dout[28] dout[29] dout[30] dout[31] dout[32] dout[33] dout[34] dout[35] dout[36] dout[37] dout[38] dout[39] dout[40] dout[41] dout[42] dout[43] dout[44] dout[45] dout[46] dout[47] dout[48] dout[49] dout[50] dout[51] dout[52] dout[53] dout[54] dout[55] dout[56] dout[57] dout[58] dout[59] dout[60] dout[61] dout[62] dout[63]

  Xwmask_dffs vdd vss clk rstb wmask[0] wmask[1] wmask[2] wmask[3] wmask[4] wmask[5] wmask[6] wmask[7] wmask_in[0] wmask_in[1] wmask_in[2] wmask_in[3] wmask_in[4] wmask_in[5] wmask_in[6] wmask_in[7] wmask_in_b[0] wmask_in_b[1] wmask_in_b[2] wmask_in_b[3] wmask_in_b[4] wmask_in_b[5] wmask_in_b[6] wmask_in_b[7] dff_array_8
  Xwmask_and_0 vdd vss we_i[0] we_ib[0] we wmask_in[0] decoder_stage_7
  Xwmask_and_1 vdd vss we_i[1] we_ib[1] we wmask_in[1] decoder_stage_7
  Xwmask_and_2 vdd vss we_i[2] we_ib[2] we wmask_in[2] decoder_stage_7
  Xwmask_and_3 vdd vss we_i[3] we_ib[3] we wmask_in[3] decoder_stage_7
  Xwmask_and_4 vdd vss we_i[4] we_ib[4] we wmask_in[4] decoder_stage_7
  Xwmask_and_5 vdd vss we_i[5] we_ib[5] we wmask_in[5] decoder_stage_7
  Xwmask_and_6 vdd vss we_i[6] we_ib[6] we wmask_in[6] decoder_stage_7
  Xwmask_and_7 vdd vss we_i[7] we_ib[7] we wmask_in[7] decoder_stage_7
  Xcol_group_0 clk rstb vdd vss bl[0] bl[1] bl[2] bl[3] br[0] br[1] br[2] br[3] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[0] we_ib[0] din[0] dout[0] sense_en column
  Xcol_group_1 clk rstb vdd vss bl[4] bl[5] bl[6] bl[7] br[4] br[5] br[6] br[7] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[0] we_ib[0] din[1] dout[1] sense_en column
  Xcol_group_2 clk rstb vdd vss bl[8] bl[9] bl[10] bl[11] br[8] br[9] br[10] br[11] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[0] we_ib[0] din[2] dout[2] sense_en column
  Xcol_group_3 clk rstb vdd vss bl[12] bl[13] bl[14] bl[15] br[12] br[13] br[14] br[15] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[0] we_ib[0] din[3] dout[3] sense_en column
  Xcol_group_4 clk rstb vdd vss bl[16] bl[17] bl[18] bl[19] br[16] br[17] br[18] br[19] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[0] we_ib[0] din[4] dout[4] sense_en column
  Xcol_group_5 clk rstb vdd vss bl[20] bl[21] bl[22] bl[23] br[20] br[21] br[22] br[23] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[0] we_ib[0] din[5] dout[5] sense_en column
  Xcol_group_6 clk rstb vdd vss bl[24] bl[25] bl[26] bl[27] br[24] br[25] br[26] br[27] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[0] we_ib[0] din[6] dout[6] sense_en column
  Xcol_group_7 clk rstb vdd vss bl[28] bl[29] bl[30] bl[31] br[28] br[29] br[30] br[31] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[0] we_ib[0] din[7] dout[7] sense_en column
  Xcol_group_8 clk rstb vdd vss bl[32] bl[33] bl[34] bl[35] br[32] br[33] br[34] br[35] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[1] we_ib[1] din[8] dout[8] sense_en column
  Xcol_group_9 clk rstb vdd vss bl[36] bl[37] bl[38] bl[39] br[36] br[37] br[38] br[39] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[1] we_ib[1] din[9] dout[9] sense_en column
  Xcol_group_10 clk rstb vdd vss bl[40] bl[41] bl[42] bl[43] br[40] br[41] br[42] br[43] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[1] we_ib[1] din[10] dout[10] sense_en column
  Xcol_group_11 clk rstb vdd vss bl[44] bl[45] bl[46] bl[47] br[44] br[45] br[46] br[47] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[1] we_ib[1] din[11] dout[11] sense_en column
  Xcol_group_12 clk rstb vdd vss bl[48] bl[49] bl[50] bl[51] br[48] br[49] br[50] br[51] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[1] we_ib[1] din[12] dout[12] sense_en column
  Xcol_group_13 clk rstb vdd vss bl[52] bl[53] bl[54] bl[55] br[52] br[53] br[54] br[55] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[1] we_ib[1] din[13] dout[13] sense_en column
  Xcol_group_14 clk rstb vdd vss bl[56] bl[57] bl[58] bl[59] br[56] br[57] br[58] br[59] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[1] we_ib[1] din[14] dout[14] sense_en column
  Xcol_group_15 clk rstb vdd vss bl[60] bl[61] bl[62] bl[63] br[60] br[61] br[62] br[63] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[1] we_ib[1] din[15] dout[15] sense_en column
  Xcol_group_16 clk rstb vdd vss bl[64] bl[65] bl[66] bl[67] br[64] br[65] br[66] br[67] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[2] we_ib[2] din[16] dout[16] sense_en column
  Xcol_group_17 clk rstb vdd vss bl[68] bl[69] bl[70] bl[71] br[68] br[69] br[70] br[71] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[2] we_ib[2] din[17] dout[17] sense_en column
  Xcol_group_18 clk rstb vdd vss bl[72] bl[73] bl[74] bl[75] br[72] br[73] br[74] br[75] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[2] we_ib[2] din[18] dout[18] sense_en column
  Xcol_group_19 clk rstb vdd vss bl[76] bl[77] bl[78] bl[79] br[76] br[77] br[78] br[79] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[2] we_ib[2] din[19] dout[19] sense_en column
  Xcol_group_20 clk rstb vdd vss bl[80] bl[81] bl[82] bl[83] br[80] br[81] br[82] br[83] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[2] we_ib[2] din[20] dout[20] sense_en column
  Xcol_group_21 clk rstb vdd vss bl[84] bl[85] bl[86] bl[87] br[84] br[85] br[86] br[87] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[2] we_ib[2] din[21] dout[21] sense_en column
  Xcol_group_22 clk rstb vdd vss bl[88] bl[89] bl[90] bl[91] br[88] br[89] br[90] br[91] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[2] we_ib[2] din[22] dout[22] sense_en column
  Xcol_group_23 clk rstb vdd vss bl[92] bl[93] bl[94] bl[95] br[92] br[93] br[94] br[95] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[2] we_ib[2] din[23] dout[23] sense_en column
  Xcol_group_24 clk rstb vdd vss bl[96] bl[97] bl[98] bl[99] br[96] br[97] br[98] br[99] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[3] we_ib[3] din[24] dout[24] sense_en column
  Xcol_group_25 clk rstb vdd vss bl[100] bl[101] bl[102] bl[103] br[100] br[101] br[102] br[103] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[3] we_ib[3] din[25] dout[25] sense_en column
  Xcol_group_26 clk rstb vdd vss bl[104] bl[105] bl[106] bl[107] br[104] br[105] br[106] br[107] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[3] we_ib[3] din[26] dout[26] sense_en column
  Xcol_group_27 clk rstb vdd vss bl[108] bl[109] bl[110] bl[111] br[108] br[109] br[110] br[111] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[3] we_ib[3] din[27] dout[27] sense_en column
  Xcol_group_28 clk rstb vdd vss bl[112] bl[113] bl[114] bl[115] br[112] br[113] br[114] br[115] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[3] we_ib[3] din[28] dout[28] sense_en column
  Xcol_group_29 clk rstb vdd vss bl[116] bl[117] bl[118] bl[119] br[116] br[117] br[118] br[119] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[3] we_ib[3] din[29] dout[29] sense_en column
  Xcol_group_30 clk rstb vdd vss bl[120] bl[121] bl[122] bl[123] br[120] br[121] br[122] br[123] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[3] we_ib[3] din[30] dout[30] sense_en column
  Xcol_group_31 clk rstb vdd vss bl[124] bl[125] bl[126] bl[127] br[124] br[125] br[126] br[127] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[3] we_ib[3] din[31] dout[31] sense_en column
  Xcol_group_32 clk rstb vdd vss bl[128] bl[129] bl[130] bl[131] br[128] br[129] br[130] br[131] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[4] we_ib[4] din[32] dout[32] sense_en column
  Xcol_group_33 clk rstb vdd vss bl[132] bl[133] bl[134] bl[135] br[132] br[133] br[134] br[135] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[4] we_ib[4] din[33] dout[33] sense_en column
  Xcol_group_34 clk rstb vdd vss bl[136] bl[137] bl[138] bl[139] br[136] br[137] br[138] br[139] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[4] we_ib[4] din[34] dout[34] sense_en column
  Xcol_group_35 clk rstb vdd vss bl[140] bl[141] bl[142] bl[143] br[140] br[141] br[142] br[143] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[4] we_ib[4] din[35] dout[35] sense_en column
  Xcol_group_36 clk rstb vdd vss bl[144] bl[145] bl[146] bl[147] br[144] br[145] br[146] br[147] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[4] we_ib[4] din[36] dout[36] sense_en column
  Xcol_group_37 clk rstb vdd vss bl[148] bl[149] bl[150] bl[151] br[148] br[149] br[150] br[151] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[4] we_ib[4] din[37] dout[37] sense_en column
  Xcol_group_38 clk rstb vdd vss bl[152] bl[153] bl[154] bl[155] br[152] br[153] br[154] br[155] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[4] we_ib[4] din[38] dout[38] sense_en column
  Xcol_group_39 clk rstb vdd vss bl[156] bl[157] bl[158] bl[159] br[156] br[157] br[158] br[159] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[4] we_ib[4] din[39] dout[39] sense_en column
  Xcol_group_40 clk rstb vdd vss bl[160] bl[161] bl[162] bl[163] br[160] br[161] br[162] br[163] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[5] we_ib[5] din[40] dout[40] sense_en column
  Xcol_group_41 clk rstb vdd vss bl[164] bl[165] bl[166] bl[167] br[164] br[165] br[166] br[167] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[5] we_ib[5] din[41] dout[41] sense_en column
  Xcol_group_42 clk rstb vdd vss bl[168] bl[169] bl[170] bl[171] br[168] br[169] br[170] br[171] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[5] we_ib[5] din[42] dout[42] sense_en column
  Xcol_group_43 clk rstb vdd vss bl[172] bl[173] bl[174] bl[175] br[172] br[173] br[174] br[175] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[5] we_ib[5] din[43] dout[43] sense_en column
  Xcol_group_44 clk rstb vdd vss bl[176] bl[177] bl[178] bl[179] br[176] br[177] br[178] br[179] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[5] we_ib[5] din[44] dout[44] sense_en column
  Xcol_group_45 clk rstb vdd vss bl[180] bl[181] bl[182] bl[183] br[180] br[181] br[182] br[183] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[5] we_ib[5] din[45] dout[45] sense_en column
  Xcol_group_46 clk rstb vdd vss bl[184] bl[185] bl[186] bl[187] br[184] br[185] br[186] br[187] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[5] we_ib[5] din[46] dout[46] sense_en column
  Xcol_group_47 clk rstb vdd vss bl[188] bl[189] bl[190] bl[191] br[188] br[189] br[190] br[191] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[5] we_ib[5] din[47] dout[47] sense_en column
  Xcol_group_48 clk rstb vdd vss bl[192] bl[193] bl[194] bl[195] br[192] br[193] br[194] br[195] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[6] we_ib[6] din[48] dout[48] sense_en column
  Xcol_group_49 clk rstb vdd vss bl[196] bl[197] bl[198] bl[199] br[196] br[197] br[198] br[199] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[6] we_ib[6] din[49] dout[49] sense_en column
  Xcol_group_50 clk rstb vdd vss bl[200] bl[201] bl[202] bl[203] br[200] br[201] br[202] br[203] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[6] we_ib[6] din[50] dout[50] sense_en column
  Xcol_group_51 clk rstb vdd vss bl[204] bl[205] bl[206] bl[207] br[204] br[205] br[206] br[207] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[6] we_ib[6] din[51] dout[51] sense_en column
  Xcol_group_52 clk rstb vdd vss bl[208] bl[209] bl[210] bl[211] br[208] br[209] br[210] br[211] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[6] we_ib[6] din[52] dout[52] sense_en column
  Xcol_group_53 clk rstb vdd vss bl[212] bl[213] bl[214] bl[215] br[212] br[213] br[214] br[215] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[6] we_ib[6] din[53] dout[53] sense_en column
  Xcol_group_54 clk rstb vdd vss bl[216] bl[217] bl[218] bl[219] br[216] br[217] br[218] br[219] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[6] we_ib[6] din[54] dout[54] sense_en column
  Xcol_group_55 clk rstb vdd vss bl[220] bl[221] bl[222] bl[223] br[220] br[221] br[222] br[223] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[6] we_ib[6] din[55] dout[55] sense_en column
  Xcol_group_56 clk rstb vdd vss bl[224] bl[225] bl[226] bl[227] br[224] br[225] br[226] br[227] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[7] we_ib[7] din[56] dout[56] sense_en column
  Xcol_group_57 clk rstb vdd vss bl[228] bl[229] bl[230] bl[231] br[228] br[229] br[230] br[231] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[7] we_ib[7] din[57] dout[57] sense_en column
  Xcol_group_58 clk rstb vdd vss bl[232] bl[233] bl[234] bl[235] br[232] br[233] br[234] br[235] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[7] we_ib[7] din[58] dout[58] sense_en column
  Xcol_group_59 clk rstb vdd vss bl[236] bl[237] bl[238] bl[239] br[236] br[237] br[238] br[239] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[7] we_ib[7] din[59] dout[59] sense_en column
  Xcol_group_60 clk rstb vdd vss bl[240] bl[241] bl[242] bl[243] br[240] br[241] br[242] br[243] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[7] we_ib[7] din[60] dout[60] sense_en column
  Xcol_group_61 clk rstb vdd vss bl[244] bl[245] bl[246] bl[247] br[244] br[245] br[246] br[247] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[7] we_ib[7] din[61] dout[61] sense_en column
  Xcol_group_62 clk rstb vdd vss bl[248] bl[249] bl[250] bl[251] br[248] br[249] br[250] br[251] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[7] we_ib[7] din[62] dout[62] sense_en column
  Xcol_group_63 clk rstb vdd vss bl[252] bl[253] bl[254] bl[255] br[252] br[253] br[254] br[255] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[7] we_ib[7] din[63] dout[63] sense_en column

.ENDS col_peripherals

.SUBCKT mos_w850_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.850


.ENDS mos_w850_l150_m1_nf1_id1

.SUBCKT mos_w500_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.500


.ENDS mos_w500_l150_m1_nf1_id1

.SUBCKT precharge vdd bl br en_b

  Xbl_pull_up bl en_b vdd vdd mos_w850_l150_m1_nf1_id1
  Xbr_pull_up br en_b vdd vdd mos_w850_l150_m1_nf1_id1
  Xequalizer bl en_b br vdd mos_w500_l150_m1_nf1_id1

.ENDS precharge

.SUBCKT mos_w800_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.800


.ENDS mos_w800_l150_m1_nf1_id0

.SUBCKT mos_w1600_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.600


.ENDS mos_w1600_l150_m1_nf1_id0

.SUBCKT mos_w2250_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.250


.ENDS mos_w2250_l150_m1_nf1_id1

.SUBCKT column_mos vdd vss bl

  Xgate_nmos vss bl vss vss mos_w800_l150_m1_nf1_id0
  Xdrain_nmos bl vss vss vss mos_w1600_l150_m1_nf1_id0
  Xdrain_pmos bl vdd vdd vdd mos_w2250_l150_m1_nf1_id1

.ENDS column_mos

.SUBCKT column_mos_1 vdd vss bl

  Xdrain_nmos bl vss vss vss mos_w1600_l150_m1_nf1_id0
  Xdrain_pmos bl vdd vdd vdd mos_w2250_l150_m1_nf1_id1

.ENDS column_mos_1

.SUBCKT replica_column_mos vdd vss bl

  Xunit0 vdd vss bl column_mos
  Xunit1 vdd vss bl column_mos_1
  Xunit2 vdd vss bl column_mos_1

.ENDS replica_column_mos

.SUBCKT sram22_inner vdd vss clk we ce rstb addr[0] addr[1] addr[2] addr[3] addr[4] addr[5] addr[6] addr[7] addr[8] wmask[0] wmask[1] wmask[2] wmask[3] wmask[4] wmask[5] wmask[6] wmask[7] din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] din[8] din[9] din[10] din[11] din[12] din[13] din[14] din[15] din[16] din[17] din[18] din[19] din[20] din[21] din[22] din[23] din[24] din[25] din[26] din[27] din[28] din[29] din[30] din[31] din[32] din[33] din[34] din[35] din[36] din[37] din[38] din[39] din[40] din[41] din[42] din[43] din[44] din[45] din[46] din[47] din[48] din[49] din[50] din[51] din[52] din[53] din[54] din[55] din[56] din[57] din[58] din[59] din[60] din[61] din[62] din[63] dout[0] dout[1] dout[2] dout[3] dout[4] dout[5] dout[6] dout[7] dout[8] dout[9] dout[10] dout[11] dout[12] dout[13] dout[14] dout[15] dout[16] dout[17] dout[18] dout[19] dout[20] dout[21] dout[22] dout[23] dout[24] dout[25] dout[26] dout[27] dout[28] dout[29] dout[30] dout[31] dout[32] dout[33] dout[34] dout[35] dout[36] dout[37] dout[38] dout[39] dout[40] dout[41] dout[42] dout[43] dout[44] dout[45] dout[46] dout[47] dout[48] dout[49] dout[50] dout[51] dout[52] dout[53] dout[54] dout[55] dout[56] dout[57] dout[58] dout[59] dout[60] dout[61] dout[62] dout[63]

  Xaddr_gate vdd vss addr_gated[0] addr_gated[1] addr_gated[2] addr_gated[3] addr_gated[4] addr_gated[5] addr_gated[6] addr_b_gated[0] addr_b_gated[1] addr_b_gated[2] addr_b_gated[3] addr_b_gated[4] addr_b_gated[5] addr_b_gated[6] addr_gate_y_b_noconn[0] addr_gate_y_b_noconn[1] addr_gate_y_b_noconn[2] addr_gate_y_b_noconn[3] addr_gate_y_b_noconn[4] addr_gate_y_b_noconn[5] addr_gate_y_b_noconn[6] addr_gate_y_b_noconn[7] addr_gate_y_b_noconn[8] addr_gate_y_b_noconn[9] addr_gate_y_b_noconn[10] addr_gate_y_b_noconn[11] addr_gate_y_b_noconn[12] addr_gate_y_b_noconn[13] wl_en addr_in[2] addr_in[3] addr_in[4] addr_in[5] addr_in[6] addr_in[7] addr_in[8] addr_in_b[2] addr_in_b[3] addr_in_b[4] addr_in_b[5] addr_in_b[6] addr_in_b[7] addr_in_b[8] decoder_stage
  Xdecoder vdd vss wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] wl_b[0] wl_b[1] wl_b[2] wl_b[3] wl_b[4] wl_b[5] wl_b[6] wl_b[7] wl_b[8] wl_b[9] wl_b[10] wl_b[11] wl_b[12] wl_b[13] wl_b[14] wl_b[15] wl_b[16] wl_b[17] wl_b[18] wl_b[19] wl_b[20] wl_b[21] wl_b[22] wl_b[23] wl_b[24] wl_b[25] wl_b[26] wl_b[27] wl_b[28] wl_b[29] wl_b[30] wl_b[31] wl_b[32] wl_b[33] wl_b[34] wl_b[35] wl_b[36] wl_b[37] wl_b[38] wl_b[39] wl_b[40] wl_b[41] wl_b[42] wl_b[43] wl_b[44] wl_b[45] wl_b[46] wl_b[47] wl_b[48] wl_b[49] wl_b[50] wl_b[51] wl_b[52] wl_b[53] wl_b[54] wl_b[55] wl_b[56] wl_b[57] wl_b[58] wl_b[59] wl_b[60] wl_b[61] wl_b[62] wl_b[63] wl_b[64] wl_b[65] wl_b[66] wl_b[67] wl_b[68] wl_b[69] wl_b[70] wl_b[71] wl_b[72] wl_b[73] wl_b[74] wl_b[75] wl_b[76] wl_b[77] wl_b[78] wl_b[79] wl_b[80] wl_b[81] wl_b[82] wl_b[83] wl_b[84] wl_b[85] wl_b[86] wl_b[87] wl_b[88] wl_b[89] wl_b[90] wl_b[91] wl_b[92] wl_b[93] wl_b[94] wl_b[95] wl_b[96] wl_b[97] wl_b[98] wl_b[99] wl_b[100] wl_b[101] wl_b[102] wl_b[103] wl_b[104] wl_b[105] wl_b[106] wl_b[107] wl_b[108] wl_b[109] wl_b[110] wl_b[111] wl_b[112] wl_b[113] wl_b[114] wl_b[115] wl_b[116] wl_b[117] wl_b[118] wl_b[119] wl_b[120] wl_b[121] wl_b[122] wl_b[123] wl_b[124] wl_b[125] wl_b[126] wl_b[127] addr_b_gated[0] addr_gated[0] addr_b_gated[1] addr_gated[1] addr_b_gated[2] addr_gated[2] addr_b_gated[3] addr_gated[3] addr_b_gated[4] addr_gated[4] addr_b_gated[5] addr_gated[5] addr_b_gated[6] addr_gated[6] decoder
  Xcolumn_decoder vdd vss col_sel[0] col_sel[1] col_sel[2] col_sel[3] col_sel_b[0] col_sel_b[1] col_sel_b[2] col_sel_b[3] addr_in_b[0] addr_in[0] addr_in_b[1] addr_in[1] decoder_1
  Xcontrol_logic clk ce_in we_in rstb rbl sense_en0 pc_b0 rwl wl_en0 write_driver_en0 vdd vss control_logic_replica_v2
  Xpc_b_buffer vdd vss pc_b pc pc_b0 decoder_stage_1
  Xwlen_buffer vdd vss wl_en wl_en_b wl_en0 decoder_stage_2
  Xwrite_driver_en_buffer vdd vss write_driver_en write_driver_en_b write_driver_en0 decoder_stage_3
  Xsense_en_buffer vdd vss sense_en sense_en_b sense_en0 decoder_stage_4
  Xaddr_we_ce_dffs vdd vss clk rstb addr[0] addr[1] addr[2] addr[3] addr[4] addr[5] addr[6] addr[7] addr[8] we ce addr_in[0] addr_in[1] addr_in[2] addr_in[3] addr_in[4] addr_in[5] addr_in[6] addr_in[7] addr_in[8] we_in ce_in addr_in_b[0] addr_in_b[1] addr_in_b[2] addr_in_b[3] addr_in_b[4] addr_in_b[5] addr_in_b[6] addr_in_b[7] addr_in_b[8] we_in_b ce_in_b dff_array_11
  Xbitcell_array vdd vss vdd vdd bl[0] bl[1] bl[2] bl[3] bl[4] bl[5] bl[6] bl[7] bl[8] bl[9] bl[10] bl[11] bl[12] bl[13] bl[14] bl[15] bl[16] bl[17] bl[18] bl[19] bl[20] bl[21] bl[22] bl[23] bl[24] bl[25] bl[26] bl[27] bl[28] bl[29] bl[30] bl[31] bl[32] bl[33] bl[34] bl[35] bl[36] bl[37] bl[38] bl[39] bl[40] bl[41] bl[42] bl[43] bl[44] bl[45] bl[46] bl[47] bl[48] bl[49] bl[50] bl[51] bl[52] bl[53] bl[54] bl[55] bl[56] bl[57] bl[58] bl[59] bl[60] bl[61] bl[62] bl[63] bl[64] bl[65] bl[66] bl[67] bl[68] bl[69] bl[70] bl[71] bl[72] bl[73] bl[74] bl[75] bl[76] bl[77] bl[78] bl[79] bl[80] bl[81] bl[82] bl[83] bl[84] bl[85] bl[86] bl[87] bl[88] bl[89] bl[90] bl[91] bl[92] bl[93] bl[94] bl[95] bl[96] bl[97] bl[98] bl[99] bl[100] bl[101] bl[102] bl[103] bl[104] bl[105] bl[106] bl[107] bl[108] bl[109] bl[110] bl[111] bl[112] bl[113] bl[114] bl[115] bl[116] bl[117] bl[118] bl[119] bl[120] bl[121] bl[122] bl[123] bl[124] bl[125] bl[126] bl[127] bl[128] bl[129] bl[130] bl[131] bl[132] bl[133] bl[134] bl[135] bl[136] bl[137] bl[138] bl[139] bl[140] bl[141] bl[142] bl[143] bl[144] bl[145] bl[146] bl[147] bl[148] bl[149] bl[150] bl[151] bl[152] bl[153] bl[154] bl[155] bl[156] bl[157] bl[158] bl[159] bl[160] bl[161] bl[162] bl[163] bl[164] bl[165] bl[166] bl[167] bl[168] bl[169] bl[170] bl[171] bl[172] bl[173] bl[174] bl[175] bl[176] bl[177] bl[178] bl[179] bl[180] bl[181] bl[182] bl[183] bl[184] bl[185] bl[186] bl[187] bl[188] bl[189] bl[190] bl[191] bl[192] bl[193] bl[194] bl[195] bl[196] bl[197] bl[198] bl[199] bl[200] bl[201] bl[202] bl[203] bl[204] bl[205] bl[206] bl[207] bl[208] bl[209] bl[210] bl[211] bl[212] bl[213] bl[214] bl[215] bl[216] bl[217] bl[218] bl[219] bl[220] bl[221] bl[222] bl[223] bl[224] bl[225] bl[226] bl[227] bl[228] bl[229] bl[230] bl[231] bl[232] bl[233] bl[234] bl[235] bl[236] bl[237] bl[238] bl[239] bl[240] bl[241] bl[242] bl[243] bl[244] bl[245] bl[246] bl[247] bl[248] bl[249] bl[250] bl[251] bl[252] bl[253] bl[254] bl[255] br[0] br[1] br[2] br[3] br[4] br[5] br[6] br[7] br[8] br[9] br[10] br[11] br[12] br[13] br[14] br[15] br[16] br[17] br[18] br[19] br[20] br[21] br[22] br[23] br[24] br[25] br[26] br[27] br[28] br[29] br[30] br[31] br[32] br[33] br[34] br[35] br[36] br[37] br[38] br[39] br[40] br[41] br[42] br[43] br[44] br[45] br[46] br[47] br[48] br[49] br[50] br[51] br[52] br[53] br[54] br[55] br[56] br[57] br[58] br[59] br[60] br[61] br[62] br[63] br[64] br[65] br[66] br[67] br[68] br[69] br[70] br[71] br[72] br[73] br[74] br[75] br[76] br[77] br[78] br[79] br[80] br[81] br[82] br[83] br[84] br[85] br[86] br[87] br[88] br[89] br[90] br[91] br[92] br[93] br[94] br[95] br[96] br[97] br[98] br[99] br[100] br[101] br[102] br[103] br[104] br[105] br[106] br[107] br[108] br[109] br[110] br[111] br[112] br[113] br[114] br[115] br[116] br[117] br[118] br[119] br[120] br[121] br[122] br[123] br[124] br[125] br[126] br[127] br[128] br[129] br[130] br[131] br[132] br[133] br[134] br[135] br[136] br[137] br[138] br[139] br[140] br[141] br[142] br[143] br[144] br[145] br[146] br[147] br[148] br[149] br[150] br[151] br[152] br[153] br[154] br[155] br[156] br[157] br[158] br[159] br[160] br[161] br[162] br[163] br[164] br[165] br[166] br[167] br[168] br[169] br[170] br[171] br[172] br[173] br[174] br[175] br[176] br[177] br[178] br[179] br[180] br[181] br[182] br[183] br[184] br[185] br[186] br[187] br[188] br[189] br[190] br[191] br[192] br[193] br[194] br[195] br[196] br[197] br[198] br[199] br[200] br[201] br[202] br[203] br[204] br[205] br[206] br[207] br[208] br[209] br[210] br[211] br[212] br[213] br[214] br[215] br[216] br[217] br[218] br[219] br[220] br[221] br[222] br[223] br[224] br[225] br[226] br[227] br[228] br[229] br[230] br[231] br[232] br[233] br[234] br[235] br[236] br[237] br[238] br[239] br[240] br[241] br[242] br[243] br[244] br[245] br[246] br[247] br[248] br[249] br[250] br[251] br[252] br[253] br[254] br[255] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] sp_cell_array
  Xreplica_bitcell_array vdd vss rbl rbr rwl replica_cell_array
  Xcol_circuitry clk rstb vdd vss sense_en bl[0] bl[1] bl[2] bl[3] bl[4] bl[5] bl[6] bl[7] bl[8] bl[9] bl[10] bl[11] bl[12] bl[13] bl[14] bl[15] bl[16] bl[17] bl[18] bl[19] bl[20] bl[21] bl[22] bl[23] bl[24] bl[25] bl[26] bl[27] bl[28] bl[29] bl[30] bl[31] bl[32] bl[33] bl[34] bl[35] bl[36] bl[37] bl[38] bl[39] bl[40] bl[41] bl[42] bl[43] bl[44] bl[45] bl[46] bl[47] bl[48] bl[49] bl[50] bl[51] bl[52] bl[53] bl[54] bl[55] bl[56] bl[57] bl[58] bl[59] bl[60] bl[61] bl[62] bl[63] bl[64] bl[65] bl[66] bl[67] bl[68] bl[69] bl[70] bl[71] bl[72] bl[73] bl[74] bl[75] bl[76] bl[77] bl[78] bl[79] bl[80] bl[81] bl[82] bl[83] bl[84] bl[85] bl[86] bl[87] bl[88] bl[89] bl[90] bl[91] bl[92] bl[93] bl[94] bl[95] bl[96] bl[97] bl[98] bl[99] bl[100] bl[101] bl[102] bl[103] bl[104] bl[105] bl[106] bl[107] bl[108] bl[109] bl[110] bl[111] bl[112] bl[113] bl[114] bl[115] bl[116] bl[117] bl[118] bl[119] bl[120] bl[121] bl[122] bl[123] bl[124] bl[125] bl[126] bl[127] bl[128] bl[129] bl[130] bl[131] bl[132] bl[133] bl[134] bl[135] bl[136] bl[137] bl[138] bl[139] bl[140] bl[141] bl[142] bl[143] bl[144] bl[145] bl[146] bl[147] bl[148] bl[149] bl[150] bl[151] bl[152] bl[153] bl[154] bl[155] bl[156] bl[157] bl[158] bl[159] bl[160] bl[161] bl[162] bl[163] bl[164] bl[165] bl[166] bl[167] bl[168] bl[169] bl[170] bl[171] bl[172] bl[173] bl[174] bl[175] bl[176] bl[177] bl[178] bl[179] bl[180] bl[181] bl[182] bl[183] bl[184] bl[185] bl[186] bl[187] bl[188] bl[189] bl[190] bl[191] bl[192] bl[193] bl[194] bl[195] bl[196] bl[197] bl[198] bl[199] bl[200] bl[201] bl[202] bl[203] bl[204] bl[205] bl[206] bl[207] bl[208] bl[209] bl[210] bl[211] bl[212] bl[213] bl[214] bl[215] bl[216] bl[217] bl[218] bl[219] bl[220] bl[221] bl[222] bl[223] bl[224] bl[225] bl[226] bl[227] bl[228] bl[229] bl[230] bl[231] bl[232] bl[233] bl[234] bl[235] bl[236] bl[237] bl[238] bl[239] bl[240] bl[241] bl[242] bl[243] bl[244] bl[245] bl[246] bl[247] bl[248] bl[249] bl[250] bl[251] bl[252] bl[253] bl[254] bl[255] br[0] br[1] br[2] br[3] br[4] br[5] br[6] br[7] br[8] br[9] br[10] br[11] br[12] br[13] br[14] br[15] br[16] br[17] br[18] br[19] br[20] br[21] br[22] br[23] br[24] br[25] br[26] br[27] br[28] br[29] br[30] br[31] br[32] br[33] br[34] br[35] br[36] br[37] br[38] br[39] br[40] br[41] br[42] br[43] br[44] br[45] br[46] br[47] br[48] br[49] br[50] br[51] br[52] br[53] br[54] br[55] br[56] br[57] br[58] br[59] br[60] br[61] br[62] br[63] br[64] br[65] br[66] br[67] br[68] br[69] br[70] br[71] br[72] br[73] br[74] br[75] br[76] br[77] br[78] br[79] br[80] br[81] br[82] br[83] br[84] br[85] br[86] br[87] br[88] br[89] br[90] br[91] br[92] br[93] br[94] br[95] br[96] br[97] br[98] br[99] br[100] br[101] br[102] br[103] br[104] br[105] br[106] br[107] br[108] br[109] br[110] br[111] br[112] br[113] br[114] br[115] br[116] br[117] br[118] br[119] br[120] br[121] br[122] br[123] br[124] br[125] br[126] br[127] br[128] br[129] br[130] br[131] br[132] br[133] br[134] br[135] br[136] br[137] br[138] br[139] br[140] br[141] br[142] br[143] br[144] br[145] br[146] br[147] br[148] br[149] br[150] br[151] br[152] br[153] br[154] br[155] br[156] br[157] br[158] br[159] br[160] br[161] br[162] br[163] br[164] br[165] br[166] br[167] br[168] br[169] br[170] br[171] br[172] br[173] br[174] br[175] br[176] br[177] br[178] br[179] br[180] br[181] br[182] br[183] br[184] br[185] br[186] br[187] br[188] br[189] br[190] br[191] br[192] br[193] br[194] br[195] br[196] br[197] br[198] br[199] br[200] br[201] br[202] br[203] br[204] br[205] br[206] br[207] br[208] br[209] br[210] br[211] br[212] br[213] br[214] br[215] br[216] br[217] br[218] br[219] br[220] br[221] br[222] br[223] br[224] br[225] br[226] br[227] br[228] br[229] br[230] br[231] br[232] br[233] br[234] br[235] br[236] br[237] br[238] br[239] br[240] br[241] br[242] br[243] br[244] br[245] br[246] br[247] br[248] br[249] br[250] br[251] br[252] br[253] br[254] br[255] pc_b col_sel[0] col_sel[1] col_sel[2] col_sel[3] col_sel_b[0] col_sel_b[1] col_sel_b[2] col_sel_b[3] write_driver_en wmask[0] wmask[1] wmask[2] wmask[3] wmask[4] wmask[5] wmask[6] wmask[7] din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] din[8] din[9] din[10] din[11] din[12] din[13] din[14] din[15] din[16] din[17] din[18] din[19] din[20] din[21] din[22] din[23] din[24] din[25] din[26] din[27] din[28] din[29] din[30] din[31] din[32] din[33] din[34] din[35] din[36] din[37] din[38] din[39] din[40] din[41] din[42] din[43] din[44] din[45] din[46] din[47] din[48] din[49] din[50] din[51] din[52] din[53] din[54] din[55] din[56] din[57] din[58] din[59] din[60] din[61] din[62] din[63] dout[0] dout[1] dout[2] dout[3] dout[4] dout[5] dout[6] dout[7] dout[8] dout[9] dout[10] dout[11] dout[12] dout[13] dout[14] dout[15] dout[16] dout[17] dout[18] dout[19] dout[20] dout[21] dout[22] dout[23] dout[24] dout[25] dout[26] dout[27] dout[28] dout[29] dout[30] dout[31] dout[32] dout[33] dout[34] dout[35] dout[36] dout[37] dout[38] dout[39] dout[40] dout[41] dout[42] dout[43] dout[44] dout[45] dout[46] dout[47] dout[48] dout[49] dout[50] dout[51] dout[52] dout[53] dout[54] dout[55] dout[56] dout[57] dout[58] dout[59] dout[60] dout[61] dout[62] dout[63] col_peripherals
  Xreplica_precharge_0 vdd rbl rbr pc_b0 precharge
  Xreplica_precharge_1 vdd rbl rbr pc_b0 precharge
  Xreplica_mos vdd vss rbl replica_column_mos

.ENDS sram22_inner

.SUBCKT sram22_512x64m4w8 vdd vss clk we ce rstb addr[0] addr[1] addr[2] addr[3] addr[4] addr[5] addr[6] addr[7] addr[8] wmask[0] wmask[1] wmask[2] wmask[3] wmask[4] wmask[5] wmask[6] wmask[7] din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] din[8] din[9] din[10] din[11] din[12] din[13] din[14] din[15] din[16] din[17] din[18] din[19] din[20] din[21] din[22] din[23] din[24] din[25] din[26] din[27] din[28] din[29] din[30] din[31] din[32] din[33] din[34] din[35] din[36] din[37] din[38] din[39] din[40] din[41] din[42] din[43] din[44] din[45] din[46] din[47] din[48] din[49] din[50] din[51] din[52] din[53] din[54] din[55] din[56] din[57] din[58] din[59] din[60] din[61] din[62] din[63] dout[0] dout[1] dout[2] dout[3] dout[4] dout[5] dout[6] dout[7] dout[8] dout[9] dout[10] dout[11] dout[12] dout[13] dout[14] dout[15] dout[16] dout[17] dout[18] dout[19] dout[20] dout[21] dout[22] dout[23] dout[24] dout[25] dout[26] dout[27] dout[28] dout[29] dout[30] dout[31] dout[32] dout[33] dout[34] dout[35] dout[36] dout[37] dout[38] dout[39] dout[40] dout[41] dout[42] dout[43] dout[44] dout[45] dout[46] dout[47] dout[48] dout[49] dout[50] dout[51] dout[52] dout[53] dout[54] dout[55] dout[56] dout[57] dout[58] dout[59] dout[60] dout[61] dout[62] dout[63]

  X0 vdd vss clk we ce rstb addr[0] addr[1] addr[2] addr[3] addr[4] addr[5] addr[6] addr[7] addr[8] wmask[0] wmask[1] wmask[2] wmask[3] wmask[4] wmask[5] wmask[6] wmask[7] din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] din[8] din[9] din[10] din[11] din[12] din[13] din[14] din[15] din[16] din[17] din[18] din[19] din[20] din[21] din[22] din[23] din[24] din[25] din[26] din[27] din[28] din[29] din[30] din[31] din[32] din[33] din[34] din[35] din[36] din[37] din[38] din[39] din[40] din[41] din[42] din[43] din[44] din[45] din[46] din[47] din[48] din[49] din[50] din[51] din[52] din[53] din[54] din[55] din[56] din[57] din[58] din[59] din[60] din[61] din[62] din[63] dout[0] dout[1] dout[2] dout[3] dout[4] dout[5] dout[6] dout[7] dout[8] dout[9] dout[10] dout[11] dout[12] dout[13] dout[14] dout[15] dout[16] dout[17] dout[18] dout[19] dout[20] dout[21] dout[22] dout[23] dout[24] dout[25] dout[26] dout[27] dout[28] dout[29] dout[30] dout[31] dout[32] dout[33] dout[34] dout[35] dout[36] dout[37] dout[38] dout[39] dout[40] dout[41] dout[42] dout[43] dout[44] dout[45] dout[46] dout[47] dout[48] dout[49] dout[50] dout[51] dout[52] dout[53] dout[54] dout[55] dout[56] dout[57] dout[58] dout[59] dout[60] dout[61] dout[62] dout[63] sram22_inner

.ENDS sram22_512x64m4w8

