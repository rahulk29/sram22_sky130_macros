VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram22_256x32m4w8
  CLASS BLOCK ;
  ORIGIN 76.825 224.365 ;
  FOREIGN sram22_256x32m4w8 -76.825 -224.365 ;
  SIZE 292.37 BY 358.29 ;
  SYMMETRY X Y R90 ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 206.555 132.52 206.885 133.65 ;
        RECT 206.555 128.355 206.885 128.685 ;
        RECT 206.555 126.995 206.885 127.325 ;
        RECT 206.555 125.635 206.885 125.965 ;
        RECT 206.555 124.275 206.885 124.605 ;
        RECT 206.555 121.41 206.885 121.74 ;
        RECT 206.555 119.235 206.885 119.565 ;
        RECT 206.555 117.655 206.885 117.985 ;
        RECT 206.555 116.805 206.885 117.135 ;
        RECT 206.555 114.495 206.885 114.825 ;
        RECT 206.555 113.645 206.885 113.975 ;
        RECT 206.555 111.335 206.885 111.665 ;
        RECT 206.555 110.485 206.885 110.815 ;
        RECT 206.555 108.175 206.885 108.505 ;
        RECT 206.555 107.325 206.885 107.655 ;
        RECT 206.555 105.015 206.885 105.345 ;
        RECT 206.555 103.435 206.885 103.765 ;
        RECT 206.555 102.585 206.885 102.915 ;
        RECT 206.555 100.275 206.885 100.605 ;
        RECT 206.555 99.425 206.885 99.755 ;
        RECT 206.555 97.115 206.885 97.445 ;
        RECT 206.555 96.265 206.885 96.595 ;
        RECT 206.555 93.955 206.885 94.285 ;
        RECT 206.555 93.105 206.885 93.435 ;
        RECT 206.555 90.795 206.885 91.125 ;
        RECT 206.555 89.215 206.885 89.545 ;
        RECT 206.555 88.365 206.885 88.695 ;
        RECT 206.555 86.055 206.885 86.385 ;
        RECT 206.555 85.205 206.885 85.535 ;
        RECT 206.555 82.895 206.885 83.225 ;
        RECT 206.555 82.045 206.885 82.375 ;
        RECT 206.555 79.735 206.885 80.065 ;
        RECT 206.555 78.885 206.885 79.215 ;
        RECT 206.555 76.575 206.885 76.905 ;
        RECT 206.555 74.995 206.885 75.325 ;
        RECT 206.555 74.145 206.885 74.475 ;
        RECT 206.555 71.835 206.885 72.165 ;
        RECT 206.555 70.985 206.885 71.315 ;
        RECT 206.555 68.675 206.885 69.005 ;
        RECT 206.555 67.825 206.885 68.155 ;
        RECT 206.555 65.515 206.885 65.845 ;
        RECT 206.555 64.665 206.885 64.995 ;
        RECT 206.555 62.355 206.885 62.685 ;
        RECT 206.555 60.775 206.885 61.105 ;
        RECT 206.555 59.925 206.885 60.255 ;
        RECT 206.555 57.615 206.885 57.945 ;
        RECT 206.555 56.765 206.885 57.095 ;
        RECT 206.555 54.455 206.885 54.785 ;
        RECT 206.555 53.605 206.885 53.935 ;
        RECT 206.555 51.295 206.885 51.625 ;
        RECT 206.555 50.445 206.885 50.775 ;
        RECT 206.555 48.135 206.885 48.465 ;
        RECT 206.555 46.555 206.885 46.885 ;
        RECT 206.555 45.705 206.885 46.035 ;
        RECT 206.555 43.395 206.885 43.725 ;
        RECT 206.555 42.545 206.885 42.875 ;
        RECT 206.555 40.235 206.885 40.565 ;
        RECT 206.555 39.385 206.885 39.715 ;
        RECT 206.555 37.075 206.885 37.405 ;
        RECT 206.555 36.225 206.885 36.555 ;
        RECT 206.555 33.915 206.885 34.245 ;
        RECT 206.555 32.335 206.885 32.665 ;
        RECT 206.555 31.485 206.885 31.815 ;
        RECT 206.555 29.175 206.885 29.505 ;
        RECT 206.555 28.325 206.885 28.655 ;
        RECT 206.555 26.015 206.885 26.345 ;
        RECT 206.555 25.165 206.885 25.495 ;
        RECT 206.555 22.855 206.885 23.185 ;
        RECT 206.555 22.005 206.885 22.335 ;
        RECT 206.555 19.695 206.885 20.025 ;
        RECT 206.555 18.115 206.885 18.445 ;
        RECT 206.555 17.265 206.885 17.595 ;
        RECT 206.555 14.955 206.885 15.285 ;
        RECT 206.555 14.105 206.885 14.435 ;
        RECT 206.555 11.795 206.885 12.125 ;
        RECT 206.555 10.945 206.885 11.275 ;
        RECT 206.555 8.635 206.885 8.965 ;
        RECT 206.555 7.785 206.885 8.115 ;
        RECT 206.555 5.475 206.885 5.805 ;
        RECT 206.555 3.895 206.885 4.225 ;
        RECT 206.555 3.045 206.885 3.375 ;
        RECT 206.555 0.87 206.885 1.2 ;
        RECT 206.555 -0.845 206.885 -0.515 ;
        RECT 206.555 -2.205 206.885 -1.875 ;
        RECT 206.555 -3.565 206.885 -3.235 ;
        RECT 206.555 -4.925 206.885 -4.595 ;
        RECT 206.555 -6.285 206.885 -5.955 ;
        RECT 206.555 -7.645 206.885 -7.315 ;
        RECT 206.555 -9.005 206.885 -8.675 ;
        RECT 206.555 -10.365 206.885 -10.035 ;
        RECT 206.555 -11.725 206.885 -11.395 ;
        RECT 206.555 -13.085 206.885 -12.755 ;
        RECT 206.555 -14.445 206.885 -14.115 ;
        RECT 206.555 -15.805 206.885 -15.475 ;
        RECT 206.555 -17.165 206.885 -16.835 ;
        RECT 206.555 -18.525 206.885 -18.195 ;
        RECT 206.555 -19.885 206.885 -19.555 ;
        RECT 206.555 -21.245 206.885 -20.915 ;
        RECT 206.555 -22.605 206.885 -22.275 ;
        RECT 206.555 -23.965 206.885 -23.635 ;
        RECT 206.555 -25.325 206.885 -24.995 ;
        RECT 206.555 -26.685 206.885 -26.355 ;
        RECT 206.555 -28.045 206.885 -27.715 ;
        RECT 206.555 -29.405 206.885 -29.075 ;
        RECT 206.555 -30.765 206.885 -30.435 ;
        RECT 206.555 -32.125 206.885 -31.795 ;
        RECT 206.555 -33.485 206.885 -33.155 ;
        RECT 206.555 -34.845 206.885 -34.515 ;
        RECT 206.555 -36.205 206.885 -35.875 ;
        RECT 206.555 -37.565 206.885 -37.235 ;
        RECT 206.555 -38.925 206.885 -38.595 ;
        RECT 206.555 -40.285 206.885 -39.955 ;
        RECT 206.555 -41.645 206.885 -41.315 ;
        RECT 206.555 -43.005 206.885 -42.675 ;
        RECT 206.555 -44.365 206.885 -44.035 ;
        RECT 206.555 -45.725 206.885 -45.395 ;
        RECT 206.555 -47.085 206.885 -46.755 ;
        RECT 206.555 -48.445 206.885 -48.115 ;
        RECT 206.555 -49.805 206.885 -49.475 ;
        RECT 206.555 -51.165 206.885 -50.835 ;
        RECT 206.555 -52.525 206.885 -52.195 ;
        RECT 206.555 -53.885 206.885 -53.555 ;
        RECT 206.555 -55.245 206.885 -54.915 ;
        RECT 206.555 -56.605 206.885 -56.275 ;
        RECT 206.555 -57.965 206.885 -57.635 ;
        RECT 206.555 -59.325 206.885 -58.995 ;
        RECT 206.555 -60.685 206.885 -60.355 ;
        RECT 206.555 -62.045 206.885 -61.715 ;
        RECT 206.555 -63.405 206.885 -63.075 ;
        RECT 206.555 -64.765 206.885 -64.435 ;
        RECT 206.555 -66.125 206.885 -65.795 ;
        RECT 206.555 -67.485 206.885 -67.155 ;
        RECT 206.555 -68.845 206.885 -68.515 ;
        RECT 206.555 -70.205 206.885 -69.875 ;
        RECT 206.555 -71.565 206.885 -71.235 ;
        RECT 206.555 -72.925 206.885 -72.595 ;
        RECT 206.555 -74.285 206.885 -73.955 ;
        RECT 206.555 -75.645 206.885 -75.315 ;
        RECT 206.555 -77.005 206.885 -76.675 ;
        RECT 206.555 -78.365 206.885 -78.035 ;
        RECT 206.555 -79.725 206.885 -79.395 ;
        RECT 206.555 -81.085 206.885 -80.755 ;
        RECT 206.555 -82.445 206.885 -82.115 ;
        RECT 206.555 -83.805 206.885 -83.475 ;
        RECT 206.555 -85.165 206.885 -84.835 ;
        RECT 206.555 -86.525 206.885 -86.195 ;
        RECT 206.555 -87.885 206.885 -87.555 ;
        RECT 206.555 -89.245 206.885 -88.915 ;
        RECT 206.555 -90.605 206.885 -90.275 ;
        RECT 206.555 -91.965 206.885 -91.635 ;
        RECT 206.555 -93.325 206.885 -92.995 ;
        RECT 206.555 -94.685 206.885 -94.355 ;
        RECT 206.555 -96.045 206.885 -95.715 ;
        RECT 206.555 -97.405 206.885 -97.075 ;
        RECT 206.555 -98.765 206.885 -98.435 ;
        RECT 206.555 -100.125 206.885 -99.795 ;
        RECT 206.555 -101.485 206.885 -101.155 ;
        RECT 206.555 -102.845 206.885 -102.515 ;
        RECT 206.555 -104.205 206.885 -103.875 ;
        RECT 206.555 -105.565 206.885 -105.235 ;
        RECT 206.555 -106.925 206.885 -106.595 ;
        RECT 206.555 -108.285 206.885 -107.955 ;
        RECT 206.555 -109.645 206.885 -109.315 ;
        RECT 206.555 -111.005 206.885 -110.675 ;
        RECT 206.555 -112.365 206.885 -112.035 ;
        RECT 206.555 -113.725 206.885 -113.395 ;
        RECT 206.555 -115.085 206.885 -114.755 ;
        RECT 206.555 -116.445 206.885 -116.115 ;
        RECT 206.555 -117.805 206.885 -117.475 ;
        RECT 206.555 -119.165 206.885 -118.835 ;
        RECT 206.555 -120.525 206.885 -120.195 ;
        RECT 206.555 -121.885 206.885 -121.555 ;
        RECT 206.555 -123.245 206.885 -122.915 ;
        RECT 206.555 -124.605 206.885 -124.275 ;
        RECT 206.555 -125.965 206.885 -125.635 ;
        RECT 206.555 -127.325 206.885 -126.995 ;
        RECT 206.555 -128.685 206.885 -128.355 ;
        RECT 206.555 -130.045 206.885 -129.715 ;
        RECT 206.555 -131.405 206.885 -131.075 ;
        RECT 206.555 -132.765 206.885 -132.435 ;
        RECT 206.555 -134.125 206.885 -133.795 ;
        RECT 206.555 -135.485 206.885 -135.155 ;
        RECT 206.555 -136.845 206.885 -136.515 ;
        RECT 206.555 -138.205 206.885 -137.875 ;
        RECT 206.555 -139.565 206.885 -139.235 ;
        RECT 206.555 -140.925 206.885 -140.595 ;
        RECT 206.555 -142.285 206.885 -141.955 ;
        RECT 206.555 -143.645 206.885 -143.315 ;
        RECT 206.555 -145.005 206.885 -144.675 ;
        RECT 206.555 -146.365 206.885 -146.035 ;
        RECT 206.555 -147.725 206.885 -147.395 ;
        RECT 206.555 -149.085 206.885 -148.755 ;
        RECT 206.555 -150.445 206.885 -150.115 ;
        RECT 206.555 -151.805 206.885 -151.475 ;
        RECT 206.555 -153.165 206.885 -152.835 ;
        RECT 206.555 -154.525 206.885 -154.195 ;
        RECT 206.555 -155.885 206.885 -155.555 ;
        RECT 206.555 -157.245 206.885 -156.915 ;
        RECT 206.555 -158.605 206.885 -158.275 ;
        RECT 206.555 -159.965 206.885 -159.635 ;
        RECT 206.555 -161.325 206.885 -160.995 ;
        RECT 206.555 -162.685 206.885 -162.355 ;
        RECT 206.555 -164.045 206.885 -163.715 ;
        RECT 206.555 -165.405 206.885 -165.075 ;
        RECT 206.555 -166.765 206.885 -166.435 ;
        RECT 206.555 -168.125 206.885 -167.795 ;
        RECT 206.555 -169.485 206.885 -169.155 ;
        RECT 206.555 -170.845 206.885 -170.515 ;
        RECT 206.555 -172.205 206.885 -171.875 ;
        RECT 206.555 -173.565 206.885 -173.235 ;
        RECT 206.555 -174.925 206.885 -174.595 ;
        RECT 206.555 -176.285 206.885 -175.955 ;
        RECT 206.555 -177.645 206.885 -177.315 ;
        RECT 206.555 -179.005 206.885 -178.675 ;
        RECT 206.555 -180.365 206.885 -180.035 ;
        RECT 206.555 -181.725 206.885 -181.395 ;
        RECT 206.555 -183.085 206.885 -182.755 ;
        RECT 206.555 -184.445 206.885 -184.115 ;
        RECT 206.555 -185.805 206.885 -185.475 ;
        RECT 206.555 -187.165 206.885 -186.835 ;
        RECT 206.555 -188.525 206.885 -188.195 ;
        RECT 206.555 -189.885 206.885 -189.555 ;
        RECT 206.555 -191.245 206.885 -190.915 ;
        RECT 206.555 -192.605 206.885 -192.275 ;
        RECT 206.555 -193.965 206.885 -193.635 ;
        RECT 206.555 -195.325 206.885 -194.995 ;
        RECT 206.555 -196.685 206.885 -196.355 ;
        RECT 206.555 -198.045 206.885 -197.715 ;
        RECT 206.555 -199.405 206.885 -199.075 ;
        RECT 206.555 -200.765 206.885 -200.435 ;
        RECT 206.555 -202.125 206.885 -201.795 ;
        RECT 206.555 -203.485 206.885 -203.155 ;
        RECT 206.555 -204.845 206.885 -204.515 ;
        RECT 206.555 -206.205 206.885 -205.875 ;
        RECT 206.555 -207.565 206.885 -207.235 ;
        RECT 206.555 -208.925 206.885 -208.595 ;
        RECT 206.555 -210.285 206.885 -209.955 ;
        RECT 206.555 -211.645 206.885 -211.315 ;
        RECT 206.555 -213.005 206.885 -212.675 ;
        RECT 206.555 -214.365 206.885 -214.035 ;
        RECT 206.555 -215.725 206.885 -215.395 ;
        RECT 206.555 -217.085 206.885 -216.755 ;
        RECT 206.555 -218.445 206.885 -218.115 ;
        RECT 206.555 -224.09 206.885 -222.96 ;
        RECT 206.56 -224.205 206.88 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.915 132.52 208.245 133.65 ;
        RECT 207.915 128.355 208.245 128.685 ;
        RECT 207.915 126.995 208.245 127.325 ;
        RECT 207.915 125.635 208.245 125.965 ;
        RECT 207.915 124.275 208.245 124.605 ;
        RECT 207.915 122.915 208.245 123.245 ;
        RECT 207.915 121.555 208.245 121.885 ;
        RECT 207.915 120.195 208.245 120.525 ;
        RECT 207.915 118.835 208.245 119.165 ;
        RECT 207.915 117.475 208.245 117.805 ;
        RECT 207.915 116.115 208.245 116.445 ;
        RECT 207.915 114.755 208.245 115.085 ;
        RECT 207.915 113.395 208.245 113.725 ;
        RECT 207.915 112.035 208.245 112.365 ;
        RECT 207.915 110.675 208.245 111.005 ;
        RECT 207.915 109.315 208.245 109.645 ;
        RECT 207.915 107.955 208.245 108.285 ;
        RECT 207.915 106.595 208.245 106.925 ;
        RECT 207.915 105.235 208.245 105.565 ;
        RECT 207.915 103.875 208.245 104.205 ;
        RECT 207.915 102.515 208.245 102.845 ;
        RECT 207.915 101.155 208.245 101.485 ;
        RECT 207.915 99.795 208.245 100.125 ;
        RECT 207.915 98.435 208.245 98.765 ;
        RECT 207.915 97.075 208.245 97.405 ;
        RECT 207.915 95.715 208.245 96.045 ;
        RECT 207.915 94.355 208.245 94.685 ;
        RECT 207.915 92.995 208.245 93.325 ;
        RECT 207.915 91.635 208.245 91.965 ;
        RECT 207.915 90.275 208.245 90.605 ;
        RECT 207.915 88.915 208.245 89.245 ;
        RECT 207.915 87.555 208.245 87.885 ;
        RECT 207.915 86.195 208.245 86.525 ;
        RECT 207.915 84.835 208.245 85.165 ;
        RECT 207.915 83.475 208.245 83.805 ;
        RECT 207.915 82.115 208.245 82.445 ;
        RECT 207.915 80.755 208.245 81.085 ;
        RECT 207.915 79.395 208.245 79.725 ;
        RECT 207.915 78.035 208.245 78.365 ;
        RECT 207.915 76.675 208.245 77.005 ;
        RECT 207.915 75.315 208.245 75.645 ;
        RECT 207.915 73.955 208.245 74.285 ;
        RECT 207.915 72.595 208.245 72.925 ;
        RECT 207.915 71.235 208.245 71.565 ;
        RECT 207.915 69.875 208.245 70.205 ;
        RECT 207.915 68.515 208.245 68.845 ;
        RECT 207.915 67.155 208.245 67.485 ;
        RECT 207.915 65.795 208.245 66.125 ;
        RECT 207.915 64.435 208.245 64.765 ;
        RECT 207.915 63.075 208.245 63.405 ;
        RECT 207.915 61.715 208.245 62.045 ;
        RECT 207.915 60.355 208.245 60.685 ;
        RECT 207.915 58.995 208.245 59.325 ;
        RECT 207.915 57.635 208.245 57.965 ;
        RECT 207.915 56.275 208.245 56.605 ;
        RECT 207.915 54.915 208.245 55.245 ;
        RECT 207.915 53.555 208.245 53.885 ;
        RECT 207.915 52.195 208.245 52.525 ;
        RECT 207.915 50.835 208.245 51.165 ;
        RECT 207.915 49.475 208.245 49.805 ;
        RECT 207.915 48.115 208.245 48.445 ;
        RECT 207.915 46.755 208.245 47.085 ;
        RECT 207.915 45.395 208.245 45.725 ;
        RECT 207.915 44.035 208.245 44.365 ;
        RECT 207.915 42.675 208.245 43.005 ;
        RECT 207.915 41.315 208.245 41.645 ;
        RECT 207.915 39.955 208.245 40.285 ;
        RECT 207.915 38.595 208.245 38.925 ;
        RECT 207.915 37.235 208.245 37.565 ;
        RECT 207.915 35.875 208.245 36.205 ;
        RECT 207.915 34.515 208.245 34.845 ;
        RECT 207.915 33.155 208.245 33.485 ;
        RECT 207.915 31.795 208.245 32.125 ;
        RECT 207.915 30.435 208.245 30.765 ;
        RECT 207.915 29.075 208.245 29.405 ;
        RECT 207.915 27.715 208.245 28.045 ;
        RECT 207.915 26.355 208.245 26.685 ;
        RECT 207.915 24.995 208.245 25.325 ;
        RECT 207.915 23.635 208.245 23.965 ;
        RECT 207.915 22.275 208.245 22.605 ;
        RECT 207.915 20.915 208.245 21.245 ;
        RECT 207.915 19.555 208.245 19.885 ;
        RECT 207.915 18.195 208.245 18.525 ;
        RECT 207.915 16.835 208.245 17.165 ;
        RECT 207.915 15.475 208.245 15.805 ;
        RECT 207.915 14.115 208.245 14.445 ;
        RECT 207.915 12.755 208.245 13.085 ;
        RECT 207.915 11.395 208.245 11.725 ;
        RECT 207.915 10.035 208.245 10.365 ;
        RECT 207.915 8.675 208.245 9.005 ;
        RECT 207.915 7.315 208.245 7.645 ;
        RECT 207.915 5.955 208.245 6.285 ;
        RECT 207.915 4.595 208.245 4.925 ;
        RECT 207.915 3.235 208.245 3.565 ;
        RECT 207.915 1.875 208.245 2.205 ;
        RECT 207.915 0.515 208.245 0.845 ;
        RECT 207.915 -0.845 208.245 -0.515 ;
        RECT 207.915 -2.205 208.245 -1.875 ;
        RECT 207.915 -3.565 208.245 -3.235 ;
        RECT 207.915 -4.925 208.245 -4.595 ;
        RECT 207.915 -6.285 208.245 -5.955 ;
        RECT 207.915 -7.645 208.245 -7.315 ;
        RECT 207.915 -9.005 208.245 -8.675 ;
        RECT 207.915 -10.365 208.245 -10.035 ;
        RECT 207.915 -11.725 208.245 -11.395 ;
        RECT 207.915 -13.085 208.245 -12.755 ;
        RECT 207.915 -14.445 208.245 -14.115 ;
        RECT 207.915 -15.805 208.245 -15.475 ;
        RECT 207.915 -17.165 208.245 -16.835 ;
        RECT 207.915 -18.525 208.245 -18.195 ;
        RECT 207.915 -19.885 208.245 -19.555 ;
        RECT 207.915 -21.245 208.245 -20.915 ;
        RECT 207.915 -22.605 208.245 -22.275 ;
        RECT 207.915 -23.965 208.245 -23.635 ;
        RECT 207.915 -25.325 208.245 -24.995 ;
        RECT 207.915 -26.685 208.245 -26.355 ;
        RECT 207.915 -28.045 208.245 -27.715 ;
        RECT 207.915 -29.405 208.245 -29.075 ;
        RECT 207.915 -30.765 208.245 -30.435 ;
        RECT 207.915 -32.125 208.245 -31.795 ;
        RECT 207.915 -33.485 208.245 -33.155 ;
        RECT 207.915 -34.845 208.245 -34.515 ;
        RECT 207.915 -36.205 208.245 -35.875 ;
        RECT 207.915 -37.565 208.245 -37.235 ;
        RECT 207.915 -38.925 208.245 -38.595 ;
        RECT 207.915 -40.285 208.245 -39.955 ;
        RECT 207.915 -41.645 208.245 -41.315 ;
        RECT 207.915 -43.005 208.245 -42.675 ;
        RECT 207.915 -44.365 208.245 -44.035 ;
        RECT 207.915 -45.725 208.245 -45.395 ;
        RECT 207.915 -47.085 208.245 -46.755 ;
        RECT 207.915 -48.445 208.245 -48.115 ;
        RECT 207.915 -49.805 208.245 -49.475 ;
        RECT 207.915 -51.165 208.245 -50.835 ;
        RECT 207.915 -52.525 208.245 -52.195 ;
        RECT 207.915 -53.885 208.245 -53.555 ;
        RECT 207.915 -55.245 208.245 -54.915 ;
        RECT 207.915 -56.605 208.245 -56.275 ;
        RECT 207.915 -57.965 208.245 -57.635 ;
        RECT 207.915 -59.325 208.245 -58.995 ;
        RECT 207.915 -60.685 208.245 -60.355 ;
        RECT 207.915 -62.045 208.245 -61.715 ;
        RECT 207.915 -63.405 208.245 -63.075 ;
        RECT 207.915 -64.765 208.245 -64.435 ;
        RECT 207.915 -66.125 208.245 -65.795 ;
        RECT 207.915 -67.485 208.245 -67.155 ;
        RECT 207.915 -68.845 208.245 -68.515 ;
        RECT 207.915 -70.205 208.245 -69.875 ;
        RECT 207.915 -71.565 208.245 -71.235 ;
        RECT 207.915 -72.925 208.245 -72.595 ;
        RECT 207.915 -74.285 208.245 -73.955 ;
        RECT 207.915 -75.645 208.245 -75.315 ;
        RECT 207.915 -77.005 208.245 -76.675 ;
        RECT 207.915 -78.365 208.245 -78.035 ;
        RECT 207.915 -79.725 208.245 -79.395 ;
        RECT 207.915 -81.085 208.245 -80.755 ;
        RECT 207.915 -82.445 208.245 -82.115 ;
        RECT 207.915 -83.805 208.245 -83.475 ;
        RECT 207.915 -85.165 208.245 -84.835 ;
        RECT 207.915 -86.525 208.245 -86.195 ;
        RECT 207.915 -87.885 208.245 -87.555 ;
        RECT 207.915 -89.245 208.245 -88.915 ;
        RECT 207.915 -90.605 208.245 -90.275 ;
        RECT 207.915 -91.965 208.245 -91.635 ;
        RECT 207.915 -93.325 208.245 -92.995 ;
        RECT 207.915 -94.685 208.245 -94.355 ;
        RECT 207.915 -96.045 208.245 -95.715 ;
        RECT 207.915 -97.405 208.245 -97.075 ;
        RECT 207.915 -98.765 208.245 -98.435 ;
        RECT 207.915 -100.125 208.245 -99.795 ;
        RECT 207.915 -101.485 208.245 -101.155 ;
        RECT 207.915 -102.845 208.245 -102.515 ;
        RECT 207.915 -104.205 208.245 -103.875 ;
        RECT 207.915 -105.565 208.245 -105.235 ;
        RECT 207.915 -106.925 208.245 -106.595 ;
        RECT 207.915 -108.285 208.245 -107.955 ;
        RECT 207.915 -109.645 208.245 -109.315 ;
        RECT 207.915 -111.005 208.245 -110.675 ;
        RECT 207.915 -112.365 208.245 -112.035 ;
        RECT 207.915 -113.725 208.245 -113.395 ;
        RECT 207.915 -115.085 208.245 -114.755 ;
        RECT 207.915 -116.445 208.245 -116.115 ;
        RECT 207.915 -117.805 208.245 -117.475 ;
        RECT 207.915 -119.165 208.245 -118.835 ;
        RECT 207.915 -120.525 208.245 -120.195 ;
        RECT 207.915 -121.885 208.245 -121.555 ;
        RECT 207.915 -123.245 208.245 -122.915 ;
        RECT 207.915 -124.605 208.245 -124.275 ;
        RECT 207.915 -125.965 208.245 -125.635 ;
        RECT 207.915 -127.325 208.245 -126.995 ;
        RECT 207.915 -128.685 208.245 -128.355 ;
        RECT 207.915 -130.045 208.245 -129.715 ;
        RECT 207.915 -131.405 208.245 -131.075 ;
        RECT 207.915 -132.765 208.245 -132.435 ;
        RECT 207.915 -134.125 208.245 -133.795 ;
        RECT 207.915 -135.485 208.245 -135.155 ;
        RECT 207.915 -136.845 208.245 -136.515 ;
        RECT 207.915 -138.205 208.245 -137.875 ;
        RECT 207.915 -139.565 208.245 -139.235 ;
        RECT 207.915 -140.925 208.245 -140.595 ;
        RECT 207.915 -142.285 208.245 -141.955 ;
        RECT 207.915 -143.645 208.245 -143.315 ;
        RECT 207.915 -145.005 208.245 -144.675 ;
        RECT 207.915 -146.365 208.245 -146.035 ;
        RECT 207.915 -147.725 208.245 -147.395 ;
        RECT 207.915 -149.085 208.245 -148.755 ;
        RECT 207.915 -150.445 208.245 -150.115 ;
        RECT 207.915 -151.805 208.245 -151.475 ;
        RECT 207.915 -153.165 208.245 -152.835 ;
        RECT 207.915 -154.525 208.245 -154.195 ;
        RECT 207.915 -155.885 208.245 -155.555 ;
        RECT 207.915 -157.245 208.245 -156.915 ;
        RECT 207.915 -158.605 208.245 -158.275 ;
        RECT 207.915 -159.965 208.245 -159.635 ;
        RECT 207.915 -161.325 208.245 -160.995 ;
        RECT 207.915 -162.685 208.245 -162.355 ;
        RECT 207.915 -164.045 208.245 -163.715 ;
        RECT 207.915 -165.405 208.245 -165.075 ;
        RECT 207.915 -166.765 208.245 -166.435 ;
        RECT 207.915 -168.125 208.245 -167.795 ;
        RECT 207.915 -169.485 208.245 -169.155 ;
        RECT 207.915 -170.845 208.245 -170.515 ;
        RECT 207.915 -172.205 208.245 -171.875 ;
        RECT 207.915 -173.565 208.245 -173.235 ;
        RECT 207.915 -174.925 208.245 -174.595 ;
        RECT 207.915 -176.285 208.245 -175.955 ;
        RECT 207.915 -177.645 208.245 -177.315 ;
        RECT 207.915 -179.005 208.245 -178.675 ;
        RECT 207.915 -180.365 208.245 -180.035 ;
        RECT 207.915 -181.725 208.245 -181.395 ;
        RECT 207.915 -183.085 208.245 -182.755 ;
        RECT 207.915 -184.445 208.245 -184.115 ;
        RECT 207.915 -185.805 208.245 -185.475 ;
        RECT 207.915 -187.165 208.245 -186.835 ;
        RECT 207.915 -188.525 208.245 -188.195 ;
        RECT 207.915 -189.885 208.245 -189.555 ;
        RECT 207.915 -191.245 208.245 -190.915 ;
        RECT 207.915 -192.605 208.245 -192.275 ;
        RECT 207.915 -193.965 208.245 -193.635 ;
        RECT 207.915 -195.325 208.245 -194.995 ;
        RECT 207.915 -196.685 208.245 -196.355 ;
        RECT 207.915 -198.045 208.245 -197.715 ;
        RECT 207.915 -199.405 208.245 -199.075 ;
        RECT 207.915 -200.765 208.245 -200.435 ;
        RECT 207.915 -202.125 208.245 -201.795 ;
        RECT 207.915 -203.485 208.245 -203.155 ;
        RECT 207.915 -204.845 208.245 -204.515 ;
        RECT 207.915 -206.205 208.245 -205.875 ;
        RECT 207.915 -207.565 208.245 -207.235 ;
        RECT 207.915 -208.925 208.245 -208.595 ;
        RECT 207.915 -210.285 208.245 -209.955 ;
        RECT 207.915 -211.645 208.245 -211.315 ;
        RECT 207.915 -213.005 208.245 -212.675 ;
        RECT 207.915 -214.365 208.245 -214.035 ;
        RECT 207.915 -215.725 208.245 -215.395 ;
        RECT 207.915 -217.085 208.245 -216.755 ;
        RECT 207.915 -218.445 208.245 -218.115 ;
        RECT 207.915 -224.09 208.245 -222.96 ;
        RECT 207.92 -224.205 208.24 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.275 132.52 209.605 133.65 ;
        RECT 209.275 128.355 209.605 128.685 ;
        RECT 209.275 126.995 209.605 127.325 ;
        RECT 209.275 125.635 209.605 125.965 ;
        RECT 209.275 124.275 209.605 124.605 ;
        RECT 209.275 122.915 209.605 123.245 ;
        RECT 209.275 121.555 209.605 121.885 ;
        RECT 209.275 120.195 209.605 120.525 ;
        RECT 209.275 118.835 209.605 119.165 ;
        RECT 209.275 117.475 209.605 117.805 ;
        RECT 209.275 116.115 209.605 116.445 ;
        RECT 209.275 114.755 209.605 115.085 ;
        RECT 209.275 113.395 209.605 113.725 ;
        RECT 209.275 112.035 209.605 112.365 ;
        RECT 209.275 110.675 209.605 111.005 ;
        RECT 209.275 109.315 209.605 109.645 ;
        RECT 209.275 107.955 209.605 108.285 ;
        RECT 209.275 106.595 209.605 106.925 ;
        RECT 209.275 105.235 209.605 105.565 ;
        RECT 209.275 103.875 209.605 104.205 ;
        RECT 209.275 102.515 209.605 102.845 ;
        RECT 209.275 101.155 209.605 101.485 ;
        RECT 209.275 99.795 209.605 100.125 ;
        RECT 209.275 98.435 209.605 98.765 ;
        RECT 209.275 97.075 209.605 97.405 ;
        RECT 209.275 95.715 209.605 96.045 ;
        RECT 209.275 94.355 209.605 94.685 ;
        RECT 209.275 92.995 209.605 93.325 ;
        RECT 209.275 91.635 209.605 91.965 ;
        RECT 209.275 90.275 209.605 90.605 ;
        RECT 209.275 88.915 209.605 89.245 ;
        RECT 209.275 87.555 209.605 87.885 ;
        RECT 209.275 86.195 209.605 86.525 ;
        RECT 209.275 84.835 209.605 85.165 ;
        RECT 209.275 83.475 209.605 83.805 ;
        RECT 209.275 82.115 209.605 82.445 ;
        RECT 209.275 80.755 209.605 81.085 ;
        RECT 209.275 79.395 209.605 79.725 ;
        RECT 209.275 78.035 209.605 78.365 ;
        RECT 209.275 76.675 209.605 77.005 ;
        RECT 209.275 75.315 209.605 75.645 ;
        RECT 209.275 73.955 209.605 74.285 ;
        RECT 209.275 72.595 209.605 72.925 ;
        RECT 209.275 71.235 209.605 71.565 ;
        RECT 209.275 69.875 209.605 70.205 ;
        RECT 209.275 68.515 209.605 68.845 ;
        RECT 209.275 67.155 209.605 67.485 ;
        RECT 209.275 65.795 209.605 66.125 ;
        RECT 209.275 64.435 209.605 64.765 ;
        RECT 209.275 63.075 209.605 63.405 ;
        RECT 209.275 61.715 209.605 62.045 ;
        RECT 209.275 60.355 209.605 60.685 ;
        RECT 209.275 58.995 209.605 59.325 ;
        RECT 209.275 57.635 209.605 57.965 ;
        RECT 209.275 56.275 209.605 56.605 ;
        RECT 209.275 54.915 209.605 55.245 ;
        RECT 209.275 53.555 209.605 53.885 ;
        RECT 209.275 52.195 209.605 52.525 ;
        RECT 209.275 50.835 209.605 51.165 ;
        RECT 209.275 49.475 209.605 49.805 ;
        RECT 209.275 48.115 209.605 48.445 ;
        RECT 209.275 46.755 209.605 47.085 ;
        RECT 209.275 45.395 209.605 45.725 ;
        RECT 209.275 44.035 209.605 44.365 ;
        RECT 209.275 42.675 209.605 43.005 ;
        RECT 209.275 41.315 209.605 41.645 ;
        RECT 209.275 39.955 209.605 40.285 ;
        RECT 209.275 38.595 209.605 38.925 ;
        RECT 209.275 37.235 209.605 37.565 ;
        RECT 209.275 35.875 209.605 36.205 ;
        RECT 209.275 34.515 209.605 34.845 ;
        RECT 209.275 33.155 209.605 33.485 ;
        RECT 209.275 31.795 209.605 32.125 ;
        RECT 209.275 30.435 209.605 30.765 ;
        RECT 209.275 29.075 209.605 29.405 ;
        RECT 209.275 27.715 209.605 28.045 ;
        RECT 209.275 26.355 209.605 26.685 ;
        RECT 209.275 24.995 209.605 25.325 ;
        RECT 209.275 23.635 209.605 23.965 ;
        RECT 209.275 22.275 209.605 22.605 ;
        RECT 209.275 20.915 209.605 21.245 ;
        RECT 209.275 19.555 209.605 19.885 ;
        RECT 209.275 18.195 209.605 18.525 ;
        RECT 209.275 16.835 209.605 17.165 ;
        RECT 209.275 15.475 209.605 15.805 ;
        RECT 209.275 14.115 209.605 14.445 ;
        RECT 209.275 12.755 209.605 13.085 ;
        RECT 209.275 11.395 209.605 11.725 ;
        RECT 209.275 10.035 209.605 10.365 ;
        RECT 209.275 8.675 209.605 9.005 ;
        RECT 209.275 7.315 209.605 7.645 ;
        RECT 209.275 5.955 209.605 6.285 ;
        RECT 209.275 4.595 209.605 4.925 ;
        RECT 209.275 3.235 209.605 3.565 ;
        RECT 209.275 1.875 209.605 2.205 ;
        RECT 209.275 0.515 209.605 0.845 ;
        RECT 209.275 -0.845 209.605 -0.515 ;
        RECT 209.275 -2.205 209.605 -1.875 ;
        RECT 209.275 -3.565 209.605 -3.235 ;
        RECT 209.275 -4.925 209.605 -4.595 ;
        RECT 209.275 -6.285 209.605 -5.955 ;
        RECT 209.275 -7.645 209.605 -7.315 ;
        RECT 209.275 -9.005 209.605 -8.675 ;
        RECT 209.275 -10.365 209.605 -10.035 ;
        RECT 209.275 -11.725 209.605 -11.395 ;
        RECT 209.275 -13.085 209.605 -12.755 ;
        RECT 209.275 -14.445 209.605 -14.115 ;
        RECT 209.275 -15.805 209.605 -15.475 ;
        RECT 209.275 -17.165 209.605 -16.835 ;
        RECT 209.275 -18.525 209.605 -18.195 ;
        RECT 209.275 -19.885 209.605 -19.555 ;
        RECT 209.275 -21.245 209.605 -20.915 ;
        RECT 209.275 -22.605 209.605 -22.275 ;
        RECT 209.275 -23.965 209.605 -23.635 ;
        RECT 209.275 -25.325 209.605 -24.995 ;
        RECT 209.275 -26.685 209.605 -26.355 ;
        RECT 209.275 -28.045 209.605 -27.715 ;
        RECT 209.275 -29.405 209.605 -29.075 ;
        RECT 209.275 -30.765 209.605 -30.435 ;
        RECT 209.275 -32.125 209.605 -31.795 ;
        RECT 209.275 -33.485 209.605 -33.155 ;
        RECT 209.275 -34.845 209.605 -34.515 ;
        RECT 209.275 -36.205 209.605 -35.875 ;
        RECT 209.275 -37.565 209.605 -37.235 ;
        RECT 209.275 -38.925 209.605 -38.595 ;
        RECT 209.275 -40.285 209.605 -39.955 ;
        RECT 209.275 -41.645 209.605 -41.315 ;
        RECT 209.275 -43.005 209.605 -42.675 ;
        RECT 209.275 -44.365 209.605 -44.035 ;
        RECT 209.275 -45.725 209.605 -45.395 ;
        RECT 209.275 -47.085 209.605 -46.755 ;
        RECT 209.275 -48.445 209.605 -48.115 ;
        RECT 209.275 -49.805 209.605 -49.475 ;
        RECT 209.275 -51.165 209.605 -50.835 ;
        RECT 209.275 -52.525 209.605 -52.195 ;
        RECT 209.275 -53.885 209.605 -53.555 ;
        RECT 209.275 -55.245 209.605 -54.915 ;
        RECT 209.275 -56.605 209.605 -56.275 ;
        RECT 209.275 -57.965 209.605 -57.635 ;
        RECT 209.275 -59.325 209.605 -58.995 ;
        RECT 209.275 -60.685 209.605 -60.355 ;
        RECT 209.275 -62.045 209.605 -61.715 ;
        RECT 209.275 -63.405 209.605 -63.075 ;
        RECT 209.275 -64.765 209.605 -64.435 ;
        RECT 209.275 -66.125 209.605 -65.795 ;
        RECT 209.275 -67.485 209.605 -67.155 ;
        RECT 209.275 -68.845 209.605 -68.515 ;
        RECT 209.275 -70.205 209.605 -69.875 ;
        RECT 209.275 -71.565 209.605 -71.235 ;
        RECT 209.275 -72.925 209.605 -72.595 ;
        RECT 209.275 -74.285 209.605 -73.955 ;
        RECT 209.275 -75.645 209.605 -75.315 ;
        RECT 209.275 -77.005 209.605 -76.675 ;
        RECT 209.275 -78.365 209.605 -78.035 ;
        RECT 209.275 -79.725 209.605 -79.395 ;
        RECT 209.275 -81.085 209.605 -80.755 ;
        RECT 209.275 -82.445 209.605 -82.115 ;
        RECT 209.275 -83.805 209.605 -83.475 ;
        RECT 209.275 -85.165 209.605 -84.835 ;
        RECT 209.275 -86.525 209.605 -86.195 ;
        RECT 209.275 -87.885 209.605 -87.555 ;
        RECT 209.275 -89.245 209.605 -88.915 ;
        RECT 209.275 -90.605 209.605 -90.275 ;
        RECT 209.275 -91.965 209.605 -91.635 ;
        RECT 209.275 -93.325 209.605 -92.995 ;
        RECT 209.275 -94.685 209.605 -94.355 ;
        RECT 209.275 -96.045 209.605 -95.715 ;
        RECT 209.275 -97.405 209.605 -97.075 ;
        RECT 209.275 -98.765 209.605 -98.435 ;
        RECT 209.275 -100.125 209.605 -99.795 ;
        RECT 209.275 -101.485 209.605 -101.155 ;
        RECT 209.275 -102.845 209.605 -102.515 ;
        RECT 209.275 -104.205 209.605 -103.875 ;
        RECT 209.275 -105.565 209.605 -105.235 ;
        RECT 209.275 -106.925 209.605 -106.595 ;
        RECT 209.275 -108.285 209.605 -107.955 ;
        RECT 209.275 -109.645 209.605 -109.315 ;
        RECT 209.275 -111.005 209.605 -110.675 ;
        RECT 209.275 -112.365 209.605 -112.035 ;
        RECT 209.275 -113.725 209.605 -113.395 ;
        RECT 209.275 -115.085 209.605 -114.755 ;
        RECT 209.275 -116.445 209.605 -116.115 ;
        RECT 209.275 -117.805 209.605 -117.475 ;
        RECT 209.275 -119.165 209.605 -118.835 ;
        RECT 209.275 -120.525 209.605 -120.195 ;
        RECT 209.275 -121.885 209.605 -121.555 ;
        RECT 209.275 -123.245 209.605 -122.915 ;
        RECT 209.275 -124.605 209.605 -124.275 ;
        RECT 209.275 -125.965 209.605 -125.635 ;
        RECT 209.275 -127.325 209.605 -126.995 ;
        RECT 209.275 -128.685 209.605 -128.355 ;
        RECT 209.275 -130.045 209.605 -129.715 ;
        RECT 209.275 -131.405 209.605 -131.075 ;
        RECT 209.275 -132.765 209.605 -132.435 ;
        RECT 209.275 -134.125 209.605 -133.795 ;
        RECT 209.275 -135.485 209.605 -135.155 ;
        RECT 209.275 -136.845 209.605 -136.515 ;
        RECT 209.275 -138.205 209.605 -137.875 ;
        RECT 209.275 -139.565 209.605 -139.235 ;
        RECT 209.275 -140.925 209.605 -140.595 ;
        RECT 209.275 -142.285 209.605 -141.955 ;
        RECT 209.275 -143.645 209.605 -143.315 ;
        RECT 209.275 -145.005 209.605 -144.675 ;
        RECT 209.275 -146.365 209.605 -146.035 ;
        RECT 209.275 -147.725 209.605 -147.395 ;
        RECT 209.275 -149.085 209.605 -148.755 ;
        RECT 209.275 -150.445 209.605 -150.115 ;
        RECT 209.275 -151.805 209.605 -151.475 ;
        RECT 209.275 -153.165 209.605 -152.835 ;
        RECT 209.275 -154.525 209.605 -154.195 ;
        RECT 209.275 -155.885 209.605 -155.555 ;
        RECT 209.275 -157.245 209.605 -156.915 ;
        RECT 209.275 -158.605 209.605 -158.275 ;
        RECT 209.275 -159.965 209.605 -159.635 ;
        RECT 209.275 -161.325 209.605 -160.995 ;
        RECT 209.275 -162.685 209.605 -162.355 ;
        RECT 209.275 -164.045 209.605 -163.715 ;
        RECT 209.275 -165.405 209.605 -165.075 ;
        RECT 209.275 -166.765 209.605 -166.435 ;
        RECT 209.275 -168.125 209.605 -167.795 ;
        RECT 209.275 -169.485 209.605 -169.155 ;
        RECT 209.275 -170.845 209.605 -170.515 ;
        RECT 209.275 -172.205 209.605 -171.875 ;
        RECT 209.275 -173.565 209.605 -173.235 ;
        RECT 209.275 -174.925 209.605 -174.595 ;
        RECT 209.275 -176.285 209.605 -175.955 ;
        RECT 209.275 -177.645 209.605 -177.315 ;
        RECT 209.275 -179.005 209.605 -178.675 ;
        RECT 209.275 -180.365 209.605 -180.035 ;
        RECT 209.275 -181.725 209.605 -181.395 ;
        RECT 209.275 -183.085 209.605 -182.755 ;
        RECT 209.275 -184.445 209.605 -184.115 ;
        RECT 209.275 -185.805 209.605 -185.475 ;
        RECT 209.275 -187.165 209.605 -186.835 ;
        RECT 209.275 -188.525 209.605 -188.195 ;
        RECT 209.275 -189.885 209.605 -189.555 ;
        RECT 209.275 -191.245 209.605 -190.915 ;
        RECT 209.275 -192.605 209.605 -192.275 ;
        RECT 209.275 -193.965 209.605 -193.635 ;
        RECT 209.275 -195.325 209.605 -194.995 ;
        RECT 209.275 -196.685 209.605 -196.355 ;
        RECT 209.275 -198.045 209.605 -197.715 ;
        RECT 209.275 -199.405 209.605 -199.075 ;
        RECT 209.275 -200.765 209.605 -200.435 ;
        RECT 209.275 -202.125 209.605 -201.795 ;
        RECT 209.275 -203.485 209.605 -203.155 ;
        RECT 209.275 -204.845 209.605 -204.515 ;
        RECT 209.275 -206.205 209.605 -205.875 ;
        RECT 209.275 -207.565 209.605 -207.235 ;
        RECT 209.275 -208.925 209.605 -208.595 ;
        RECT 209.275 -210.285 209.605 -209.955 ;
        RECT 209.275 -211.645 209.605 -211.315 ;
        RECT 209.275 -213.005 209.605 -212.675 ;
        RECT 209.275 -214.365 209.605 -214.035 ;
        RECT 209.275 -215.725 209.605 -215.395 ;
        RECT 209.275 -217.085 209.605 -216.755 ;
        RECT 209.275 -218.445 209.605 -218.115 ;
        RECT 209.275 -224.09 209.605 -222.96 ;
        RECT 209.28 -224.205 209.6 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 191.76 -121.535 192.09 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.955 132.52 193.285 133.65 ;
        RECT 192.955 128.355 193.285 128.685 ;
        RECT 192.955 126.995 193.285 127.325 ;
        RECT 192.955 125.635 193.285 125.965 ;
        RECT 192.955 124.275 193.285 124.605 ;
        RECT 192.96 123.6 193.28 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.315 132.52 194.645 133.65 ;
        RECT 194.315 128.355 194.645 128.685 ;
        RECT 194.315 126.995 194.645 127.325 ;
        RECT 194.315 125.635 194.645 125.965 ;
        RECT 194.315 124.275 194.645 124.605 ;
        RECT 194.32 123.6 194.64 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.315 -0.845 194.645 -0.515 ;
        RECT 194.315 -2.205 194.645 -1.875 ;
        RECT 194.315 -3.565 194.645 -3.235 ;
        RECT 194.32 -3.565 194.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.675 132.52 196.005 133.65 ;
        RECT 195.675 128.355 196.005 128.685 ;
        RECT 195.675 126.995 196.005 127.325 ;
        RECT 195.675 125.635 196.005 125.965 ;
        RECT 195.675 124.275 196.005 124.605 ;
        RECT 195.68 123.6 196 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.675 -0.845 196.005 -0.515 ;
        RECT 195.675 -2.205 196.005 -1.875 ;
        RECT 195.675 -3.565 196.005 -3.235 ;
        RECT 195.68 -3.565 196 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.675 -119.165 196.005 -118.835 ;
        RECT 195.675 -120.525 196.005 -120.195 ;
        RECT 195.675 -121.885 196.005 -121.555 ;
        RECT 195.675 -123.245 196.005 -122.915 ;
        RECT 195.675 -124.605 196.005 -124.275 ;
        RECT 195.675 -125.965 196.005 -125.635 ;
        RECT 195.675 -127.325 196.005 -126.995 ;
        RECT 195.675 -128.685 196.005 -128.355 ;
        RECT 195.675 -130.045 196.005 -129.715 ;
        RECT 195.675 -131.405 196.005 -131.075 ;
        RECT 195.675 -132.765 196.005 -132.435 ;
        RECT 195.675 -134.125 196.005 -133.795 ;
        RECT 195.675 -135.485 196.005 -135.155 ;
        RECT 195.675 -136.845 196.005 -136.515 ;
        RECT 195.675 -138.205 196.005 -137.875 ;
        RECT 195.675 -139.565 196.005 -139.235 ;
        RECT 195.675 -140.925 196.005 -140.595 ;
        RECT 195.675 -142.285 196.005 -141.955 ;
        RECT 195.675 -143.645 196.005 -143.315 ;
        RECT 195.675 -145.005 196.005 -144.675 ;
        RECT 195.675 -146.365 196.005 -146.035 ;
        RECT 195.675 -147.725 196.005 -147.395 ;
        RECT 195.675 -149.085 196.005 -148.755 ;
        RECT 195.675 -150.445 196.005 -150.115 ;
        RECT 195.675 -151.805 196.005 -151.475 ;
        RECT 195.675 -153.165 196.005 -152.835 ;
        RECT 195.675 -154.525 196.005 -154.195 ;
        RECT 195.675 -155.885 196.005 -155.555 ;
        RECT 195.675 -157.245 196.005 -156.915 ;
        RECT 195.675 -158.605 196.005 -158.275 ;
        RECT 195.675 -159.965 196.005 -159.635 ;
        RECT 195.675 -161.325 196.005 -160.995 ;
        RECT 195.675 -162.685 196.005 -162.355 ;
        RECT 195.675 -164.045 196.005 -163.715 ;
        RECT 195.675 -165.405 196.005 -165.075 ;
        RECT 195.675 -166.765 196.005 -166.435 ;
        RECT 195.675 -168.125 196.005 -167.795 ;
        RECT 195.675 -169.485 196.005 -169.155 ;
        RECT 195.675 -170.845 196.005 -170.515 ;
        RECT 195.675 -172.205 196.005 -171.875 ;
        RECT 195.675 -173.565 196.005 -173.235 ;
        RECT 195.675 -174.925 196.005 -174.595 ;
        RECT 195.675 -176.285 196.005 -175.955 ;
        RECT 195.675 -177.645 196.005 -177.315 ;
        RECT 195.675 -179.005 196.005 -178.675 ;
        RECT 195.675 -180.365 196.005 -180.035 ;
        RECT 195.675 -181.725 196.005 -181.395 ;
        RECT 195.675 -183.085 196.005 -182.755 ;
        RECT 195.675 -184.445 196.005 -184.115 ;
        RECT 195.675 -185.805 196.005 -185.475 ;
        RECT 195.675 -187.165 196.005 -186.835 ;
        RECT 195.675 -188.525 196.005 -188.195 ;
        RECT 195.675 -189.885 196.005 -189.555 ;
        RECT 195.675 -191.245 196.005 -190.915 ;
        RECT 195.675 -192.605 196.005 -192.275 ;
        RECT 195.675 -193.965 196.005 -193.635 ;
        RECT 195.675 -195.325 196.005 -194.995 ;
        RECT 195.675 -196.685 196.005 -196.355 ;
        RECT 195.675 -198.045 196.005 -197.715 ;
        RECT 195.675 -199.405 196.005 -199.075 ;
        RECT 195.675 -200.765 196.005 -200.435 ;
        RECT 195.675 -202.125 196.005 -201.795 ;
        RECT 195.675 -203.485 196.005 -203.155 ;
        RECT 195.675 -204.845 196.005 -204.515 ;
        RECT 195.675 -206.205 196.005 -205.875 ;
        RECT 195.675 -207.565 196.005 -207.235 ;
        RECT 195.675 -208.925 196.005 -208.595 ;
        RECT 195.675 -210.285 196.005 -209.955 ;
        RECT 195.675 -211.645 196.005 -211.315 ;
        RECT 195.675 -213.005 196.005 -212.675 ;
        RECT 195.675 -214.365 196.005 -214.035 ;
        RECT 195.675 -215.725 196.005 -215.395 ;
        RECT 195.675 -217.085 196.005 -216.755 ;
        RECT 195.675 -218.445 196.005 -218.115 ;
        RECT 195.675 -224.09 196.005 -222.96 ;
        RECT 195.68 -224.205 196 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.035 132.52 197.365 133.65 ;
        RECT 197.035 128.355 197.365 128.685 ;
        RECT 197.035 126.995 197.365 127.325 ;
        RECT 197.035 125.635 197.365 125.965 ;
        RECT 197.035 124.275 197.365 124.605 ;
        RECT 197.04 123.6 197.36 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.035 -0.845 197.365 -0.515 ;
        RECT 197.035 -2.205 197.365 -1.875 ;
        RECT 197.035 -3.565 197.365 -3.235 ;
        RECT 197.04 -3.565 197.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.035 -119.165 197.365 -118.835 ;
        RECT 197.035 -120.525 197.365 -120.195 ;
        RECT 197.035 -121.885 197.365 -121.555 ;
        RECT 197.035 -123.245 197.365 -122.915 ;
        RECT 197.035 -124.605 197.365 -124.275 ;
        RECT 197.035 -125.965 197.365 -125.635 ;
        RECT 197.035 -127.325 197.365 -126.995 ;
        RECT 197.035 -128.685 197.365 -128.355 ;
        RECT 197.035 -130.045 197.365 -129.715 ;
        RECT 197.035 -131.405 197.365 -131.075 ;
        RECT 197.035 -132.765 197.365 -132.435 ;
        RECT 197.035 -134.125 197.365 -133.795 ;
        RECT 197.035 -135.485 197.365 -135.155 ;
        RECT 197.035 -136.845 197.365 -136.515 ;
        RECT 197.035 -138.205 197.365 -137.875 ;
        RECT 197.035 -139.565 197.365 -139.235 ;
        RECT 197.035 -140.925 197.365 -140.595 ;
        RECT 197.035 -142.285 197.365 -141.955 ;
        RECT 197.035 -143.645 197.365 -143.315 ;
        RECT 197.035 -145.005 197.365 -144.675 ;
        RECT 197.035 -146.365 197.365 -146.035 ;
        RECT 197.035 -147.725 197.365 -147.395 ;
        RECT 197.035 -149.085 197.365 -148.755 ;
        RECT 197.035 -150.445 197.365 -150.115 ;
        RECT 197.035 -151.805 197.365 -151.475 ;
        RECT 197.035 -153.165 197.365 -152.835 ;
        RECT 197.035 -154.525 197.365 -154.195 ;
        RECT 197.035 -155.885 197.365 -155.555 ;
        RECT 197.035 -157.245 197.365 -156.915 ;
        RECT 197.035 -158.605 197.365 -158.275 ;
        RECT 197.035 -159.965 197.365 -159.635 ;
        RECT 197.035 -161.325 197.365 -160.995 ;
        RECT 197.035 -162.685 197.365 -162.355 ;
        RECT 197.035 -164.045 197.365 -163.715 ;
        RECT 197.035 -165.405 197.365 -165.075 ;
        RECT 197.035 -166.765 197.365 -166.435 ;
        RECT 197.035 -168.125 197.365 -167.795 ;
        RECT 197.035 -169.485 197.365 -169.155 ;
        RECT 197.035 -170.845 197.365 -170.515 ;
        RECT 197.035 -172.205 197.365 -171.875 ;
        RECT 197.035 -173.565 197.365 -173.235 ;
        RECT 197.035 -174.925 197.365 -174.595 ;
        RECT 197.035 -176.285 197.365 -175.955 ;
        RECT 197.035 -177.645 197.365 -177.315 ;
        RECT 197.035 -179.005 197.365 -178.675 ;
        RECT 197.035 -180.365 197.365 -180.035 ;
        RECT 197.035 -181.725 197.365 -181.395 ;
        RECT 197.035 -183.085 197.365 -182.755 ;
        RECT 197.035 -184.445 197.365 -184.115 ;
        RECT 197.035 -185.805 197.365 -185.475 ;
        RECT 197.035 -187.165 197.365 -186.835 ;
        RECT 197.035 -188.525 197.365 -188.195 ;
        RECT 197.035 -189.885 197.365 -189.555 ;
        RECT 197.035 -191.245 197.365 -190.915 ;
        RECT 197.035 -192.605 197.365 -192.275 ;
        RECT 197.035 -193.965 197.365 -193.635 ;
        RECT 197.035 -195.325 197.365 -194.995 ;
        RECT 197.035 -196.685 197.365 -196.355 ;
        RECT 197.035 -198.045 197.365 -197.715 ;
        RECT 197.035 -199.405 197.365 -199.075 ;
        RECT 197.035 -200.765 197.365 -200.435 ;
        RECT 197.035 -202.125 197.365 -201.795 ;
        RECT 197.035 -203.485 197.365 -203.155 ;
        RECT 197.035 -204.845 197.365 -204.515 ;
        RECT 197.035 -206.205 197.365 -205.875 ;
        RECT 197.035 -207.565 197.365 -207.235 ;
        RECT 197.035 -208.925 197.365 -208.595 ;
        RECT 197.035 -210.285 197.365 -209.955 ;
        RECT 197.035 -211.645 197.365 -211.315 ;
        RECT 197.035 -213.005 197.365 -212.675 ;
        RECT 197.035 -214.365 197.365 -214.035 ;
        RECT 197.035 -215.725 197.365 -215.395 ;
        RECT 197.035 -217.085 197.365 -216.755 ;
        RECT 197.035 -218.445 197.365 -218.115 ;
        RECT 197.035 -224.09 197.365 -222.96 ;
        RECT 197.04 -224.205 197.36 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.395 132.52 198.725 133.65 ;
        RECT 198.395 128.355 198.725 128.685 ;
        RECT 198.395 126.995 198.725 127.325 ;
        RECT 198.395 125.635 198.725 125.965 ;
        RECT 198.395 124.275 198.725 124.605 ;
        RECT 198.4 123.6 198.72 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.395 -123.245 198.725 -122.915 ;
        RECT 198.395 -124.605 198.725 -124.275 ;
        RECT 198.395 -125.965 198.725 -125.635 ;
        RECT 198.395 -127.325 198.725 -126.995 ;
        RECT 198.395 -128.685 198.725 -128.355 ;
        RECT 198.395 -130.045 198.725 -129.715 ;
        RECT 198.395 -131.405 198.725 -131.075 ;
        RECT 198.395 -132.765 198.725 -132.435 ;
        RECT 198.395 -134.125 198.725 -133.795 ;
        RECT 198.395 -135.485 198.725 -135.155 ;
        RECT 198.395 -136.845 198.725 -136.515 ;
        RECT 198.395 -138.205 198.725 -137.875 ;
        RECT 198.395 -139.565 198.725 -139.235 ;
        RECT 198.395 -140.925 198.725 -140.595 ;
        RECT 198.395 -142.285 198.725 -141.955 ;
        RECT 198.395 -143.645 198.725 -143.315 ;
        RECT 198.395 -145.005 198.725 -144.675 ;
        RECT 198.395 -146.365 198.725 -146.035 ;
        RECT 198.395 -147.725 198.725 -147.395 ;
        RECT 198.395 -149.085 198.725 -148.755 ;
        RECT 198.395 -150.445 198.725 -150.115 ;
        RECT 198.395 -151.805 198.725 -151.475 ;
        RECT 198.395 -153.165 198.725 -152.835 ;
        RECT 198.395 -154.525 198.725 -154.195 ;
        RECT 198.395 -155.885 198.725 -155.555 ;
        RECT 198.395 -157.245 198.725 -156.915 ;
        RECT 198.395 -158.605 198.725 -158.275 ;
        RECT 198.395 -159.965 198.725 -159.635 ;
        RECT 198.395 -161.325 198.725 -160.995 ;
        RECT 198.395 -162.685 198.725 -162.355 ;
        RECT 198.395 -164.045 198.725 -163.715 ;
        RECT 198.395 -165.405 198.725 -165.075 ;
        RECT 198.395 -166.765 198.725 -166.435 ;
        RECT 198.395 -168.125 198.725 -167.795 ;
        RECT 198.395 -169.485 198.725 -169.155 ;
        RECT 198.395 -170.845 198.725 -170.515 ;
        RECT 198.395 -172.205 198.725 -171.875 ;
        RECT 198.395 -173.565 198.725 -173.235 ;
        RECT 198.395 -174.925 198.725 -174.595 ;
        RECT 198.395 -176.285 198.725 -175.955 ;
        RECT 198.395 -177.645 198.725 -177.315 ;
        RECT 198.395 -179.005 198.725 -178.675 ;
        RECT 198.395 -180.365 198.725 -180.035 ;
        RECT 198.395 -181.725 198.725 -181.395 ;
        RECT 198.395 -183.085 198.725 -182.755 ;
        RECT 198.395 -184.445 198.725 -184.115 ;
        RECT 198.395 -185.805 198.725 -185.475 ;
        RECT 198.395 -187.165 198.725 -186.835 ;
        RECT 198.395 -188.525 198.725 -188.195 ;
        RECT 198.395 -189.885 198.725 -189.555 ;
        RECT 198.395 -191.245 198.725 -190.915 ;
        RECT 198.395 -192.605 198.725 -192.275 ;
        RECT 198.395 -193.965 198.725 -193.635 ;
        RECT 198.395 -195.325 198.725 -194.995 ;
        RECT 198.395 -196.685 198.725 -196.355 ;
        RECT 198.395 -198.045 198.725 -197.715 ;
        RECT 198.395 -199.405 198.725 -199.075 ;
        RECT 198.395 -200.765 198.725 -200.435 ;
        RECT 198.395 -202.125 198.725 -201.795 ;
        RECT 198.395 -203.485 198.725 -203.155 ;
        RECT 198.395 -204.845 198.725 -204.515 ;
        RECT 198.395 -206.205 198.725 -205.875 ;
        RECT 198.395 -207.565 198.725 -207.235 ;
        RECT 198.395 -208.925 198.725 -208.595 ;
        RECT 198.395 -210.285 198.725 -209.955 ;
        RECT 198.395 -211.645 198.725 -211.315 ;
        RECT 198.395 -213.005 198.725 -212.675 ;
        RECT 198.395 -214.365 198.725 -214.035 ;
        RECT 198.395 -215.725 198.725 -215.395 ;
        RECT 198.395 -217.085 198.725 -216.755 ;
        RECT 198.395 -218.445 198.725 -218.115 ;
        RECT 198.395 -224.09 198.725 -222.96 ;
        RECT 198.4 -224.205 198.72 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.51 -121.535 198.84 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.755 132.52 200.085 133.65 ;
        RECT 199.755 128.355 200.085 128.685 ;
        RECT 199.755 126.995 200.085 127.325 ;
        RECT 199.755 125.635 200.085 125.965 ;
        RECT 199.755 124.275 200.085 124.605 ;
        RECT 199.76 123.6 200.08 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.755 -0.845 200.085 -0.515 ;
        RECT 199.755 -2.205 200.085 -1.875 ;
        RECT 199.755 -3.565 200.085 -3.235 ;
        RECT 199.76 -3.565 200.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.755 -119.165 200.085 -118.835 ;
        RECT 199.755 -120.525 200.085 -120.195 ;
        RECT 199.755 -121.885 200.085 -121.555 ;
        RECT 199.755 -123.245 200.085 -122.915 ;
        RECT 199.755 -124.605 200.085 -124.275 ;
        RECT 199.755 -125.965 200.085 -125.635 ;
        RECT 199.755 -127.325 200.085 -126.995 ;
        RECT 199.755 -128.685 200.085 -128.355 ;
        RECT 199.755 -130.045 200.085 -129.715 ;
        RECT 199.755 -131.405 200.085 -131.075 ;
        RECT 199.755 -132.765 200.085 -132.435 ;
        RECT 199.755 -134.125 200.085 -133.795 ;
        RECT 199.755 -135.485 200.085 -135.155 ;
        RECT 199.755 -136.845 200.085 -136.515 ;
        RECT 199.755 -138.205 200.085 -137.875 ;
        RECT 199.755 -139.565 200.085 -139.235 ;
        RECT 199.755 -140.925 200.085 -140.595 ;
        RECT 199.755 -142.285 200.085 -141.955 ;
        RECT 199.755 -143.645 200.085 -143.315 ;
        RECT 199.755 -145.005 200.085 -144.675 ;
        RECT 199.755 -146.365 200.085 -146.035 ;
        RECT 199.755 -147.725 200.085 -147.395 ;
        RECT 199.755 -149.085 200.085 -148.755 ;
        RECT 199.755 -150.445 200.085 -150.115 ;
        RECT 199.755 -151.805 200.085 -151.475 ;
        RECT 199.755 -153.165 200.085 -152.835 ;
        RECT 199.755 -154.525 200.085 -154.195 ;
        RECT 199.755 -155.885 200.085 -155.555 ;
        RECT 199.755 -157.245 200.085 -156.915 ;
        RECT 199.755 -158.605 200.085 -158.275 ;
        RECT 199.755 -159.965 200.085 -159.635 ;
        RECT 199.755 -161.325 200.085 -160.995 ;
        RECT 199.755 -162.685 200.085 -162.355 ;
        RECT 199.755 -164.045 200.085 -163.715 ;
        RECT 199.755 -165.405 200.085 -165.075 ;
        RECT 199.755 -166.765 200.085 -166.435 ;
        RECT 199.755 -168.125 200.085 -167.795 ;
        RECT 199.755 -169.485 200.085 -169.155 ;
        RECT 199.755 -170.845 200.085 -170.515 ;
        RECT 199.755 -172.205 200.085 -171.875 ;
        RECT 199.755 -173.565 200.085 -173.235 ;
        RECT 199.755 -174.925 200.085 -174.595 ;
        RECT 199.755 -176.285 200.085 -175.955 ;
        RECT 199.755 -177.645 200.085 -177.315 ;
        RECT 199.755 -179.005 200.085 -178.675 ;
        RECT 199.755 -180.365 200.085 -180.035 ;
        RECT 199.755 -181.725 200.085 -181.395 ;
        RECT 199.755 -183.085 200.085 -182.755 ;
        RECT 199.755 -184.445 200.085 -184.115 ;
        RECT 199.755 -185.805 200.085 -185.475 ;
        RECT 199.755 -187.165 200.085 -186.835 ;
        RECT 199.755 -188.525 200.085 -188.195 ;
        RECT 199.755 -189.885 200.085 -189.555 ;
        RECT 199.755 -191.245 200.085 -190.915 ;
        RECT 199.755 -192.605 200.085 -192.275 ;
        RECT 199.755 -193.965 200.085 -193.635 ;
        RECT 199.755 -195.325 200.085 -194.995 ;
        RECT 199.755 -196.685 200.085 -196.355 ;
        RECT 199.755 -198.045 200.085 -197.715 ;
        RECT 199.755 -199.405 200.085 -199.075 ;
        RECT 199.755 -200.765 200.085 -200.435 ;
        RECT 199.755 -202.125 200.085 -201.795 ;
        RECT 199.755 -203.485 200.085 -203.155 ;
        RECT 199.755 -204.845 200.085 -204.515 ;
        RECT 199.755 -206.205 200.085 -205.875 ;
        RECT 199.755 -207.565 200.085 -207.235 ;
        RECT 199.755 -208.925 200.085 -208.595 ;
        RECT 199.755 -210.285 200.085 -209.955 ;
        RECT 199.755 -211.645 200.085 -211.315 ;
        RECT 199.755 -213.005 200.085 -212.675 ;
        RECT 199.755 -214.365 200.085 -214.035 ;
        RECT 199.755 -215.725 200.085 -215.395 ;
        RECT 199.755 -217.085 200.085 -216.755 ;
        RECT 199.755 -218.445 200.085 -218.115 ;
        RECT 199.755 -224.09 200.085 -222.96 ;
        RECT 199.76 -224.205 200.08 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.115 132.52 201.445 133.65 ;
        RECT 201.115 128.355 201.445 128.685 ;
        RECT 201.115 126.995 201.445 127.325 ;
        RECT 201.115 125.635 201.445 125.965 ;
        RECT 201.115 124.275 201.445 124.605 ;
        RECT 201.12 123.6 201.44 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.115 -0.845 201.445 -0.515 ;
        RECT 201.115 -2.205 201.445 -1.875 ;
        RECT 201.115 -3.565 201.445 -3.235 ;
        RECT 201.12 -3.565 201.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.115 -119.165 201.445 -118.835 ;
        RECT 201.115 -120.525 201.445 -120.195 ;
        RECT 201.115 -121.885 201.445 -121.555 ;
        RECT 201.115 -123.245 201.445 -122.915 ;
        RECT 201.115 -124.605 201.445 -124.275 ;
        RECT 201.115 -125.965 201.445 -125.635 ;
        RECT 201.115 -127.325 201.445 -126.995 ;
        RECT 201.115 -128.685 201.445 -128.355 ;
        RECT 201.115 -130.045 201.445 -129.715 ;
        RECT 201.115 -131.405 201.445 -131.075 ;
        RECT 201.115 -132.765 201.445 -132.435 ;
        RECT 201.115 -134.125 201.445 -133.795 ;
        RECT 201.115 -135.485 201.445 -135.155 ;
        RECT 201.115 -136.845 201.445 -136.515 ;
        RECT 201.115 -138.205 201.445 -137.875 ;
        RECT 201.115 -139.565 201.445 -139.235 ;
        RECT 201.115 -140.925 201.445 -140.595 ;
        RECT 201.115 -142.285 201.445 -141.955 ;
        RECT 201.115 -143.645 201.445 -143.315 ;
        RECT 201.115 -145.005 201.445 -144.675 ;
        RECT 201.115 -146.365 201.445 -146.035 ;
        RECT 201.115 -147.725 201.445 -147.395 ;
        RECT 201.115 -149.085 201.445 -148.755 ;
        RECT 201.115 -150.445 201.445 -150.115 ;
        RECT 201.115 -151.805 201.445 -151.475 ;
        RECT 201.115 -153.165 201.445 -152.835 ;
        RECT 201.115 -154.525 201.445 -154.195 ;
        RECT 201.115 -155.885 201.445 -155.555 ;
        RECT 201.115 -157.245 201.445 -156.915 ;
        RECT 201.115 -158.605 201.445 -158.275 ;
        RECT 201.115 -159.965 201.445 -159.635 ;
        RECT 201.115 -161.325 201.445 -160.995 ;
        RECT 201.115 -162.685 201.445 -162.355 ;
        RECT 201.115 -164.045 201.445 -163.715 ;
        RECT 201.115 -165.405 201.445 -165.075 ;
        RECT 201.115 -166.765 201.445 -166.435 ;
        RECT 201.115 -168.125 201.445 -167.795 ;
        RECT 201.115 -169.485 201.445 -169.155 ;
        RECT 201.115 -170.845 201.445 -170.515 ;
        RECT 201.115 -172.205 201.445 -171.875 ;
        RECT 201.115 -173.565 201.445 -173.235 ;
        RECT 201.115 -174.925 201.445 -174.595 ;
        RECT 201.115 -176.285 201.445 -175.955 ;
        RECT 201.115 -177.645 201.445 -177.315 ;
        RECT 201.115 -179.005 201.445 -178.675 ;
        RECT 201.115 -180.365 201.445 -180.035 ;
        RECT 201.115 -181.725 201.445 -181.395 ;
        RECT 201.115 -183.085 201.445 -182.755 ;
        RECT 201.115 -184.445 201.445 -184.115 ;
        RECT 201.115 -185.805 201.445 -185.475 ;
        RECT 201.115 -187.165 201.445 -186.835 ;
        RECT 201.115 -188.525 201.445 -188.195 ;
        RECT 201.115 -189.885 201.445 -189.555 ;
        RECT 201.115 -191.245 201.445 -190.915 ;
        RECT 201.115 -192.605 201.445 -192.275 ;
        RECT 201.115 -193.965 201.445 -193.635 ;
        RECT 201.115 -195.325 201.445 -194.995 ;
        RECT 201.115 -196.685 201.445 -196.355 ;
        RECT 201.115 -198.045 201.445 -197.715 ;
        RECT 201.115 -199.405 201.445 -199.075 ;
        RECT 201.115 -200.765 201.445 -200.435 ;
        RECT 201.115 -202.125 201.445 -201.795 ;
        RECT 201.115 -203.485 201.445 -203.155 ;
        RECT 201.115 -204.845 201.445 -204.515 ;
        RECT 201.115 -206.205 201.445 -205.875 ;
        RECT 201.115 -207.565 201.445 -207.235 ;
        RECT 201.115 -208.925 201.445 -208.595 ;
        RECT 201.115 -210.285 201.445 -209.955 ;
        RECT 201.115 -211.645 201.445 -211.315 ;
        RECT 201.115 -213.005 201.445 -212.675 ;
        RECT 201.115 -214.365 201.445 -214.035 ;
        RECT 201.115 -215.725 201.445 -215.395 ;
        RECT 201.115 -217.085 201.445 -216.755 ;
        RECT 201.115 -218.445 201.445 -218.115 ;
        RECT 201.115 -224.09 201.445 -222.96 ;
        RECT 201.12 -224.205 201.44 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 202.475 132.52 202.805 133.65 ;
        RECT 202.475 128.355 202.805 128.685 ;
        RECT 202.475 126.995 202.805 127.325 ;
        RECT 202.475 125.635 202.805 125.965 ;
        RECT 202.475 124.275 202.805 124.605 ;
        RECT 202.475 121.41 202.805 121.74 ;
        RECT 202.475 119.235 202.805 119.565 ;
        RECT 202.475 117.655 202.805 117.985 ;
        RECT 202.475 116.805 202.805 117.135 ;
        RECT 202.475 114.495 202.805 114.825 ;
        RECT 202.475 113.645 202.805 113.975 ;
        RECT 202.475 111.335 202.805 111.665 ;
        RECT 202.475 110.485 202.805 110.815 ;
        RECT 202.475 108.175 202.805 108.505 ;
        RECT 202.475 107.325 202.805 107.655 ;
        RECT 202.475 105.015 202.805 105.345 ;
        RECT 202.475 103.435 202.805 103.765 ;
        RECT 202.475 102.585 202.805 102.915 ;
        RECT 202.475 100.275 202.805 100.605 ;
        RECT 202.475 99.425 202.805 99.755 ;
        RECT 202.475 97.115 202.805 97.445 ;
        RECT 202.475 96.265 202.805 96.595 ;
        RECT 202.475 93.955 202.805 94.285 ;
        RECT 202.475 93.105 202.805 93.435 ;
        RECT 202.475 90.795 202.805 91.125 ;
        RECT 202.475 89.215 202.805 89.545 ;
        RECT 202.475 88.365 202.805 88.695 ;
        RECT 202.475 86.055 202.805 86.385 ;
        RECT 202.475 85.205 202.805 85.535 ;
        RECT 202.475 82.895 202.805 83.225 ;
        RECT 202.475 82.045 202.805 82.375 ;
        RECT 202.475 79.735 202.805 80.065 ;
        RECT 202.475 78.885 202.805 79.215 ;
        RECT 202.475 76.575 202.805 76.905 ;
        RECT 202.475 74.995 202.805 75.325 ;
        RECT 202.475 74.145 202.805 74.475 ;
        RECT 202.475 71.835 202.805 72.165 ;
        RECT 202.475 70.985 202.805 71.315 ;
        RECT 202.475 68.675 202.805 69.005 ;
        RECT 202.475 67.825 202.805 68.155 ;
        RECT 202.475 65.515 202.805 65.845 ;
        RECT 202.475 64.665 202.805 64.995 ;
        RECT 202.475 62.355 202.805 62.685 ;
        RECT 202.475 60.775 202.805 61.105 ;
        RECT 202.475 59.925 202.805 60.255 ;
        RECT 202.475 57.615 202.805 57.945 ;
        RECT 202.475 56.765 202.805 57.095 ;
        RECT 202.475 54.455 202.805 54.785 ;
        RECT 202.475 53.605 202.805 53.935 ;
        RECT 202.475 51.295 202.805 51.625 ;
        RECT 202.475 50.445 202.805 50.775 ;
        RECT 202.475 48.135 202.805 48.465 ;
        RECT 202.475 46.555 202.805 46.885 ;
        RECT 202.475 45.705 202.805 46.035 ;
        RECT 202.475 43.395 202.805 43.725 ;
        RECT 202.475 42.545 202.805 42.875 ;
        RECT 202.475 40.235 202.805 40.565 ;
        RECT 202.475 39.385 202.805 39.715 ;
        RECT 202.475 37.075 202.805 37.405 ;
        RECT 202.475 36.225 202.805 36.555 ;
        RECT 202.475 33.915 202.805 34.245 ;
        RECT 202.475 32.335 202.805 32.665 ;
        RECT 202.475 31.485 202.805 31.815 ;
        RECT 202.475 29.175 202.805 29.505 ;
        RECT 202.475 28.325 202.805 28.655 ;
        RECT 202.475 26.015 202.805 26.345 ;
        RECT 202.475 25.165 202.805 25.495 ;
        RECT 202.475 22.855 202.805 23.185 ;
        RECT 202.475 22.005 202.805 22.335 ;
        RECT 202.475 19.695 202.805 20.025 ;
        RECT 202.475 18.115 202.805 18.445 ;
        RECT 202.475 17.265 202.805 17.595 ;
        RECT 202.475 14.955 202.805 15.285 ;
        RECT 202.475 14.105 202.805 14.435 ;
        RECT 202.475 11.795 202.805 12.125 ;
        RECT 202.475 10.945 202.805 11.275 ;
        RECT 202.475 8.635 202.805 8.965 ;
        RECT 202.475 7.785 202.805 8.115 ;
        RECT 202.475 5.475 202.805 5.805 ;
        RECT 202.475 3.895 202.805 4.225 ;
        RECT 202.475 3.045 202.805 3.375 ;
        RECT 202.475 0.87 202.805 1.2 ;
        RECT 202.475 -0.845 202.805 -0.515 ;
        RECT 202.475 -2.205 202.805 -1.875 ;
        RECT 202.475 -3.565 202.805 -3.235 ;
        RECT 202.475 -4.925 202.805 -4.595 ;
        RECT 202.475 -6.285 202.805 -5.955 ;
        RECT 202.475 -7.645 202.805 -7.315 ;
        RECT 202.475 -9.005 202.805 -8.675 ;
        RECT 202.475 -10.365 202.805 -10.035 ;
        RECT 202.475 -11.725 202.805 -11.395 ;
        RECT 202.475 -13.085 202.805 -12.755 ;
        RECT 202.475 -14.445 202.805 -14.115 ;
        RECT 202.475 -15.805 202.805 -15.475 ;
        RECT 202.475 -17.165 202.805 -16.835 ;
        RECT 202.475 -18.525 202.805 -18.195 ;
        RECT 202.475 -19.885 202.805 -19.555 ;
        RECT 202.475 -21.245 202.805 -20.915 ;
        RECT 202.475 -22.605 202.805 -22.275 ;
        RECT 202.475 -23.965 202.805 -23.635 ;
        RECT 202.475 -25.325 202.805 -24.995 ;
        RECT 202.475 -26.685 202.805 -26.355 ;
        RECT 202.475 -28.045 202.805 -27.715 ;
        RECT 202.475 -29.405 202.805 -29.075 ;
        RECT 202.475 -30.765 202.805 -30.435 ;
        RECT 202.475 -32.125 202.805 -31.795 ;
        RECT 202.475 -33.485 202.805 -33.155 ;
        RECT 202.475 -34.845 202.805 -34.515 ;
        RECT 202.475 -36.205 202.805 -35.875 ;
        RECT 202.475 -37.565 202.805 -37.235 ;
        RECT 202.475 -38.925 202.805 -38.595 ;
        RECT 202.475 -40.285 202.805 -39.955 ;
        RECT 202.475 -41.645 202.805 -41.315 ;
        RECT 202.475 -43.005 202.805 -42.675 ;
        RECT 202.475 -44.365 202.805 -44.035 ;
        RECT 202.475 -45.725 202.805 -45.395 ;
        RECT 202.475 -47.085 202.805 -46.755 ;
        RECT 202.475 -48.445 202.805 -48.115 ;
        RECT 202.475 -49.805 202.805 -49.475 ;
        RECT 202.475 -51.165 202.805 -50.835 ;
        RECT 202.475 -52.525 202.805 -52.195 ;
        RECT 202.475 -53.885 202.805 -53.555 ;
        RECT 202.475 -55.245 202.805 -54.915 ;
        RECT 202.475 -56.605 202.805 -56.275 ;
        RECT 202.475 -57.965 202.805 -57.635 ;
        RECT 202.475 -59.325 202.805 -58.995 ;
        RECT 202.475 -60.685 202.805 -60.355 ;
        RECT 202.475 -62.045 202.805 -61.715 ;
        RECT 202.475 -63.405 202.805 -63.075 ;
        RECT 202.475 -64.765 202.805 -64.435 ;
        RECT 202.475 -66.125 202.805 -65.795 ;
        RECT 202.475 -67.485 202.805 -67.155 ;
        RECT 202.475 -68.845 202.805 -68.515 ;
        RECT 202.475 -70.205 202.805 -69.875 ;
        RECT 202.475 -71.565 202.805 -71.235 ;
        RECT 202.475 -72.925 202.805 -72.595 ;
        RECT 202.475 -74.285 202.805 -73.955 ;
        RECT 202.475 -75.645 202.805 -75.315 ;
        RECT 202.475 -77.005 202.805 -76.675 ;
        RECT 202.475 -78.365 202.805 -78.035 ;
        RECT 202.475 -79.725 202.805 -79.395 ;
        RECT 202.475 -81.085 202.805 -80.755 ;
        RECT 202.475 -82.445 202.805 -82.115 ;
        RECT 202.475 -83.805 202.805 -83.475 ;
        RECT 202.475 -85.165 202.805 -84.835 ;
        RECT 202.475 -86.525 202.805 -86.195 ;
        RECT 202.475 -87.885 202.805 -87.555 ;
        RECT 202.475 -89.245 202.805 -88.915 ;
        RECT 202.475 -90.605 202.805 -90.275 ;
        RECT 202.475 -91.965 202.805 -91.635 ;
        RECT 202.475 -93.325 202.805 -92.995 ;
        RECT 202.475 -94.685 202.805 -94.355 ;
        RECT 202.475 -96.045 202.805 -95.715 ;
        RECT 202.475 -97.405 202.805 -97.075 ;
        RECT 202.475 -98.765 202.805 -98.435 ;
        RECT 202.475 -100.125 202.805 -99.795 ;
        RECT 202.475 -101.485 202.805 -101.155 ;
        RECT 202.475 -102.845 202.805 -102.515 ;
        RECT 202.475 -104.205 202.805 -103.875 ;
        RECT 202.475 -105.565 202.805 -105.235 ;
        RECT 202.475 -106.925 202.805 -106.595 ;
        RECT 202.475 -108.285 202.805 -107.955 ;
        RECT 202.475 -109.645 202.805 -109.315 ;
        RECT 202.475 -111.005 202.805 -110.675 ;
        RECT 202.475 -112.365 202.805 -112.035 ;
        RECT 202.475 -113.725 202.805 -113.395 ;
        RECT 202.475 -115.085 202.805 -114.755 ;
        RECT 202.475 -116.445 202.805 -116.115 ;
        RECT 202.475 -117.805 202.805 -117.475 ;
        RECT 202.475 -119.165 202.805 -118.835 ;
        RECT 202.475 -120.525 202.805 -120.195 ;
        RECT 202.475 -121.885 202.805 -121.555 ;
        RECT 202.475 -123.245 202.805 -122.915 ;
        RECT 202.475 -124.605 202.805 -124.275 ;
        RECT 202.475 -125.965 202.805 -125.635 ;
        RECT 202.475 -127.325 202.805 -126.995 ;
        RECT 202.475 -128.685 202.805 -128.355 ;
        RECT 202.475 -130.045 202.805 -129.715 ;
        RECT 202.475 -131.405 202.805 -131.075 ;
        RECT 202.475 -132.765 202.805 -132.435 ;
        RECT 202.475 -134.125 202.805 -133.795 ;
        RECT 202.475 -135.485 202.805 -135.155 ;
        RECT 202.475 -136.845 202.805 -136.515 ;
        RECT 202.475 -138.205 202.805 -137.875 ;
        RECT 202.475 -139.565 202.805 -139.235 ;
        RECT 202.475 -140.925 202.805 -140.595 ;
        RECT 202.475 -142.285 202.805 -141.955 ;
        RECT 202.475 -143.645 202.805 -143.315 ;
        RECT 202.475 -145.005 202.805 -144.675 ;
        RECT 202.475 -146.365 202.805 -146.035 ;
        RECT 202.475 -147.725 202.805 -147.395 ;
        RECT 202.475 -149.085 202.805 -148.755 ;
        RECT 202.475 -150.445 202.805 -150.115 ;
        RECT 202.475 -151.805 202.805 -151.475 ;
        RECT 202.475 -153.165 202.805 -152.835 ;
        RECT 202.475 -154.525 202.805 -154.195 ;
        RECT 202.475 -155.885 202.805 -155.555 ;
        RECT 202.475 -157.245 202.805 -156.915 ;
        RECT 202.475 -158.605 202.805 -158.275 ;
        RECT 202.475 -159.965 202.805 -159.635 ;
        RECT 202.475 -161.325 202.805 -160.995 ;
        RECT 202.475 -162.685 202.805 -162.355 ;
        RECT 202.475 -164.045 202.805 -163.715 ;
        RECT 202.475 -165.405 202.805 -165.075 ;
        RECT 202.475 -166.765 202.805 -166.435 ;
        RECT 202.475 -168.125 202.805 -167.795 ;
        RECT 202.475 -169.485 202.805 -169.155 ;
        RECT 202.475 -170.845 202.805 -170.515 ;
        RECT 202.475 -172.205 202.805 -171.875 ;
        RECT 202.475 -173.565 202.805 -173.235 ;
        RECT 202.475 -174.925 202.805 -174.595 ;
        RECT 202.475 -176.285 202.805 -175.955 ;
        RECT 202.475 -177.645 202.805 -177.315 ;
        RECT 202.475 -179.005 202.805 -178.675 ;
        RECT 202.475 -180.365 202.805 -180.035 ;
        RECT 202.475 -181.725 202.805 -181.395 ;
        RECT 202.475 -183.085 202.805 -182.755 ;
        RECT 202.475 -184.445 202.805 -184.115 ;
        RECT 202.475 -185.805 202.805 -185.475 ;
        RECT 202.475 -187.165 202.805 -186.835 ;
        RECT 202.475 -188.525 202.805 -188.195 ;
        RECT 202.475 -189.885 202.805 -189.555 ;
        RECT 202.475 -191.245 202.805 -190.915 ;
        RECT 202.475 -192.605 202.805 -192.275 ;
        RECT 202.475 -193.965 202.805 -193.635 ;
        RECT 202.475 -195.325 202.805 -194.995 ;
        RECT 202.475 -196.685 202.805 -196.355 ;
        RECT 202.475 -198.045 202.805 -197.715 ;
        RECT 202.475 -199.405 202.805 -199.075 ;
        RECT 202.475 -200.765 202.805 -200.435 ;
        RECT 202.475 -202.125 202.805 -201.795 ;
        RECT 202.475 -203.485 202.805 -203.155 ;
        RECT 202.475 -204.845 202.805 -204.515 ;
        RECT 202.475 -206.205 202.805 -205.875 ;
        RECT 202.475 -207.565 202.805 -207.235 ;
        RECT 202.475 -208.925 202.805 -208.595 ;
        RECT 202.475 -210.285 202.805 -209.955 ;
        RECT 202.475 -211.645 202.805 -211.315 ;
        RECT 202.475 -213.005 202.805 -212.675 ;
        RECT 202.475 -214.365 202.805 -214.035 ;
        RECT 202.475 -215.725 202.805 -215.395 ;
        RECT 202.475 -217.085 202.805 -216.755 ;
        RECT 202.475 -218.445 202.805 -218.115 ;
        RECT 202.475 -224.09 202.805 -222.96 ;
        RECT 202.48 -224.205 202.8 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.835 132.52 204.165 133.65 ;
        RECT 203.835 128.355 204.165 128.685 ;
        RECT 203.835 126.995 204.165 127.325 ;
        RECT 203.835 125.635 204.165 125.965 ;
        RECT 203.835 124.275 204.165 124.605 ;
        RECT 203.835 121.41 204.165 121.74 ;
        RECT 203.835 119.235 204.165 119.565 ;
        RECT 203.835 117.655 204.165 117.985 ;
        RECT 203.835 116.805 204.165 117.135 ;
        RECT 203.835 114.495 204.165 114.825 ;
        RECT 203.835 113.645 204.165 113.975 ;
        RECT 203.835 111.335 204.165 111.665 ;
        RECT 203.835 110.485 204.165 110.815 ;
        RECT 203.835 108.175 204.165 108.505 ;
        RECT 203.835 107.325 204.165 107.655 ;
        RECT 203.835 105.015 204.165 105.345 ;
        RECT 203.835 103.435 204.165 103.765 ;
        RECT 203.835 102.585 204.165 102.915 ;
        RECT 203.835 100.275 204.165 100.605 ;
        RECT 203.835 99.425 204.165 99.755 ;
        RECT 203.835 97.115 204.165 97.445 ;
        RECT 203.835 96.265 204.165 96.595 ;
        RECT 203.835 93.955 204.165 94.285 ;
        RECT 203.835 93.105 204.165 93.435 ;
        RECT 203.835 90.795 204.165 91.125 ;
        RECT 203.835 89.215 204.165 89.545 ;
        RECT 203.835 88.365 204.165 88.695 ;
        RECT 203.835 86.055 204.165 86.385 ;
        RECT 203.835 85.205 204.165 85.535 ;
        RECT 203.835 82.895 204.165 83.225 ;
        RECT 203.835 82.045 204.165 82.375 ;
        RECT 203.835 79.735 204.165 80.065 ;
        RECT 203.835 78.885 204.165 79.215 ;
        RECT 203.835 76.575 204.165 76.905 ;
        RECT 203.835 74.995 204.165 75.325 ;
        RECT 203.835 74.145 204.165 74.475 ;
        RECT 203.835 71.835 204.165 72.165 ;
        RECT 203.835 70.985 204.165 71.315 ;
        RECT 203.835 68.675 204.165 69.005 ;
        RECT 203.835 67.825 204.165 68.155 ;
        RECT 203.835 65.515 204.165 65.845 ;
        RECT 203.835 64.665 204.165 64.995 ;
        RECT 203.835 62.355 204.165 62.685 ;
        RECT 203.835 60.775 204.165 61.105 ;
        RECT 203.835 59.925 204.165 60.255 ;
        RECT 203.835 57.615 204.165 57.945 ;
        RECT 203.835 56.765 204.165 57.095 ;
        RECT 203.835 54.455 204.165 54.785 ;
        RECT 203.835 53.605 204.165 53.935 ;
        RECT 203.835 51.295 204.165 51.625 ;
        RECT 203.835 50.445 204.165 50.775 ;
        RECT 203.835 48.135 204.165 48.465 ;
        RECT 203.835 46.555 204.165 46.885 ;
        RECT 203.835 45.705 204.165 46.035 ;
        RECT 203.835 43.395 204.165 43.725 ;
        RECT 203.835 42.545 204.165 42.875 ;
        RECT 203.835 40.235 204.165 40.565 ;
        RECT 203.835 39.385 204.165 39.715 ;
        RECT 203.835 37.075 204.165 37.405 ;
        RECT 203.835 36.225 204.165 36.555 ;
        RECT 203.835 33.915 204.165 34.245 ;
        RECT 203.835 32.335 204.165 32.665 ;
        RECT 203.835 31.485 204.165 31.815 ;
        RECT 203.835 29.175 204.165 29.505 ;
        RECT 203.835 28.325 204.165 28.655 ;
        RECT 203.835 26.015 204.165 26.345 ;
        RECT 203.835 25.165 204.165 25.495 ;
        RECT 203.835 22.855 204.165 23.185 ;
        RECT 203.835 22.005 204.165 22.335 ;
        RECT 203.835 19.695 204.165 20.025 ;
        RECT 203.835 18.115 204.165 18.445 ;
        RECT 203.835 17.265 204.165 17.595 ;
        RECT 203.835 14.955 204.165 15.285 ;
        RECT 203.835 14.105 204.165 14.435 ;
        RECT 203.835 11.795 204.165 12.125 ;
        RECT 203.835 10.945 204.165 11.275 ;
        RECT 203.835 8.635 204.165 8.965 ;
        RECT 203.835 7.785 204.165 8.115 ;
        RECT 203.835 5.475 204.165 5.805 ;
        RECT 203.835 3.895 204.165 4.225 ;
        RECT 203.835 3.045 204.165 3.375 ;
        RECT 203.835 0.87 204.165 1.2 ;
        RECT 203.835 -0.845 204.165 -0.515 ;
        RECT 203.835 -2.205 204.165 -1.875 ;
        RECT 203.835 -3.565 204.165 -3.235 ;
        RECT 203.835 -4.925 204.165 -4.595 ;
        RECT 203.835 -6.285 204.165 -5.955 ;
        RECT 203.835 -7.645 204.165 -7.315 ;
        RECT 203.835 -9.005 204.165 -8.675 ;
        RECT 203.835 -10.365 204.165 -10.035 ;
        RECT 203.835 -11.725 204.165 -11.395 ;
        RECT 203.835 -13.085 204.165 -12.755 ;
        RECT 203.835 -14.445 204.165 -14.115 ;
        RECT 203.835 -15.805 204.165 -15.475 ;
        RECT 203.835 -17.165 204.165 -16.835 ;
        RECT 203.835 -18.525 204.165 -18.195 ;
        RECT 203.835 -19.885 204.165 -19.555 ;
        RECT 203.835 -21.245 204.165 -20.915 ;
        RECT 203.835 -22.605 204.165 -22.275 ;
        RECT 203.835 -23.965 204.165 -23.635 ;
        RECT 203.835 -25.325 204.165 -24.995 ;
        RECT 203.835 -26.685 204.165 -26.355 ;
        RECT 203.835 -28.045 204.165 -27.715 ;
        RECT 203.835 -29.405 204.165 -29.075 ;
        RECT 203.835 -30.765 204.165 -30.435 ;
        RECT 203.835 -32.125 204.165 -31.795 ;
        RECT 203.835 -33.485 204.165 -33.155 ;
        RECT 203.835 -34.845 204.165 -34.515 ;
        RECT 203.835 -36.205 204.165 -35.875 ;
        RECT 203.835 -37.565 204.165 -37.235 ;
        RECT 203.835 -38.925 204.165 -38.595 ;
        RECT 203.835 -40.285 204.165 -39.955 ;
        RECT 203.835 -41.645 204.165 -41.315 ;
        RECT 203.835 -43.005 204.165 -42.675 ;
        RECT 203.835 -44.365 204.165 -44.035 ;
        RECT 203.835 -45.725 204.165 -45.395 ;
        RECT 203.835 -47.085 204.165 -46.755 ;
        RECT 203.835 -48.445 204.165 -48.115 ;
        RECT 203.835 -49.805 204.165 -49.475 ;
        RECT 203.835 -51.165 204.165 -50.835 ;
        RECT 203.835 -52.525 204.165 -52.195 ;
        RECT 203.835 -53.885 204.165 -53.555 ;
        RECT 203.835 -55.245 204.165 -54.915 ;
        RECT 203.835 -56.605 204.165 -56.275 ;
        RECT 203.835 -57.965 204.165 -57.635 ;
        RECT 203.835 -59.325 204.165 -58.995 ;
        RECT 203.835 -60.685 204.165 -60.355 ;
        RECT 203.835 -62.045 204.165 -61.715 ;
        RECT 203.835 -63.405 204.165 -63.075 ;
        RECT 203.835 -64.765 204.165 -64.435 ;
        RECT 203.835 -66.125 204.165 -65.795 ;
        RECT 203.835 -67.485 204.165 -67.155 ;
        RECT 203.835 -68.845 204.165 -68.515 ;
        RECT 203.835 -70.205 204.165 -69.875 ;
        RECT 203.835 -71.565 204.165 -71.235 ;
        RECT 203.835 -72.925 204.165 -72.595 ;
        RECT 203.835 -74.285 204.165 -73.955 ;
        RECT 203.835 -75.645 204.165 -75.315 ;
        RECT 203.835 -77.005 204.165 -76.675 ;
        RECT 203.835 -78.365 204.165 -78.035 ;
        RECT 203.835 -79.725 204.165 -79.395 ;
        RECT 203.835 -81.085 204.165 -80.755 ;
        RECT 203.835 -82.445 204.165 -82.115 ;
        RECT 203.835 -83.805 204.165 -83.475 ;
        RECT 203.835 -85.165 204.165 -84.835 ;
        RECT 203.835 -86.525 204.165 -86.195 ;
        RECT 203.835 -87.885 204.165 -87.555 ;
        RECT 203.835 -89.245 204.165 -88.915 ;
        RECT 203.835 -90.605 204.165 -90.275 ;
        RECT 203.835 -91.965 204.165 -91.635 ;
        RECT 203.835 -93.325 204.165 -92.995 ;
        RECT 203.835 -94.685 204.165 -94.355 ;
        RECT 203.835 -96.045 204.165 -95.715 ;
        RECT 203.835 -97.405 204.165 -97.075 ;
        RECT 203.835 -98.765 204.165 -98.435 ;
        RECT 203.835 -100.125 204.165 -99.795 ;
        RECT 203.835 -101.485 204.165 -101.155 ;
        RECT 203.835 -102.845 204.165 -102.515 ;
        RECT 203.835 -104.205 204.165 -103.875 ;
        RECT 203.835 -105.565 204.165 -105.235 ;
        RECT 203.835 -106.925 204.165 -106.595 ;
        RECT 203.835 -108.285 204.165 -107.955 ;
        RECT 203.835 -109.645 204.165 -109.315 ;
        RECT 203.835 -111.005 204.165 -110.675 ;
        RECT 203.835 -112.365 204.165 -112.035 ;
        RECT 203.835 -113.725 204.165 -113.395 ;
        RECT 203.835 -115.085 204.165 -114.755 ;
        RECT 203.835 -116.445 204.165 -116.115 ;
        RECT 203.835 -117.805 204.165 -117.475 ;
        RECT 203.835 -119.165 204.165 -118.835 ;
        RECT 203.835 -120.525 204.165 -120.195 ;
        RECT 203.835 -121.885 204.165 -121.555 ;
        RECT 203.835 -123.245 204.165 -122.915 ;
        RECT 203.835 -124.605 204.165 -124.275 ;
        RECT 203.835 -125.965 204.165 -125.635 ;
        RECT 203.835 -127.325 204.165 -126.995 ;
        RECT 203.835 -128.685 204.165 -128.355 ;
        RECT 203.835 -130.045 204.165 -129.715 ;
        RECT 203.835 -131.405 204.165 -131.075 ;
        RECT 203.835 -132.765 204.165 -132.435 ;
        RECT 203.835 -134.125 204.165 -133.795 ;
        RECT 203.835 -135.485 204.165 -135.155 ;
        RECT 203.835 -136.845 204.165 -136.515 ;
        RECT 203.835 -138.205 204.165 -137.875 ;
        RECT 203.835 -139.565 204.165 -139.235 ;
        RECT 203.835 -140.925 204.165 -140.595 ;
        RECT 203.835 -142.285 204.165 -141.955 ;
        RECT 203.835 -143.645 204.165 -143.315 ;
        RECT 203.835 -145.005 204.165 -144.675 ;
        RECT 203.835 -146.365 204.165 -146.035 ;
        RECT 203.835 -147.725 204.165 -147.395 ;
        RECT 203.835 -149.085 204.165 -148.755 ;
        RECT 203.835 -150.445 204.165 -150.115 ;
        RECT 203.835 -151.805 204.165 -151.475 ;
        RECT 203.835 -153.165 204.165 -152.835 ;
        RECT 203.835 -154.525 204.165 -154.195 ;
        RECT 203.835 -155.885 204.165 -155.555 ;
        RECT 203.835 -157.245 204.165 -156.915 ;
        RECT 203.835 -158.605 204.165 -158.275 ;
        RECT 203.835 -159.965 204.165 -159.635 ;
        RECT 203.835 -161.325 204.165 -160.995 ;
        RECT 203.835 -162.685 204.165 -162.355 ;
        RECT 203.835 -164.045 204.165 -163.715 ;
        RECT 203.835 -165.405 204.165 -165.075 ;
        RECT 203.835 -166.765 204.165 -166.435 ;
        RECT 203.835 -168.125 204.165 -167.795 ;
        RECT 203.835 -169.485 204.165 -169.155 ;
        RECT 203.835 -170.845 204.165 -170.515 ;
        RECT 203.835 -172.205 204.165 -171.875 ;
        RECT 203.835 -173.565 204.165 -173.235 ;
        RECT 203.835 -174.925 204.165 -174.595 ;
        RECT 203.835 -176.285 204.165 -175.955 ;
        RECT 203.835 -177.645 204.165 -177.315 ;
        RECT 203.835 -179.005 204.165 -178.675 ;
        RECT 203.835 -180.365 204.165 -180.035 ;
        RECT 203.835 -181.725 204.165 -181.395 ;
        RECT 203.835 -183.085 204.165 -182.755 ;
        RECT 203.835 -184.445 204.165 -184.115 ;
        RECT 203.835 -185.805 204.165 -185.475 ;
        RECT 203.835 -187.165 204.165 -186.835 ;
        RECT 203.835 -188.525 204.165 -188.195 ;
        RECT 203.835 -189.885 204.165 -189.555 ;
        RECT 203.835 -191.245 204.165 -190.915 ;
        RECT 203.835 -192.605 204.165 -192.275 ;
        RECT 203.835 -193.965 204.165 -193.635 ;
        RECT 203.835 -195.325 204.165 -194.995 ;
        RECT 203.835 -196.685 204.165 -196.355 ;
        RECT 203.835 -198.045 204.165 -197.715 ;
        RECT 203.835 -199.405 204.165 -199.075 ;
        RECT 203.835 -200.765 204.165 -200.435 ;
        RECT 203.835 -202.125 204.165 -201.795 ;
        RECT 203.835 -203.485 204.165 -203.155 ;
        RECT 203.835 -204.845 204.165 -204.515 ;
        RECT 203.835 -206.205 204.165 -205.875 ;
        RECT 203.835 -207.565 204.165 -207.235 ;
        RECT 203.835 -208.925 204.165 -208.595 ;
        RECT 203.835 -210.285 204.165 -209.955 ;
        RECT 203.835 -211.645 204.165 -211.315 ;
        RECT 203.835 -213.005 204.165 -212.675 ;
        RECT 203.835 -214.365 204.165 -214.035 ;
        RECT 203.835 -215.725 204.165 -215.395 ;
        RECT 203.835 -217.085 204.165 -216.755 ;
        RECT 203.835 -218.445 204.165 -218.115 ;
        RECT 203.835 -224.09 204.165 -222.96 ;
        RECT 203.84 -224.205 204.16 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.195 -211.645 205.525 -211.315 ;
        RECT 205.195 -213.005 205.525 -212.675 ;
        RECT 205.195 -214.365 205.525 -214.035 ;
        RECT 205.195 -215.725 205.525 -215.395 ;
        RECT 205.195 -217.085 205.525 -216.755 ;
        RECT 205.195 -218.445 205.525 -218.115 ;
        RECT 205.195 -224.09 205.525 -222.96 ;
        RECT 205.2 -224.205 205.52 133.765 ;
        RECT 205.195 132.52 205.525 133.65 ;
        RECT 205.195 128.355 205.525 128.685 ;
        RECT 205.195 126.995 205.525 127.325 ;
        RECT 205.195 125.635 205.525 125.965 ;
        RECT 205.195 124.275 205.525 124.605 ;
        RECT 205.195 121.41 205.525 121.74 ;
        RECT 205.195 119.235 205.525 119.565 ;
        RECT 205.195 117.655 205.525 117.985 ;
        RECT 205.195 116.805 205.525 117.135 ;
        RECT 205.195 114.495 205.525 114.825 ;
        RECT 205.195 113.645 205.525 113.975 ;
        RECT 205.195 111.335 205.525 111.665 ;
        RECT 205.195 110.485 205.525 110.815 ;
        RECT 205.195 108.175 205.525 108.505 ;
        RECT 205.195 107.325 205.525 107.655 ;
        RECT 205.195 105.015 205.525 105.345 ;
        RECT 205.195 103.435 205.525 103.765 ;
        RECT 205.195 102.585 205.525 102.915 ;
        RECT 205.195 100.275 205.525 100.605 ;
        RECT 205.195 99.425 205.525 99.755 ;
        RECT 205.195 97.115 205.525 97.445 ;
        RECT 205.195 96.265 205.525 96.595 ;
        RECT 205.195 93.955 205.525 94.285 ;
        RECT 205.195 93.105 205.525 93.435 ;
        RECT 205.195 90.795 205.525 91.125 ;
        RECT 205.195 89.215 205.525 89.545 ;
        RECT 205.195 88.365 205.525 88.695 ;
        RECT 205.195 86.055 205.525 86.385 ;
        RECT 205.195 85.205 205.525 85.535 ;
        RECT 205.195 82.895 205.525 83.225 ;
        RECT 205.195 82.045 205.525 82.375 ;
        RECT 205.195 79.735 205.525 80.065 ;
        RECT 205.195 78.885 205.525 79.215 ;
        RECT 205.195 76.575 205.525 76.905 ;
        RECT 205.195 74.995 205.525 75.325 ;
        RECT 205.195 74.145 205.525 74.475 ;
        RECT 205.195 71.835 205.525 72.165 ;
        RECT 205.195 70.985 205.525 71.315 ;
        RECT 205.195 68.675 205.525 69.005 ;
        RECT 205.195 67.825 205.525 68.155 ;
        RECT 205.195 65.515 205.525 65.845 ;
        RECT 205.195 64.665 205.525 64.995 ;
        RECT 205.195 62.355 205.525 62.685 ;
        RECT 205.195 60.775 205.525 61.105 ;
        RECT 205.195 59.925 205.525 60.255 ;
        RECT 205.195 57.615 205.525 57.945 ;
        RECT 205.195 56.765 205.525 57.095 ;
        RECT 205.195 54.455 205.525 54.785 ;
        RECT 205.195 53.605 205.525 53.935 ;
        RECT 205.195 51.295 205.525 51.625 ;
        RECT 205.195 50.445 205.525 50.775 ;
        RECT 205.195 48.135 205.525 48.465 ;
        RECT 205.195 46.555 205.525 46.885 ;
        RECT 205.195 45.705 205.525 46.035 ;
        RECT 205.195 43.395 205.525 43.725 ;
        RECT 205.195 42.545 205.525 42.875 ;
        RECT 205.195 40.235 205.525 40.565 ;
        RECT 205.195 39.385 205.525 39.715 ;
        RECT 205.195 37.075 205.525 37.405 ;
        RECT 205.195 36.225 205.525 36.555 ;
        RECT 205.195 33.915 205.525 34.245 ;
        RECT 205.195 32.335 205.525 32.665 ;
        RECT 205.195 31.485 205.525 31.815 ;
        RECT 205.195 29.175 205.525 29.505 ;
        RECT 205.195 28.325 205.525 28.655 ;
        RECT 205.195 26.015 205.525 26.345 ;
        RECT 205.195 25.165 205.525 25.495 ;
        RECT 205.195 22.855 205.525 23.185 ;
        RECT 205.195 22.005 205.525 22.335 ;
        RECT 205.195 19.695 205.525 20.025 ;
        RECT 205.195 18.115 205.525 18.445 ;
        RECT 205.195 17.265 205.525 17.595 ;
        RECT 205.195 14.955 205.525 15.285 ;
        RECT 205.195 14.105 205.525 14.435 ;
        RECT 205.195 11.795 205.525 12.125 ;
        RECT 205.195 10.945 205.525 11.275 ;
        RECT 205.195 8.635 205.525 8.965 ;
        RECT 205.195 7.785 205.525 8.115 ;
        RECT 205.195 5.475 205.525 5.805 ;
        RECT 205.195 3.895 205.525 4.225 ;
        RECT 205.195 3.045 205.525 3.375 ;
        RECT 205.195 0.87 205.525 1.2 ;
        RECT 205.195 -0.845 205.525 -0.515 ;
        RECT 205.195 -2.205 205.525 -1.875 ;
        RECT 205.195 -3.565 205.525 -3.235 ;
        RECT 205.195 -4.925 205.525 -4.595 ;
        RECT 205.195 -6.285 205.525 -5.955 ;
        RECT 205.195 -7.645 205.525 -7.315 ;
        RECT 205.195 -9.005 205.525 -8.675 ;
        RECT 205.195 -10.365 205.525 -10.035 ;
        RECT 205.195 -11.725 205.525 -11.395 ;
        RECT 205.195 -13.085 205.525 -12.755 ;
        RECT 205.195 -14.445 205.525 -14.115 ;
        RECT 205.195 -15.805 205.525 -15.475 ;
        RECT 205.195 -17.165 205.525 -16.835 ;
        RECT 205.195 -18.525 205.525 -18.195 ;
        RECT 205.195 -19.885 205.525 -19.555 ;
        RECT 205.195 -21.245 205.525 -20.915 ;
        RECT 205.195 -22.605 205.525 -22.275 ;
        RECT 205.195 -23.965 205.525 -23.635 ;
        RECT 205.195 -25.325 205.525 -24.995 ;
        RECT 205.195 -26.685 205.525 -26.355 ;
        RECT 205.195 -28.045 205.525 -27.715 ;
        RECT 205.195 -29.405 205.525 -29.075 ;
        RECT 205.195 -30.765 205.525 -30.435 ;
        RECT 205.195 -32.125 205.525 -31.795 ;
        RECT 205.195 -33.485 205.525 -33.155 ;
        RECT 205.195 -34.845 205.525 -34.515 ;
        RECT 205.195 -36.205 205.525 -35.875 ;
        RECT 205.195 -37.565 205.525 -37.235 ;
        RECT 205.195 -38.925 205.525 -38.595 ;
        RECT 205.195 -40.285 205.525 -39.955 ;
        RECT 205.195 -41.645 205.525 -41.315 ;
        RECT 205.195 -43.005 205.525 -42.675 ;
        RECT 205.195 -44.365 205.525 -44.035 ;
        RECT 205.195 -45.725 205.525 -45.395 ;
        RECT 205.195 -47.085 205.525 -46.755 ;
        RECT 205.195 -48.445 205.525 -48.115 ;
        RECT 205.195 -49.805 205.525 -49.475 ;
        RECT 205.195 -51.165 205.525 -50.835 ;
        RECT 205.195 -52.525 205.525 -52.195 ;
        RECT 205.195 -53.885 205.525 -53.555 ;
        RECT 205.195 -55.245 205.525 -54.915 ;
        RECT 205.195 -56.605 205.525 -56.275 ;
        RECT 205.195 -57.965 205.525 -57.635 ;
        RECT 205.195 -59.325 205.525 -58.995 ;
        RECT 205.195 -60.685 205.525 -60.355 ;
        RECT 205.195 -62.045 205.525 -61.715 ;
        RECT 205.195 -63.405 205.525 -63.075 ;
        RECT 205.195 -64.765 205.525 -64.435 ;
        RECT 205.195 -66.125 205.525 -65.795 ;
        RECT 205.195 -67.485 205.525 -67.155 ;
        RECT 205.195 -68.845 205.525 -68.515 ;
        RECT 205.195 -70.205 205.525 -69.875 ;
        RECT 205.195 -71.565 205.525 -71.235 ;
        RECT 205.195 -72.925 205.525 -72.595 ;
        RECT 205.195 -74.285 205.525 -73.955 ;
        RECT 205.195 -75.645 205.525 -75.315 ;
        RECT 205.195 -77.005 205.525 -76.675 ;
        RECT 205.195 -78.365 205.525 -78.035 ;
        RECT 205.195 -79.725 205.525 -79.395 ;
        RECT 205.195 -81.085 205.525 -80.755 ;
        RECT 205.195 -82.445 205.525 -82.115 ;
        RECT 205.195 -83.805 205.525 -83.475 ;
        RECT 205.195 -85.165 205.525 -84.835 ;
        RECT 205.195 -86.525 205.525 -86.195 ;
        RECT 205.195 -87.885 205.525 -87.555 ;
        RECT 205.195 -89.245 205.525 -88.915 ;
        RECT 205.195 -90.605 205.525 -90.275 ;
        RECT 205.195 -91.965 205.525 -91.635 ;
        RECT 205.195 -93.325 205.525 -92.995 ;
        RECT 205.195 -94.685 205.525 -94.355 ;
        RECT 205.195 -96.045 205.525 -95.715 ;
        RECT 205.195 -97.405 205.525 -97.075 ;
        RECT 205.195 -98.765 205.525 -98.435 ;
        RECT 205.195 -100.125 205.525 -99.795 ;
        RECT 205.195 -101.485 205.525 -101.155 ;
        RECT 205.195 -102.845 205.525 -102.515 ;
        RECT 205.195 -104.205 205.525 -103.875 ;
        RECT 205.195 -105.565 205.525 -105.235 ;
        RECT 205.195 -106.925 205.525 -106.595 ;
        RECT 205.195 -108.285 205.525 -107.955 ;
        RECT 205.195 -109.645 205.525 -109.315 ;
        RECT 205.195 -111.005 205.525 -110.675 ;
        RECT 205.195 -112.365 205.525 -112.035 ;
        RECT 205.195 -113.725 205.525 -113.395 ;
        RECT 205.195 -115.085 205.525 -114.755 ;
        RECT 205.195 -116.445 205.525 -116.115 ;
        RECT 205.195 -117.805 205.525 -117.475 ;
        RECT 205.195 -119.165 205.525 -118.835 ;
        RECT 205.195 -120.525 205.525 -120.195 ;
        RECT 205.195 -121.885 205.525 -121.555 ;
        RECT 205.195 -123.245 205.525 -122.915 ;
        RECT 205.195 -124.605 205.525 -124.275 ;
        RECT 205.195 -125.965 205.525 -125.635 ;
        RECT 205.195 -127.325 205.525 -126.995 ;
        RECT 205.195 -128.685 205.525 -128.355 ;
        RECT 205.195 -130.045 205.525 -129.715 ;
        RECT 205.195 -131.405 205.525 -131.075 ;
        RECT 205.195 -132.765 205.525 -132.435 ;
        RECT 205.195 -134.125 205.525 -133.795 ;
        RECT 205.195 -135.485 205.525 -135.155 ;
        RECT 205.195 -136.845 205.525 -136.515 ;
        RECT 205.195 -138.205 205.525 -137.875 ;
        RECT 205.195 -139.565 205.525 -139.235 ;
        RECT 205.195 -140.925 205.525 -140.595 ;
        RECT 205.195 -142.285 205.525 -141.955 ;
        RECT 205.195 -143.645 205.525 -143.315 ;
        RECT 205.195 -145.005 205.525 -144.675 ;
        RECT 205.195 -146.365 205.525 -146.035 ;
        RECT 205.195 -147.725 205.525 -147.395 ;
        RECT 205.195 -149.085 205.525 -148.755 ;
        RECT 205.195 -150.445 205.525 -150.115 ;
        RECT 205.195 -151.805 205.525 -151.475 ;
        RECT 205.195 -153.165 205.525 -152.835 ;
        RECT 205.195 -154.525 205.525 -154.195 ;
        RECT 205.195 -155.885 205.525 -155.555 ;
        RECT 205.195 -157.245 205.525 -156.915 ;
        RECT 205.195 -158.605 205.525 -158.275 ;
        RECT 205.195 -159.965 205.525 -159.635 ;
        RECT 205.195 -161.325 205.525 -160.995 ;
        RECT 205.195 -162.685 205.525 -162.355 ;
        RECT 205.195 -164.045 205.525 -163.715 ;
        RECT 205.195 -165.405 205.525 -165.075 ;
        RECT 205.195 -166.765 205.525 -166.435 ;
        RECT 205.195 -168.125 205.525 -167.795 ;
        RECT 205.195 -169.485 205.525 -169.155 ;
        RECT 205.195 -170.845 205.525 -170.515 ;
        RECT 205.195 -172.205 205.525 -171.875 ;
        RECT 205.195 -173.565 205.525 -173.235 ;
        RECT 205.195 -174.925 205.525 -174.595 ;
        RECT 205.195 -176.285 205.525 -175.955 ;
        RECT 205.195 -177.645 205.525 -177.315 ;
        RECT 205.195 -179.005 205.525 -178.675 ;
        RECT 205.195 -180.365 205.525 -180.035 ;
        RECT 205.195 -181.725 205.525 -181.395 ;
        RECT 205.195 -183.085 205.525 -182.755 ;
        RECT 205.195 -184.445 205.525 -184.115 ;
        RECT 205.195 -185.805 205.525 -185.475 ;
        RECT 205.195 -187.165 205.525 -186.835 ;
        RECT 205.195 -188.525 205.525 -188.195 ;
        RECT 205.195 -189.885 205.525 -189.555 ;
        RECT 205.195 -191.245 205.525 -190.915 ;
        RECT 205.195 -192.605 205.525 -192.275 ;
        RECT 205.195 -193.965 205.525 -193.635 ;
        RECT 205.195 -195.325 205.525 -194.995 ;
        RECT 205.195 -196.685 205.525 -196.355 ;
        RECT 205.195 -198.045 205.525 -197.715 ;
        RECT 205.195 -199.405 205.525 -199.075 ;
        RECT 205.195 -200.765 205.525 -200.435 ;
        RECT 205.195 -202.125 205.525 -201.795 ;
        RECT 205.195 -203.485 205.525 -203.155 ;
        RECT 205.195 -204.845 205.525 -204.515 ;
        RECT 205.195 -206.205 205.525 -205.875 ;
        RECT 205.195 -207.565 205.525 -207.235 ;
        RECT 205.195 -208.925 205.525 -208.595 ;
        RECT 205.195 -210.285 205.525 -209.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.115 132.52 167.445 133.65 ;
        RECT 167.115 128.355 167.445 128.685 ;
        RECT 167.115 126.995 167.445 127.325 ;
        RECT 167.115 125.635 167.445 125.965 ;
        RECT 167.115 124.275 167.445 124.605 ;
        RECT 167.12 123.6 167.44 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.115 -123.245 167.445 -122.915 ;
        RECT 167.115 -124.605 167.445 -124.275 ;
        RECT 167.115 -125.965 167.445 -125.635 ;
        RECT 167.115 -127.325 167.445 -126.995 ;
        RECT 167.115 -128.685 167.445 -128.355 ;
        RECT 167.115 -130.045 167.445 -129.715 ;
        RECT 167.115 -131.405 167.445 -131.075 ;
        RECT 167.115 -132.765 167.445 -132.435 ;
        RECT 167.115 -134.125 167.445 -133.795 ;
        RECT 167.115 -135.485 167.445 -135.155 ;
        RECT 167.115 -136.845 167.445 -136.515 ;
        RECT 167.115 -138.205 167.445 -137.875 ;
        RECT 167.115 -139.565 167.445 -139.235 ;
        RECT 167.115 -140.925 167.445 -140.595 ;
        RECT 167.115 -142.285 167.445 -141.955 ;
        RECT 167.115 -143.645 167.445 -143.315 ;
        RECT 167.115 -145.005 167.445 -144.675 ;
        RECT 167.115 -146.365 167.445 -146.035 ;
        RECT 167.115 -147.725 167.445 -147.395 ;
        RECT 167.115 -149.085 167.445 -148.755 ;
        RECT 167.115 -150.445 167.445 -150.115 ;
        RECT 167.115 -151.805 167.445 -151.475 ;
        RECT 167.115 -153.165 167.445 -152.835 ;
        RECT 167.115 -154.525 167.445 -154.195 ;
        RECT 167.115 -155.885 167.445 -155.555 ;
        RECT 167.115 -157.245 167.445 -156.915 ;
        RECT 167.115 -158.605 167.445 -158.275 ;
        RECT 167.115 -159.965 167.445 -159.635 ;
        RECT 167.115 -161.325 167.445 -160.995 ;
        RECT 167.115 -162.685 167.445 -162.355 ;
        RECT 167.115 -164.045 167.445 -163.715 ;
        RECT 167.115 -165.405 167.445 -165.075 ;
        RECT 167.115 -166.765 167.445 -166.435 ;
        RECT 167.115 -168.125 167.445 -167.795 ;
        RECT 167.115 -169.485 167.445 -169.155 ;
        RECT 167.115 -170.845 167.445 -170.515 ;
        RECT 167.115 -172.205 167.445 -171.875 ;
        RECT 167.115 -173.565 167.445 -173.235 ;
        RECT 167.115 -174.925 167.445 -174.595 ;
        RECT 167.115 -176.285 167.445 -175.955 ;
        RECT 167.115 -177.645 167.445 -177.315 ;
        RECT 167.115 -179.005 167.445 -178.675 ;
        RECT 167.115 -180.365 167.445 -180.035 ;
        RECT 167.115 -181.725 167.445 -181.395 ;
        RECT 167.115 -183.085 167.445 -182.755 ;
        RECT 167.115 -184.445 167.445 -184.115 ;
        RECT 167.115 -185.805 167.445 -185.475 ;
        RECT 167.115 -187.165 167.445 -186.835 ;
        RECT 167.115 -188.525 167.445 -188.195 ;
        RECT 167.115 -189.885 167.445 -189.555 ;
        RECT 167.115 -191.245 167.445 -190.915 ;
        RECT 167.115 -192.605 167.445 -192.275 ;
        RECT 167.115 -193.965 167.445 -193.635 ;
        RECT 167.115 -195.325 167.445 -194.995 ;
        RECT 167.115 -196.685 167.445 -196.355 ;
        RECT 167.115 -198.045 167.445 -197.715 ;
        RECT 167.115 -199.405 167.445 -199.075 ;
        RECT 167.115 -200.765 167.445 -200.435 ;
        RECT 167.115 -202.125 167.445 -201.795 ;
        RECT 167.115 -203.485 167.445 -203.155 ;
        RECT 167.115 -204.845 167.445 -204.515 ;
        RECT 167.115 -206.205 167.445 -205.875 ;
        RECT 167.115 -207.565 167.445 -207.235 ;
        RECT 167.115 -208.925 167.445 -208.595 ;
        RECT 167.115 -210.285 167.445 -209.955 ;
        RECT 167.115 -211.645 167.445 -211.315 ;
        RECT 167.115 -213.005 167.445 -212.675 ;
        RECT 167.115 -214.365 167.445 -214.035 ;
        RECT 167.115 -215.725 167.445 -215.395 ;
        RECT 167.115 -217.085 167.445 -216.755 ;
        RECT 167.115 -218.445 167.445 -218.115 ;
        RECT 167.115 -224.09 167.445 -222.96 ;
        RECT 167.12 -224.205 167.44 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.36 -121.535 167.69 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.475 132.52 168.805 133.65 ;
        RECT 168.475 128.355 168.805 128.685 ;
        RECT 168.475 126.995 168.805 127.325 ;
        RECT 168.475 125.635 168.805 125.965 ;
        RECT 168.475 124.275 168.805 124.605 ;
        RECT 168.48 123.6 168.8 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.835 132.52 170.165 133.65 ;
        RECT 169.835 128.355 170.165 128.685 ;
        RECT 169.835 126.995 170.165 127.325 ;
        RECT 169.835 125.635 170.165 125.965 ;
        RECT 169.835 124.275 170.165 124.605 ;
        RECT 169.84 123.6 170.16 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.835 -0.845 170.165 -0.515 ;
        RECT 169.835 -2.205 170.165 -1.875 ;
        RECT 169.835 -3.565 170.165 -3.235 ;
        RECT 169.84 -3.565 170.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.195 132.52 171.525 133.65 ;
        RECT 171.195 128.355 171.525 128.685 ;
        RECT 171.195 126.995 171.525 127.325 ;
        RECT 171.195 125.635 171.525 125.965 ;
        RECT 171.195 124.275 171.525 124.605 ;
        RECT 171.2 123.6 171.52 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.195 -0.845 171.525 -0.515 ;
        RECT 171.195 -2.205 171.525 -1.875 ;
        RECT 171.195 -3.565 171.525 -3.235 ;
        RECT 171.2 -3.565 171.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.195 -119.165 171.525 -118.835 ;
        RECT 171.195 -120.525 171.525 -120.195 ;
        RECT 171.195 -121.885 171.525 -121.555 ;
        RECT 171.195 -123.245 171.525 -122.915 ;
        RECT 171.195 -124.605 171.525 -124.275 ;
        RECT 171.195 -125.965 171.525 -125.635 ;
        RECT 171.195 -127.325 171.525 -126.995 ;
        RECT 171.195 -128.685 171.525 -128.355 ;
        RECT 171.195 -130.045 171.525 -129.715 ;
        RECT 171.195 -131.405 171.525 -131.075 ;
        RECT 171.195 -132.765 171.525 -132.435 ;
        RECT 171.195 -134.125 171.525 -133.795 ;
        RECT 171.195 -135.485 171.525 -135.155 ;
        RECT 171.195 -136.845 171.525 -136.515 ;
        RECT 171.195 -138.205 171.525 -137.875 ;
        RECT 171.195 -139.565 171.525 -139.235 ;
        RECT 171.195 -140.925 171.525 -140.595 ;
        RECT 171.195 -142.285 171.525 -141.955 ;
        RECT 171.195 -143.645 171.525 -143.315 ;
        RECT 171.195 -145.005 171.525 -144.675 ;
        RECT 171.195 -146.365 171.525 -146.035 ;
        RECT 171.195 -147.725 171.525 -147.395 ;
        RECT 171.195 -149.085 171.525 -148.755 ;
        RECT 171.195 -150.445 171.525 -150.115 ;
        RECT 171.195 -151.805 171.525 -151.475 ;
        RECT 171.195 -153.165 171.525 -152.835 ;
        RECT 171.195 -154.525 171.525 -154.195 ;
        RECT 171.195 -155.885 171.525 -155.555 ;
        RECT 171.195 -157.245 171.525 -156.915 ;
        RECT 171.195 -158.605 171.525 -158.275 ;
        RECT 171.195 -159.965 171.525 -159.635 ;
        RECT 171.195 -161.325 171.525 -160.995 ;
        RECT 171.195 -162.685 171.525 -162.355 ;
        RECT 171.195 -164.045 171.525 -163.715 ;
        RECT 171.195 -165.405 171.525 -165.075 ;
        RECT 171.195 -166.765 171.525 -166.435 ;
        RECT 171.195 -168.125 171.525 -167.795 ;
        RECT 171.195 -169.485 171.525 -169.155 ;
        RECT 171.195 -170.845 171.525 -170.515 ;
        RECT 171.195 -172.205 171.525 -171.875 ;
        RECT 171.195 -173.565 171.525 -173.235 ;
        RECT 171.195 -174.925 171.525 -174.595 ;
        RECT 171.195 -176.285 171.525 -175.955 ;
        RECT 171.195 -177.645 171.525 -177.315 ;
        RECT 171.195 -179.005 171.525 -178.675 ;
        RECT 171.195 -180.365 171.525 -180.035 ;
        RECT 171.195 -181.725 171.525 -181.395 ;
        RECT 171.195 -183.085 171.525 -182.755 ;
        RECT 171.195 -184.445 171.525 -184.115 ;
        RECT 171.195 -185.805 171.525 -185.475 ;
        RECT 171.195 -187.165 171.525 -186.835 ;
        RECT 171.195 -188.525 171.525 -188.195 ;
        RECT 171.195 -189.885 171.525 -189.555 ;
        RECT 171.195 -191.245 171.525 -190.915 ;
        RECT 171.195 -192.605 171.525 -192.275 ;
        RECT 171.195 -193.965 171.525 -193.635 ;
        RECT 171.195 -195.325 171.525 -194.995 ;
        RECT 171.195 -196.685 171.525 -196.355 ;
        RECT 171.195 -198.045 171.525 -197.715 ;
        RECT 171.195 -199.405 171.525 -199.075 ;
        RECT 171.195 -200.765 171.525 -200.435 ;
        RECT 171.195 -202.125 171.525 -201.795 ;
        RECT 171.195 -203.485 171.525 -203.155 ;
        RECT 171.195 -204.845 171.525 -204.515 ;
        RECT 171.195 -206.205 171.525 -205.875 ;
        RECT 171.195 -207.565 171.525 -207.235 ;
        RECT 171.195 -208.925 171.525 -208.595 ;
        RECT 171.195 -210.285 171.525 -209.955 ;
        RECT 171.195 -211.645 171.525 -211.315 ;
        RECT 171.195 -213.005 171.525 -212.675 ;
        RECT 171.195 -214.365 171.525 -214.035 ;
        RECT 171.195 -215.725 171.525 -215.395 ;
        RECT 171.195 -217.085 171.525 -216.755 ;
        RECT 171.195 -218.445 171.525 -218.115 ;
        RECT 171.195 -224.09 171.525 -222.96 ;
        RECT 171.2 -224.205 171.52 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.555 132.52 172.885 133.65 ;
        RECT 172.555 128.355 172.885 128.685 ;
        RECT 172.555 126.995 172.885 127.325 ;
        RECT 172.555 125.635 172.885 125.965 ;
        RECT 172.555 124.275 172.885 124.605 ;
        RECT 172.56 123.6 172.88 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.555 -0.845 172.885 -0.515 ;
        RECT 172.555 -2.205 172.885 -1.875 ;
        RECT 172.555 -3.565 172.885 -3.235 ;
        RECT 172.56 -3.565 172.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.555 -119.165 172.885 -118.835 ;
        RECT 172.555 -120.525 172.885 -120.195 ;
        RECT 172.555 -121.885 172.885 -121.555 ;
        RECT 172.555 -123.245 172.885 -122.915 ;
        RECT 172.555 -124.605 172.885 -124.275 ;
        RECT 172.555 -125.965 172.885 -125.635 ;
        RECT 172.555 -127.325 172.885 -126.995 ;
        RECT 172.555 -128.685 172.885 -128.355 ;
        RECT 172.555 -130.045 172.885 -129.715 ;
        RECT 172.555 -131.405 172.885 -131.075 ;
        RECT 172.555 -132.765 172.885 -132.435 ;
        RECT 172.555 -134.125 172.885 -133.795 ;
        RECT 172.555 -135.485 172.885 -135.155 ;
        RECT 172.555 -136.845 172.885 -136.515 ;
        RECT 172.555 -138.205 172.885 -137.875 ;
        RECT 172.555 -139.565 172.885 -139.235 ;
        RECT 172.555 -140.925 172.885 -140.595 ;
        RECT 172.555 -142.285 172.885 -141.955 ;
        RECT 172.555 -143.645 172.885 -143.315 ;
        RECT 172.555 -145.005 172.885 -144.675 ;
        RECT 172.555 -146.365 172.885 -146.035 ;
        RECT 172.555 -147.725 172.885 -147.395 ;
        RECT 172.555 -149.085 172.885 -148.755 ;
        RECT 172.555 -150.445 172.885 -150.115 ;
        RECT 172.555 -151.805 172.885 -151.475 ;
        RECT 172.555 -153.165 172.885 -152.835 ;
        RECT 172.555 -154.525 172.885 -154.195 ;
        RECT 172.555 -155.885 172.885 -155.555 ;
        RECT 172.555 -157.245 172.885 -156.915 ;
        RECT 172.555 -158.605 172.885 -158.275 ;
        RECT 172.555 -159.965 172.885 -159.635 ;
        RECT 172.555 -161.325 172.885 -160.995 ;
        RECT 172.555 -162.685 172.885 -162.355 ;
        RECT 172.555 -164.045 172.885 -163.715 ;
        RECT 172.555 -165.405 172.885 -165.075 ;
        RECT 172.555 -166.765 172.885 -166.435 ;
        RECT 172.555 -168.125 172.885 -167.795 ;
        RECT 172.555 -169.485 172.885 -169.155 ;
        RECT 172.555 -170.845 172.885 -170.515 ;
        RECT 172.555 -172.205 172.885 -171.875 ;
        RECT 172.555 -173.565 172.885 -173.235 ;
        RECT 172.555 -174.925 172.885 -174.595 ;
        RECT 172.555 -176.285 172.885 -175.955 ;
        RECT 172.555 -177.645 172.885 -177.315 ;
        RECT 172.555 -179.005 172.885 -178.675 ;
        RECT 172.555 -180.365 172.885 -180.035 ;
        RECT 172.555 -181.725 172.885 -181.395 ;
        RECT 172.555 -183.085 172.885 -182.755 ;
        RECT 172.555 -184.445 172.885 -184.115 ;
        RECT 172.555 -185.805 172.885 -185.475 ;
        RECT 172.555 -187.165 172.885 -186.835 ;
        RECT 172.555 -188.525 172.885 -188.195 ;
        RECT 172.555 -189.885 172.885 -189.555 ;
        RECT 172.555 -191.245 172.885 -190.915 ;
        RECT 172.555 -192.605 172.885 -192.275 ;
        RECT 172.555 -193.965 172.885 -193.635 ;
        RECT 172.555 -195.325 172.885 -194.995 ;
        RECT 172.555 -196.685 172.885 -196.355 ;
        RECT 172.555 -198.045 172.885 -197.715 ;
        RECT 172.555 -199.405 172.885 -199.075 ;
        RECT 172.555 -200.765 172.885 -200.435 ;
        RECT 172.555 -202.125 172.885 -201.795 ;
        RECT 172.555 -203.485 172.885 -203.155 ;
        RECT 172.555 -204.845 172.885 -204.515 ;
        RECT 172.555 -206.205 172.885 -205.875 ;
        RECT 172.555 -207.565 172.885 -207.235 ;
        RECT 172.555 -208.925 172.885 -208.595 ;
        RECT 172.555 -210.285 172.885 -209.955 ;
        RECT 172.555 -211.645 172.885 -211.315 ;
        RECT 172.555 -213.005 172.885 -212.675 ;
        RECT 172.555 -214.365 172.885 -214.035 ;
        RECT 172.555 -215.725 172.885 -215.395 ;
        RECT 172.555 -217.085 172.885 -216.755 ;
        RECT 172.555 -218.445 172.885 -218.115 ;
        RECT 172.555 -224.09 172.885 -222.96 ;
        RECT 172.56 -224.205 172.88 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.46 -121.535 173.79 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.915 132.52 174.245 133.65 ;
        RECT 173.915 128.355 174.245 128.685 ;
        RECT 173.915 126.995 174.245 127.325 ;
        RECT 173.915 125.635 174.245 125.965 ;
        RECT 173.915 124.275 174.245 124.605 ;
        RECT 173.92 123.6 174.24 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.915 -123.245 174.245 -122.915 ;
        RECT 173.915 -124.605 174.245 -124.275 ;
        RECT 173.915 -125.965 174.245 -125.635 ;
        RECT 173.915 -127.325 174.245 -126.995 ;
        RECT 173.915 -128.685 174.245 -128.355 ;
        RECT 173.915 -130.045 174.245 -129.715 ;
        RECT 173.915 -131.405 174.245 -131.075 ;
        RECT 173.915 -132.765 174.245 -132.435 ;
        RECT 173.915 -134.125 174.245 -133.795 ;
        RECT 173.915 -135.485 174.245 -135.155 ;
        RECT 173.915 -136.845 174.245 -136.515 ;
        RECT 173.915 -138.205 174.245 -137.875 ;
        RECT 173.915 -139.565 174.245 -139.235 ;
        RECT 173.915 -140.925 174.245 -140.595 ;
        RECT 173.915 -142.285 174.245 -141.955 ;
        RECT 173.915 -143.645 174.245 -143.315 ;
        RECT 173.915 -145.005 174.245 -144.675 ;
        RECT 173.915 -146.365 174.245 -146.035 ;
        RECT 173.915 -147.725 174.245 -147.395 ;
        RECT 173.915 -149.085 174.245 -148.755 ;
        RECT 173.915 -150.445 174.245 -150.115 ;
        RECT 173.915 -151.805 174.245 -151.475 ;
        RECT 173.915 -153.165 174.245 -152.835 ;
        RECT 173.915 -154.525 174.245 -154.195 ;
        RECT 173.915 -155.885 174.245 -155.555 ;
        RECT 173.915 -157.245 174.245 -156.915 ;
        RECT 173.915 -158.605 174.245 -158.275 ;
        RECT 173.915 -159.965 174.245 -159.635 ;
        RECT 173.915 -161.325 174.245 -160.995 ;
        RECT 173.915 -162.685 174.245 -162.355 ;
        RECT 173.915 -164.045 174.245 -163.715 ;
        RECT 173.915 -165.405 174.245 -165.075 ;
        RECT 173.915 -166.765 174.245 -166.435 ;
        RECT 173.915 -168.125 174.245 -167.795 ;
        RECT 173.915 -169.485 174.245 -169.155 ;
        RECT 173.915 -170.845 174.245 -170.515 ;
        RECT 173.915 -172.205 174.245 -171.875 ;
        RECT 173.915 -173.565 174.245 -173.235 ;
        RECT 173.915 -174.925 174.245 -174.595 ;
        RECT 173.915 -176.285 174.245 -175.955 ;
        RECT 173.915 -177.645 174.245 -177.315 ;
        RECT 173.915 -179.005 174.245 -178.675 ;
        RECT 173.915 -180.365 174.245 -180.035 ;
        RECT 173.915 -181.725 174.245 -181.395 ;
        RECT 173.915 -183.085 174.245 -182.755 ;
        RECT 173.915 -184.445 174.245 -184.115 ;
        RECT 173.915 -185.805 174.245 -185.475 ;
        RECT 173.915 -187.165 174.245 -186.835 ;
        RECT 173.915 -188.525 174.245 -188.195 ;
        RECT 173.915 -189.885 174.245 -189.555 ;
        RECT 173.915 -191.245 174.245 -190.915 ;
        RECT 173.915 -192.605 174.245 -192.275 ;
        RECT 173.915 -193.965 174.245 -193.635 ;
        RECT 173.915 -195.325 174.245 -194.995 ;
        RECT 173.915 -196.685 174.245 -196.355 ;
        RECT 173.915 -198.045 174.245 -197.715 ;
        RECT 173.915 -199.405 174.245 -199.075 ;
        RECT 173.915 -200.765 174.245 -200.435 ;
        RECT 173.915 -202.125 174.245 -201.795 ;
        RECT 173.915 -203.485 174.245 -203.155 ;
        RECT 173.915 -204.845 174.245 -204.515 ;
        RECT 173.915 -206.205 174.245 -205.875 ;
        RECT 173.915 -207.565 174.245 -207.235 ;
        RECT 173.915 -208.925 174.245 -208.595 ;
        RECT 173.915 -210.285 174.245 -209.955 ;
        RECT 173.915 -211.645 174.245 -211.315 ;
        RECT 173.915 -213.005 174.245 -212.675 ;
        RECT 173.915 -214.365 174.245 -214.035 ;
        RECT 173.915 -215.725 174.245 -215.395 ;
        RECT 173.915 -217.085 174.245 -216.755 ;
        RECT 173.915 -218.445 174.245 -218.115 ;
        RECT 173.915 -224.09 174.245 -222.96 ;
        RECT 173.92 -224.205 174.24 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.275 132.52 175.605 133.65 ;
        RECT 175.275 128.355 175.605 128.685 ;
        RECT 175.275 126.995 175.605 127.325 ;
        RECT 175.275 125.635 175.605 125.965 ;
        RECT 175.275 124.275 175.605 124.605 ;
        RECT 175.28 123.6 175.6 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.275 -0.845 175.605 -0.515 ;
        RECT 175.275 -2.205 175.605 -1.875 ;
        RECT 175.275 -3.565 175.605 -3.235 ;
        RECT 175.28 -3.565 175.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 176.635 132.52 176.965 133.65 ;
        RECT 176.635 128.355 176.965 128.685 ;
        RECT 176.635 126.995 176.965 127.325 ;
        RECT 176.635 125.635 176.965 125.965 ;
        RECT 176.635 124.275 176.965 124.605 ;
        RECT 176.64 123.6 176.96 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 176.635 -0.845 176.965 -0.515 ;
        RECT 176.635 -2.205 176.965 -1.875 ;
        RECT 176.635 -3.565 176.965 -3.235 ;
        RECT 176.64 -3.565 176.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.995 132.52 178.325 133.65 ;
        RECT 177.995 128.355 178.325 128.685 ;
        RECT 177.995 126.995 178.325 127.325 ;
        RECT 177.995 125.635 178.325 125.965 ;
        RECT 177.995 124.275 178.325 124.605 ;
        RECT 178 123.6 178.32 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.995 -0.845 178.325 -0.515 ;
        RECT 177.995 -2.205 178.325 -1.875 ;
        RECT 177.995 -3.565 178.325 -3.235 ;
        RECT 178 -3.565 178.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.995 -119.165 178.325 -118.835 ;
        RECT 177.995 -120.525 178.325 -120.195 ;
        RECT 177.995 -121.885 178.325 -121.555 ;
        RECT 177.995 -123.245 178.325 -122.915 ;
        RECT 177.995 -124.605 178.325 -124.275 ;
        RECT 177.995 -125.965 178.325 -125.635 ;
        RECT 177.995 -127.325 178.325 -126.995 ;
        RECT 177.995 -128.685 178.325 -128.355 ;
        RECT 177.995 -130.045 178.325 -129.715 ;
        RECT 177.995 -131.405 178.325 -131.075 ;
        RECT 177.995 -132.765 178.325 -132.435 ;
        RECT 177.995 -134.125 178.325 -133.795 ;
        RECT 177.995 -135.485 178.325 -135.155 ;
        RECT 177.995 -136.845 178.325 -136.515 ;
        RECT 177.995 -138.205 178.325 -137.875 ;
        RECT 177.995 -139.565 178.325 -139.235 ;
        RECT 177.995 -140.925 178.325 -140.595 ;
        RECT 177.995 -142.285 178.325 -141.955 ;
        RECT 177.995 -143.645 178.325 -143.315 ;
        RECT 177.995 -145.005 178.325 -144.675 ;
        RECT 177.995 -146.365 178.325 -146.035 ;
        RECT 177.995 -147.725 178.325 -147.395 ;
        RECT 177.995 -149.085 178.325 -148.755 ;
        RECT 177.995 -150.445 178.325 -150.115 ;
        RECT 177.995 -151.805 178.325 -151.475 ;
        RECT 177.995 -153.165 178.325 -152.835 ;
        RECT 177.995 -154.525 178.325 -154.195 ;
        RECT 177.995 -155.885 178.325 -155.555 ;
        RECT 177.995 -157.245 178.325 -156.915 ;
        RECT 177.995 -158.605 178.325 -158.275 ;
        RECT 177.995 -159.965 178.325 -159.635 ;
        RECT 177.995 -161.325 178.325 -160.995 ;
        RECT 177.995 -162.685 178.325 -162.355 ;
        RECT 177.995 -164.045 178.325 -163.715 ;
        RECT 177.995 -165.405 178.325 -165.075 ;
        RECT 177.995 -166.765 178.325 -166.435 ;
        RECT 177.995 -168.125 178.325 -167.795 ;
        RECT 177.995 -169.485 178.325 -169.155 ;
        RECT 177.995 -170.845 178.325 -170.515 ;
        RECT 177.995 -172.205 178.325 -171.875 ;
        RECT 177.995 -173.565 178.325 -173.235 ;
        RECT 177.995 -174.925 178.325 -174.595 ;
        RECT 177.995 -176.285 178.325 -175.955 ;
        RECT 177.995 -177.645 178.325 -177.315 ;
        RECT 177.995 -179.005 178.325 -178.675 ;
        RECT 177.995 -180.365 178.325 -180.035 ;
        RECT 177.995 -181.725 178.325 -181.395 ;
        RECT 177.995 -183.085 178.325 -182.755 ;
        RECT 177.995 -184.445 178.325 -184.115 ;
        RECT 177.995 -185.805 178.325 -185.475 ;
        RECT 177.995 -187.165 178.325 -186.835 ;
        RECT 177.995 -188.525 178.325 -188.195 ;
        RECT 177.995 -189.885 178.325 -189.555 ;
        RECT 177.995 -191.245 178.325 -190.915 ;
        RECT 177.995 -192.605 178.325 -192.275 ;
        RECT 177.995 -193.965 178.325 -193.635 ;
        RECT 177.995 -195.325 178.325 -194.995 ;
        RECT 177.995 -196.685 178.325 -196.355 ;
        RECT 177.995 -198.045 178.325 -197.715 ;
        RECT 177.995 -199.405 178.325 -199.075 ;
        RECT 177.995 -200.765 178.325 -200.435 ;
        RECT 177.995 -202.125 178.325 -201.795 ;
        RECT 177.995 -203.485 178.325 -203.155 ;
        RECT 177.995 -204.845 178.325 -204.515 ;
        RECT 177.995 -206.205 178.325 -205.875 ;
        RECT 177.995 -207.565 178.325 -207.235 ;
        RECT 177.995 -208.925 178.325 -208.595 ;
        RECT 177.995 -210.285 178.325 -209.955 ;
        RECT 177.995 -211.645 178.325 -211.315 ;
        RECT 177.995 -213.005 178.325 -212.675 ;
        RECT 177.995 -214.365 178.325 -214.035 ;
        RECT 177.995 -215.725 178.325 -215.395 ;
        RECT 177.995 -217.085 178.325 -216.755 ;
        RECT 177.995 -218.445 178.325 -218.115 ;
        RECT 177.995 -224.09 178.325 -222.96 ;
        RECT 178 -224.205 178.32 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.355 132.52 179.685 133.65 ;
        RECT 179.355 128.355 179.685 128.685 ;
        RECT 179.355 126.995 179.685 127.325 ;
        RECT 179.355 125.635 179.685 125.965 ;
        RECT 179.355 124.275 179.685 124.605 ;
        RECT 179.36 123.6 179.68 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.355 -123.245 179.685 -122.915 ;
        RECT 179.355 -124.605 179.685 -124.275 ;
        RECT 179.355 -125.965 179.685 -125.635 ;
        RECT 179.355 -127.325 179.685 -126.995 ;
        RECT 179.355 -128.685 179.685 -128.355 ;
        RECT 179.355 -130.045 179.685 -129.715 ;
        RECT 179.355 -131.405 179.685 -131.075 ;
        RECT 179.355 -132.765 179.685 -132.435 ;
        RECT 179.355 -134.125 179.685 -133.795 ;
        RECT 179.355 -135.485 179.685 -135.155 ;
        RECT 179.355 -136.845 179.685 -136.515 ;
        RECT 179.355 -138.205 179.685 -137.875 ;
        RECT 179.355 -139.565 179.685 -139.235 ;
        RECT 179.355 -140.925 179.685 -140.595 ;
        RECT 179.355 -142.285 179.685 -141.955 ;
        RECT 179.355 -143.645 179.685 -143.315 ;
        RECT 179.355 -145.005 179.685 -144.675 ;
        RECT 179.355 -146.365 179.685 -146.035 ;
        RECT 179.355 -147.725 179.685 -147.395 ;
        RECT 179.355 -149.085 179.685 -148.755 ;
        RECT 179.355 -150.445 179.685 -150.115 ;
        RECT 179.355 -151.805 179.685 -151.475 ;
        RECT 179.355 -153.165 179.685 -152.835 ;
        RECT 179.355 -154.525 179.685 -154.195 ;
        RECT 179.355 -155.885 179.685 -155.555 ;
        RECT 179.355 -157.245 179.685 -156.915 ;
        RECT 179.355 -158.605 179.685 -158.275 ;
        RECT 179.355 -159.965 179.685 -159.635 ;
        RECT 179.355 -161.325 179.685 -160.995 ;
        RECT 179.355 -162.685 179.685 -162.355 ;
        RECT 179.355 -164.045 179.685 -163.715 ;
        RECT 179.355 -165.405 179.685 -165.075 ;
        RECT 179.355 -166.765 179.685 -166.435 ;
        RECT 179.355 -168.125 179.685 -167.795 ;
        RECT 179.355 -169.485 179.685 -169.155 ;
        RECT 179.355 -170.845 179.685 -170.515 ;
        RECT 179.355 -172.205 179.685 -171.875 ;
        RECT 179.355 -173.565 179.685 -173.235 ;
        RECT 179.355 -174.925 179.685 -174.595 ;
        RECT 179.355 -176.285 179.685 -175.955 ;
        RECT 179.355 -177.645 179.685 -177.315 ;
        RECT 179.355 -179.005 179.685 -178.675 ;
        RECT 179.355 -180.365 179.685 -180.035 ;
        RECT 179.355 -181.725 179.685 -181.395 ;
        RECT 179.355 -183.085 179.685 -182.755 ;
        RECT 179.355 -184.445 179.685 -184.115 ;
        RECT 179.355 -185.805 179.685 -185.475 ;
        RECT 179.355 -187.165 179.685 -186.835 ;
        RECT 179.355 -188.525 179.685 -188.195 ;
        RECT 179.355 -189.885 179.685 -189.555 ;
        RECT 179.355 -191.245 179.685 -190.915 ;
        RECT 179.355 -192.605 179.685 -192.275 ;
        RECT 179.355 -193.965 179.685 -193.635 ;
        RECT 179.355 -195.325 179.685 -194.995 ;
        RECT 179.355 -196.685 179.685 -196.355 ;
        RECT 179.355 -198.045 179.685 -197.715 ;
        RECT 179.355 -199.405 179.685 -199.075 ;
        RECT 179.355 -200.765 179.685 -200.435 ;
        RECT 179.355 -202.125 179.685 -201.795 ;
        RECT 179.355 -203.485 179.685 -203.155 ;
        RECT 179.355 -204.845 179.685 -204.515 ;
        RECT 179.355 -206.205 179.685 -205.875 ;
        RECT 179.355 -207.565 179.685 -207.235 ;
        RECT 179.355 -208.925 179.685 -208.595 ;
        RECT 179.355 -210.285 179.685 -209.955 ;
        RECT 179.355 -211.645 179.685 -211.315 ;
        RECT 179.355 -213.005 179.685 -212.675 ;
        RECT 179.355 -214.365 179.685 -214.035 ;
        RECT 179.355 -215.725 179.685 -215.395 ;
        RECT 179.355 -217.085 179.685 -216.755 ;
        RECT 179.355 -218.445 179.685 -218.115 ;
        RECT 179.355 -224.09 179.685 -222.96 ;
        RECT 179.36 -224.205 179.68 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.56 -121.535 179.89 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.715 132.52 181.045 133.65 ;
        RECT 180.715 128.355 181.045 128.685 ;
        RECT 180.715 126.995 181.045 127.325 ;
        RECT 180.715 125.635 181.045 125.965 ;
        RECT 180.715 124.275 181.045 124.605 ;
        RECT 180.72 123.6 181.04 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.075 132.52 182.405 133.65 ;
        RECT 182.075 128.355 182.405 128.685 ;
        RECT 182.075 126.995 182.405 127.325 ;
        RECT 182.075 125.635 182.405 125.965 ;
        RECT 182.075 124.275 182.405 124.605 ;
        RECT 182.08 123.6 182.4 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.075 -0.845 182.405 -0.515 ;
        RECT 182.075 -2.205 182.405 -1.875 ;
        RECT 182.075 -3.565 182.405 -3.235 ;
        RECT 182.08 -3.565 182.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.435 132.52 183.765 133.65 ;
        RECT 183.435 128.355 183.765 128.685 ;
        RECT 183.435 126.995 183.765 127.325 ;
        RECT 183.435 125.635 183.765 125.965 ;
        RECT 183.435 124.275 183.765 124.605 ;
        RECT 183.44 123.6 183.76 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.435 -0.845 183.765 -0.515 ;
        RECT 183.435 -2.205 183.765 -1.875 ;
        RECT 183.435 -3.565 183.765 -3.235 ;
        RECT 183.44 -3.565 183.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.435 -119.165 183.765 -118.835 ;
        RECT 183.435 -120.525 183.765 -120.195 ;
        RECT 183.435 -121.885 183.765 -121.555 ;
        RECT 183.435 -123.245 183.765 -122.915 ;
        RECT 183.435 -124.605 183.765 -124.275 ;
        RECT 183.435 -125.965 183.765 -125.635 ;
        RECT 183.435 -127.325 183.765 -126.995 ;
        RECT 183.435 -128.685 183.765 -128.355 ;
        RECT 183.435 -130.045 183.765 -129.715 ;
        RECT 183.435 -131.405 183.765 -131.075 ;
        RECT 183.435 -132.765 183.765 -132.435 ;
        RECT 183.435 -134.125 183.765 -133.795 ;
        RECT 183.435 -135.485 183.765 -135.155 ;
        RECT 183.435 -136.845 183.765 -136.515 ;
        RECT 183.435 -138.205 183.765 -137.875 ;
        RECT 183.435 -139.565 183.765 -139.235 ;
        RECT 183.435 -140.925 183.765 -140.595 ;
        RECT 183.435 -142.285 183.765 -141.955 ;
        RECT 183.435 -143.645 183.765 -143.315 ;
        RECT 183.435 -145.005 183.765 -144.675 ;
        RECT 183.435 -146.365 183.765 -146.035 ;
        RECT 183.435 -147.725 183.765 -147.395 ;
        RECT 183.435 -149.085 183.765 -148.755 ;
        RECT 183.435 -150.445 183.765 -150.115 ;
        RECT 183.435 -151.805 183.765 -151.475 ;
        RECT 183.435 -153.165 183.765 -152.835 ;
        RECT 183.435 -154.525 183.765 -154.195 ;
        RECT 183.435 -155.885 183.765 -155.555 ;
        RECT 183.435 -157.245 183.765 -156.915 ;
        RECT 183.435 -158.605 183.765 -158.275 ;
        RECT 183.435 -159.965 183.765 -159.635 ;
        RECT 183.435 -161.325 183.765 -160.995 ;
        RECT 183.435 -162.685 183.765 -162.355 ;
        RECT 183.435 -164.045 183.765 -163.715 ;
        RECT 183.435 -165.405 183.765 -165.075 ;
        RECT 183.435 -166.765 183.765 -166.435 ;
        RECT 183.435 -168.125 183.765 -167.795 ;
        RECT 183.435 -169.485 183.765 -169.155 ;
        RECT 183.435 -170.845 183.765 -170.515 ;
        RECT 183.435 -172.205 183.765 -171.875 ;
        RECT 183.435 -173.565 183.765 -173.235 ;
        RECT 183.435 -174.925 183.765 -174.595 ;
        RECT 183.435 -176.285 183.765 -175.955 ;
        RECT 183.435 -177.645 183.765 -177.315 ;
        RECT 183.435 -179.005 183.765 -178.675 ;
        RECT 183.435 -180.365 183.765 -180.035 ;
        RECT 183.435 -181.725 183.765 -181.395 ;
        RECT 183.435 -183.085 183.765 -182.755 ;
        RECT 183.435 -184.445 183.765 -184.115 ;
        RECT 183.435 -185.805 183.765 -185.475 ;
        RECT 183.435 -187.165 183.765 -186.835 ;
        RECT 183.435 -188.525 183.765 -188.195 ;
        RECT 183.435 -189.885 183.765 -189.555 ;
        RECT 183.435 -191.245 183.765 -190.915 ;
        RECT 183.435 -192.605 183.765 -192.275 ;
        RECT 183.435 -193.965 183.765 -193.635 ;
        RECT 183.435 -195.325 183.765 -194.995 ;
        RECT 183.435 -196.685 183.765 -196.355 ;
        RECT 183.435 -198.045 183.765 -197.715 ;
        RECT 183.435 -199.405 183.765 -199.075 ;
        RECT 183.435 -200.765 183.765 -200.435 ;
        RECT 183.435 -202.125 183.765 -201.795 ;
        RECT 183.435 -203.485 183.765 -203.155 ;
        RECT 183.435 -204.845 183.765 -204.515 ;
        RECT 183.435 -206.205 183.765 -205.875 ;
        RECT 183.435 -207.565 183.765 -207.235 ;
        RECT 183.435 -208.925 183.765 -208.595 ;
        RECT 183.435 -210.285 183.765 -209.955 ;
        RECT 183.435 -211.645 183.765 -211.315 ;
        RECT 183.435 -213.005 183.765 -212.675 ;
        RECT 183.435 -214.365 183.765 -214.035 ;
        RECT 183.435 -215.725 183.765 -215.395 ;
        RECT 183.435 -217.085 183.765 -216.755 ;
        RECT 183.435 -218.445 183.765 -218.115 ;
        RECT 183.435 -224.09 183.765 -222.96 ;
        RECT 183.44 -224.205 183.76 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.795 132.52 185.125 133.65 ;
        RECT 184.795 128.355 185.125 128.685 ;
        RECT 184.795 126.995 185.125 127.325 ;
        RECT 184.795 125.635 185.125 125.965 ;
        RECT 184.795 124.275 185.125 124.605 ;
        RECT 184.8 123.6 185.12 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.795 -0.845 185.125 -0.515 ;
        RECT 184.795 -2.205 185.125 -1.875 ;
        RECT 184.795 -3.565 185.125 -3.235 ;
        RECT 184.8 -3.565 185.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.795 -119.165 185.125 -118.835 ;
        RECT 184.795 -120.525 185.125 -120.195 ;
        RECT 184.795 -121.885 185.125 -121.555 ;
        RECT 184.795 -123.245 185.125 -122.915 ;
        RECT 184.795 -124.605 185.125 -124.275 ;
        RECT 184.795 -125.965 185.125 -125.635 ;
        RECT 184.795 -127.325 185.125 -126.995 ;
        RECT 184.795 -128.685 185.125 -128.355 ;
        RECT 184.795 -130.045 185.125 -129.715 ;
        RECT 184.795 -131.405 185.125 -131.075 ;
        RECT 184.795 -132.765 185.125 -132.435 ;
        RECT 184.795 -134.125 185.125 -133.795 ;
        RECT 184.795 -135.485 185.125 -135.155 ;
        RECT 184.795 -136.845 185.125 -136.515 ;
        RECT 184.795 -138.205 185.125 -137.875 ;
        RECT 184.795 -139.565 185.125 -139.235 ;
        RECT 184.795 -140.925 185.125 -140.595 ;
        RECT 184.795 -142.285 185.125 -141.955 ;
        RECT 184.795 -143.645 185.125 -143.315 ;
        RECT 184.795 -145.005 185.125 -144.675 ;
        RECT 184.795 -146.365 185.125 -146.035 ;
        RECT 184.795 -147.725 185.125 -147.395 ;
        RECT 184.795 -149.085 185.125 -148.755 ;
        RECT 184.795 -150.445 185.125 -150.115 ;
        RECT 184.795 -151.805 185.125 -151.475 ;
        RECT 184.795 -153.165 185.125 -152.835 ;
        RECT 184.795 -154.525 185.125 -154.195 ;
        RECT 184.795 -155.885 185.125 -155.555 ;
        RECT 184.795 -157.245 185.125 -156.915 ;
        RECT 184.795 -158.605 185.125 -158.275 ;
        RECT 184.795 -159.965 185.125 -159.635 ;
        RECT 184.795 -161.325 185.125 -160.995 ;
        RECT 184.795 -162.685 185.125 -162.355 ;
        RECT 184.795 -164.045 185.125 -163.715 ;
        RECT 184.795 -165.405 185.125 -165.075 ;
        RECT 184.795 -166.765 185.125 -166.435 ;
        RECT 184.795 -168.125 185.125 -167.795 ;
        RECT 184.795 -169.485 185.125 -169.155 ;
        RECT 184.795 -170.845 185.125 -170.515 ;
        RECT 184.795 -172.205 185.125 -171.875 ;
        RECT 184.795 -173.565 185.125 -173.235 ;
        RECT 184.795 -174.925 185.125 -174.595 ;
        RECT 184.795 -176.285 185.125 -175.955 ;
        RECT 184.795 -177.645 185.125 -177.315 ;
        RECT 184.795 -179.005 185.125 -178.675 ;
        RECT 184.795 -180.365 185.125 -180.035 ;
        RECT 184.795 -181.725 185.125 -181.395 ;
        RECT 184.795 -183.085 185.125 -182.755 ;
        RECT 184.795 -184.445 185.125 -184.115 ;
        RECT 184.795 -185.805 185.125 -185.475 ;
        RECT 184.795 -187.165 185.125 -186.835 ;
        RECT 184.795 -188.525 185.125 -188.195 ;
        RECT 184.795 -189.885 185.125 -189.555 ;
        RECT 184.795 -191.245 185.125 -190.915 ;
        RECT 184.795 -192.605 185.125 -192.275 ;
        RECT 184.795 -193.965 185.125 -193.635 ;
        RECT 184.795 -195.325 185.125 -194.995 ;
        RECT 184.795 -196.685 185.125 -196.355 ;
        RECT 184.795 -198.045 185.125 -197.715 ;
        RECT 184.795 -199.405 185.125 -199.075 ;
        RECT 184.795 -200.765 185.125 -200.435 ;
        RECT 184.795 -202.125 185.125 -201.795 ;
        RECT 184.795 -203.485 185.125 -203.155 ;
        RECT 184.795 -204.845 185.125 -204.515 ;
        RECT 184.795 -206.205 185.125 -205.875 ;
        RECT 184.795 -207.565 185.125 -207.235 ;
        RECT 184.795 -208.925 185.125 -208.595 ;
        RECT 184.795 -210.285 185.125 -209.955 ;
        RECT 184.795 -211.645 185.125 -211.315 ;
        RECT 184.795 -213.005 185.125 -212.675 ;
        RECT 184.795 -214.365 185.125 -214.035 ;
        RECT 184.795 -215.725 185.125 -215.395 ;
        RECT 184.795 -217.085 185.125 -216.755 ;
        RECT 184.795 -218.445 185.125 -218.115 ;
        RECT 184.795 -224.09 185.125 -222.96 ;
        RECT 184.8 -224.205 185.12 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.66 -121.535 185.99 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.155 132.52 186.485 133.65 ;
        RECT 186.155 128.355 186.485 128.685 ;
        RECT 186.155 126.995 186.485 127.325 ;
        RECT 186.155 125.635 186.485 125.965 ;
        RECT 186.155 124.275 186.485 124.605 ;
        RECT 186.16 123.6 186.48 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.155 -123.245 186.485 -122.915 ;
        RECT 186.155 -124.605 186.485 -124.275 ;
        RECT 186.155 -125.965 186.485 -125.635 ;
        RECT 186.155 -127.325 186.485 -126.995 ;
        RECT 186.155 -128.685 186.485 -128.355 ;
        RECT 186.155 -130.045 186.485 -129.715 ;
        RECT 186.155 -131.405 186.485 -131.075 ;
        RECT 186.155 -132.765 186.485 -132.435 ;
        RECT 186.155 -134.125 186.485 -133.795 ;
        RECT 186.155 -135.485 186.485 -135.155 ;
        RECT 186.155 -136.845 186.485 -136.515 ;
        RECT 186.155 -138.205 186.485 -137.875 ;
        RECT 186.155 -139.565 186.485 -139.235 ;
        RECT 186.155 -140.925 186.485 -140.595 ;
        RECT 186.155 -142.285 186.485 -141.955 ;
        RECT 186.155 -143.645 186.485 -143.315 ;
        RECT 186.155 -145.005 186.485 -144.675 ;
        RECT 186.155 -146.365 186.485 -146.035 ;
        RECT 186.155 -147.725 186.485 -147.395 ;
        RECT 186.155 -149.085 186.485 -148.755 ;
        RECT 186.155 -150.445 186.485 -150.115 ;
        RECT 186.155 -151.805 186.485 -151.475 ;
        RECT 186.155 -153.165 186.485 -152.835 ;
        RECT 186.155 -154.525 186.485 -154.195 ;
        RECT 186.155 -155.885 186.485 -155.555 ;
        RECT 186.155 -157.245 186.485 -156.915 ;
        RECT 186.155 -158.605 186.485 -158.275 ;
        RECT 186.155 -159.965 186.485 -159.635 ;
        RECT 186.155 -161.325 186.485 -160.995 ;
        RECT 186.155 -162.685 186.485 -162.355 ;
        RECT 186.155 -164.045 186.485 -163.715 ;
        RECT 186.155 -165.405 186.485 -165.075 ;
        RECT 186.155 -166.765 186.485 -166.435 ;
        RECT 186.155 -168.125 186.485 -167.795 ;
        RECT 186.155 -169.485 186.485 -169.155 ;
        RECT 186.155 -170.845 186.485 -170.515 ;
        RECT 186.155 -172.205 186.485 -171.875 ;
        RECT 186.155 -173.565 186.485 -173.235 ;
        RECT 186.155 -174.925 186.485 -174.595 ;
        RECT 186.155 -176.285 186.485 -175.955 ;
        RECT 186.155 -177.645 186.485 -177.315 ;
        RECT 186.155 -179.005 186.485 -178.675 ;
        RECT 186.155 -180.365 186.485 -180.035 ;
        RECT 186.155 -181.725 186.485 -181.395 ;
        RECT 186.155 -183.085 186.485 -182.755 ;
        RECT 186.155 -184.445 186.485 -184.115 ;
        RECT 186.155 -185.805 186.485 -185.475 ;
        RECT 186.155 -187.165 186.485 -186.835 ;
        RECT 186.155 -188.525 186.485 -188.195 ;
        RECT 186.155 -189.885 186.485 -189.555 ;
        RECT 186.155 -191.245 186.485 -190.915 ;
        RECT 186.155 -192.605 186.485 -192.275 ;
        RECT 186.155 -193.965 186.485 -193.635 ;
        RECT 186.155 -195.325 186.485 -194.995 ;
        RECT 186.155 -196.685 186.485 -196.355 ;
        RECT 186.155 -198.045 186.485 -197.715 ;
        RECT 186.155 -199.405 186.485 -199.075 ;
        RECT 186.155 -200.765 186.485 -200.435 ;
        RECT 186.155 -202.125 186.485 -201.795 ;
        RECT 186.155 -203.485 186.485 -203.155 ;
        RECT 186.155 -204.845 186.485 -204.515 ;
        RECT 186.155 -206.205 186.485 -205.875 ;
        RECT 186.155 -207.565 186.485 -207.235 ;
        RECT 186.155 -208.925 186.485 -208.595 ;
        RECT 186.155 -210.285 186.485 -209.955 ;
        RECT 186.155 -211.645 186.485 -211.315 ;
        RECT 186.155 -213.005 186.485 -212.675 ;
        RECT 186.155 -214.365 186.485 -214.035 ;
        RECT 186.155 -215.725 186.485 -215.395 ;
        RECT 186.155 -217.085 186.485 -216.755 ;
        RECT 186.155 -218.445 186.485 -218.115 ;
        RECT 186.155 -224.09 186.485 -222.96 ;
        RECT 186.16 -224.205 186.48 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 187.515 132.52 187.845 133.65 ;
        RECT 187.515 128.355 187.845 128.685 ;
        RECT 187.515 126.995 187.845 127.325 ;
        RECT 187.515 125.635 187.845 125.965 ;
        RECT 187.515 124.275 187.845 124.605 ;
        RECT 187.52 123.6 187.84 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 187.515 -0.845 187.845 -0.515 ;
        RECT 187.515 -2.205 187.845 -1.875 ;
        RECT 187.515 -3.565 187.845 -3.235 ;
        RECT 187.52 -3.565 187.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.875 132.52 189.205 133.65 ;
        RECT 188.875 128.355 189.205 128.685 ;
        RECT 188.875 126.995 189.205 127.325 ;
        RECT 188.875 125.635 189.205 125.965 ;
        RECT 188.875 124.275 189.205 124.605 ;
        RECT 188.88 123.6 189.2 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.875 -0.845 189.205 -0.515 ;
        RECT 188.875 -2.205 189.205 -1.875 ;
        RECT 188.875 -3.565 189.205 -3.235 ;
        RECT 188.88 -3.565 189.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.235 132.52 190.565 133.65 ;
        RECT 190.235 128.355 190.565 128.685 ;
        RECT 190.235 126.995 190.565 127.325 ;
        RECT 190.235 125.635 190.565 125.965 ;
        RECT 190.235 124.275 190.565 124.605 ;
        RECT 190.24 123.6 190.56 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.235 -0.845 190.565 -0.515 ;
        RECT 190.235 -2.205 190.565 -1.875 ;
        RECT 190.235 -3.565 190.565 -3.235 ;
        RECT 190.24 -3.565 190.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.235 -119.165 190.565 -118.835 ;
        RECT 190.235 -120.525 190.565 -120.195 ;
        RECT 190.235 -121.885 190.565 -121.555 ;
        RECT 190.235 -123.245 190.565 -122.915 ;
        RECT 190.235 -124.605 190.565 -124.275 ;
        RECT 190.235 -125.965 190.565 -125.635 ;
        RECT 190.235 -127.325 190.565 -126.995 ;
        RECT 190.235 -128.685 190.565 -128.355 ;
        RECT 190.235 -130.045 190.565 -129.715 ;
        RECT 190.235 -131.405 190.565 -131.075 ;
        RECT 190.235 -132.765 190.565 -132.435 ;
        RECT 190.235 -134.125 190.565 -133.795 ;
        RECT 190.235 -135.485 190.565 -135.155 ;
        RECT 190.235 -136.845 190.565 -136.515 ;
        RECT 190.235 -138.205 190.565 -137.875 ;
        RECT 190.235 -139.565 190.565 -139.235 ;
        RECT 190.235 -140.925 190.565 -140.595 ;
        RECT 190.235 -142.285 190.565 -141.955 ;
        RECT 190.235 -143.645 190.565 -143.315 ;
        RECT 190.235 -145.005 190.565 -144.675 ;
        RECT 190.235 -146.365 190.565 -146.035 ;
        RECT 190.235 -147.725 190.565 -147.395 ;
        RECT 190.235 -149.085 190.565 -148.755 ;
        RECT 190.235 -150.445 190.565 -150.115 ;
        RECT 190.235 -151.805 190.565 -151.475 ;
        RECT 190.235 -153.165 190.565 -152.835 ;
        RECT 190.235 -154.525 190.565 -154.195 ;
        RECT 190.235 -155.885 190.565 -155.555 ;
        RECT 190.235 -157.245 190.565 -156.915 ;
        RECT 190.235 -158.605 190.565 -158.275 ;
        RECT 190.235 -159.965 190.565 -159.635 ;
        RECT 190.235 -161.325 190.565 -160.995 ;
        RECT 190.235 -162.685 190.565 -162.355 ;
        RECT 190.235 -164.045 190.565 -163.715 ;
        RECT 190.235 -165.405 190.565 -165.075 ;
        RECT 190.235 -166.765 190.565 -166.435 ;
        RECT 190.235 -168.125 190.565 -167.795 ;
        RECT 190.235 -169.485 190.565 -169.155 ;
        RECT 190.235 -170.845 190.565 -170.515 ;
        RECT 190.235 -172.205 190.565 -171.875 ;
        RECT 190.235 -173.565 190.565 -173.235 ;
        RECT 190.235 -174.925 190.565 -174.595 ;
        RECT 190.235 -176.285 190.565 -175.955 ;
        RECT 190.235 -177.645 190.565 -177.315 ;
        RECT 190.235 -179.005 190.565 -178.675 ;
        RECT 190.235 -180.365 190.565 -180.035 ;
        RECT 190.235 -181.725 190.565 -181.395 ;
        RECT 190.235 -183.085 190.565 -182.755 ;
        RECT 190.235 -184.445 190.565 -184.115 ;
        RECT 190.235 -185.805 190.565 -185.475 ;
        RECT 190.235 -187.165 190.565 -186.835 ;
        RECT 190.235 -188.525 190.565 -188.195 ;
        RECT 190.235 -189.885 190.565 -189.555 ;
        RECT 190.235 -191.245 190.565 -190.915 ;
        RECT 190.235 -192.605 190.565 -192.275 ;
        RECT 190.235 -193.965 190.565 -193.635 ;
        RECT 190.235 -195.325 190.565 -194.995 ;
        RECT 190.235 -196.685 190.565 -196.355 ;
        RECT 190.235 -198.045 190.565 -197.715 ;
        RECT 190.235 -199.405 190.565 -199.075 ;
        RECT 190.235 -200.765 190.565 -200.435 ;
        RECT 190.235 -202.125 190.565 -201.795 ;
        RECT 190.235 -203.485 190.565 -203.155 ;
        RECT 190.235 -204.845 190.565 -204.515 ;
        RECT 190.235 -206.205 190.565 -205.875 ;
        RECT 190.235 -207.565 190.565 -207.235 ;
        RECT 190.235 -208.925 190.565 -208.595 ;
        RECT 190.235 -210.285 190.565 -209.955 ;
        RECT 190.235 -211.645 190.565 -211.315 ;
        RECT 190.235 -213.005 190.565 -212.675 ;
        RECT 190.235 -214.365 190.565 -214.035 ;
        RECT 190.235 -215.725 190.565 -215.395 ;
        RECT 190.235 -217.085 190.565 -216.755 ;
        RECT 190.235 -218.445 190.565 -218.115 ;
        RECT 190.235 -224.09 190.565 -222.96 ;
        RECT 190.24 -224.205 190.56 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 191.595 132.52 191.925 133.65 ;
        RECT 191.595 128.355 191.925 128.685 ;
        RECT 191.595 126.995 191.925 127.325 ;
        RECT 191.595 125.635 191.925 125.965 ;
        RECT 191.595 124.275 191.925 124.605 ;
        RECT 191.6 123.6 191.92 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 191.595 -206.205 191.925 -205.875 ;
        RECT 191.595 -207.565 191.925 -207.235 ;
        RECT 191.595 -208.925 191.925 -208.595 ;
        RECT 191.595 -210.285 191.925 -209.955 ;
        RECT 191.595 -211.645 191.925 -211.315 ;
        RECT 191.595 -213.005 191.925 -212.675 ;
        RECT 191.595 -214.365 191.925 -214.035 ;
        RECT 191.595 -215.725 191.925 -215.395 ;
        RECT 191.595 -217.085 191.925 -216.755 ;
        RECT 191.595 -218.445 191.925 -218.115 ;
        RECT 191.595 -224.09 191.925 -222.96 ;
        RECT 191.6 -224.205 191.92 -122.24 ;
        RECT 191.595 -123.245 191.925 -122.915 ;
        RECT 191.595 -124.605 191.925 -124.275 ;
        RECT 191.595 -125.965 191.925 -125.635 ;
        RECT 191.595 -127.325 191.925 -126.995 ;
        RECT 191.595 -128.685 191.925 -128.355 ;
        RECT 191.595 -130.045 191.925 -129.715 ;
        RECT 191.595 -131.405 191.925 -131.075 ;
        RECT 191.595 -132.765 191.925 -132.435 ;
        RECT 191.595 -134.125 191.925 -133.795 ;
        RECT 191.595 -135.485 191.925 -135.155 ;
        RECT 191.595 -136.845 191.925 -136.515 ;
        RECT 191.595 -138.205 191.925 -137.875 ;
        RECT 191.595 -139.565 191.925 -139.235 ;
        RECT 191.595 -140.925 191.925 -140.595 ;
        RECT 191.595 -142.285 191.925 -141.955 ;
        RECT 191.595 -143.645 191.925 -143.315 ;
        RECT 191.595 -145.005 191.925 -144.675 ;
        RECT 191.595 -146.365 191.925 -146.035 ;
        RECT 191.595 -147.725 191.925 -147.395 ;
        RECT 191.595 -149.085 191.925 -148.755 ;
        RECT 191.595 -150.445 191.925 -150.115 ;
        RECT 191.595 -151.805 191.925 -151.475 ;
        RECT 191.595 -153.165 191.925 -152.835 ;
        RECT 191.595 -154.525 191.925 -154.195 ;
        RECT 191.595 -155.885 191.925 -155.555 ;
        RECT 191.595 -157.245 191.925 -156.915 ;
        RECT 191.595 -158.605 191.925 -158.275 ;
        RECT 191.595 -159.965 191.925 -159.635 ;
        RECT 191.595 -161.325 191.925 -160.995 ;
        RECT 191.595 -162.685 191.925 -162.355 ;
        RECT 191.595 -164.045 191.925 -163.715 ;
        RECT 191.595 -165.405 191.925 -165.075 ;
        RECT 191.595 -166.765 191.925 -166.435 ;
        RECT 191.595 -168.125 191.925 -167.795 ;
        RECT 191.595 -169.485 191.925 -169.155 ;
        RECT 191.595 -170.845 191.925 -170.515 ;
        RECT 191.595 -172.205 191.925 -171.875 ;
        RECT 191.595 -173.565 191.925 -173.235 ;
        RECT 191.595 -174.925 191.925 -174.595 ;
        RECT 191.595 -176.285 191.925 -175.955 ;
        RECT 191.595 -177.645 191.925 -177.315 ;
        RECT 191.595 -179.005 191.925 -178.675 ;
        RECT 191.595 -180.365 191.925 -180.035 ;
        RECT 191.595 -181.725 191.925 -181.395 ;
        RECT 191.595 -183.085 191.925 -182.755 ;
        RECT 191.595 -184.445 191.925 -184.115 ;
        RECT 191.595 -185.805 191.925 -185.475 ;
        RECT 191.595 -187.165 191.925 -186.835 ;
        RECT 191.595 -188.525 191.925 -188.195 ;
        RECT 191.595 -189.885 191.925 -189.555 ;
        RECT 191.595 -191.245 191.925 -190.915 ;
        RECT 191.595 -192.605 191.925 -192.275 ;
        RECT 191.595 -193.965 191.925 -193.635 ;
        RECT 191.595 -195.325 191.925 -194.995 ;
        RECT 191.595 -196.685 191.925 -196.355 ;
        RECT 191.595 -198.045 191.925 -197.715 ;
        RECT 191.595 -199.405 191.925 -199.075 ;
        RECT 191.595 -200.765 191.925 -200.435 ;
        RECT 191.595 -202.125 191.925 -201.795 ;
        RECT 191.595 -203.485 191.925 -203.155 ;
        RECT 191.595 -204.845 191.925 -204.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.86 -121.535 137.19 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.195 132.52 137.525 133.65 ;
        RECT 137.195 128.355 137.525 128.685 ;
        RECT 137.195 126.995 137.525 127.325 ;
        RECT 137.195 125.635 137.525 125.965 ;
        RECT 137.195 124.275 137.525 124.605 ;
        RECT 137.2 123.6 137.52 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.195 -123.245 137.525 -122.915 ;
        RECT 137.195 -124.605 137.525 -124.275 ;
        RECT 137.195 -125.965 137.525 -125.635 ;
        RECT 137.195 -127.325 137.525 -126.995 ;
        RECT 137.195 -128.685 137.525 -128.355 ;
        RECT 137.195 -130.045 137.525 -129.715 ;
        RECT 137.195 -131.405 137.525 -131.075 ;
        RECT 137.195 -132.765 137.525 -132.435 ;
        RECT 137.195 -134.125 137.525 -133.795 ;
        RECT 137.195 -135.485 137.525 -135.155 ;
        RECT 137.195 -136.845 137.525 -136.515 ;
        RECT 137.195 -138.205 137.525 -137.875 ;
        RECT 137.195 -139.565 137.525 -139.235 ;
        RECT 137.195 -140.925 137.525 -140.595 ;
        RECT 137.195 -142.285 137.525 -141.955 ;
        RECT 137.195 -143.645 137.525 -143.315 ;
        RECT 137.195 -145.005 137.525 -144.675 ;
        RECT 137.195 -146.365 137.525 -146.035 ;
        RECT 137.195 -147.725 137.525 -147.395 ;
        RECT 137.195 -149.085 137.525 -148.755 ;
        RECT 137.195 -150.445 137.525 -150.115 ;
        RECT 137.195 -151.805 137.525 -151.475 ;
        RECT 137.195 -153.165 137.525 -152.835 ;
        RECT 137.195 -154.525 137.525 -154.195 ;
        RECT 137.195 -155.885 137.525 -155.555 ;
        RECT 137.195 -157.245 137.525 -156.915 ;
        RECT 137.195 -158.605 137.525 -158.275 ;
        RECT 137.195 -159.965 137.525 -159.635 ;
        RECT 137.195 -161.325 137.525 -160.995 ;
        RECT 137.195 -162.685 137.525 -162.355 ;
        RECT 137.195 -164.045 137.525 -163.715 ;
        RECT 137.195 -165.405 137.525 -165.075 ;
        RECT 137.195 -166.765 137.525 -166.435 ;
        RECT 137.195 -168.125 137.525 -167.795 ;
        RECT 137.195 -169.485 137.525 -169.155 ;
        RECT 137.195 -170.845 137.525 -170.515 ;
        RECT 137.195 -172.205 137.525 -171.875 ;
        RECT 137.195 -173.565 137.525 -173.235 ;
        RECT 137.195 -174.925 137.525 -174.595 ;
        RECT 137.195 -176.285 137.525 -175.955 ;
        RECT 137.195 -177.645 137.525 -177.315 ;
        RECT 137.195 -179.005 137.525 -178.675 ;
        RECT 137.195 -180.365 137.525 -180.035 ;
        RECT 137.195 -181.725 137.525 -181.395 ;
        RECT 137.195 -183.085 137.525 -182.755 ;
        RECT 137.195 -184.445 137.525 -184.115 ;
        RECT 137.195 -185.805 137.525 -185.475 ;
        RECT 137.195 -187.165 137.525 -186.835 ;
        RECT 137.195 -188.525 137.525 -188.195 ;
        RECT 137.195 -189.885 137.525 -189.555 ;
        RECT 137.195 -191.245 137.525 -190.915 ;
        RECT 137.195 -192.605 137.525 -192.275 ;
        RECT 137.195 -193.965 137.525 -193.635 ;
        RECT 137.195 -195.325 137.525 -194.995 ;
        RECT 137.195 -196.685 137.525 -196.355 ;
        RECT 137.195 -198.045 137.525 -197.715 ;
        RECT 137.195 -199.405 137.525 -199.075 ;
        RECT 137.195 -200.765 137.525 -200.435 ;
        RECT 137.195 -202.125 137.525 -201.795 ;
        RECT 137.195 -203.485 137.525 -203.155 ;
        RECT 137.195 -204.845 137.525 -204.515 ;
        RECT 137.195 -206.205 137.525 -205.875 ;
        RECT 137.195 -207.565 137.525 -207.235 ;
        RECT 137.195 -208.925 137.525 -208.595 ;
        RECT 137.195 -210.285 137.525 -209.955 ;
        RECT 137.195 -211.645 137.525 -211.315 ;
        RECT 137.195 -213.005 137.525 -212.675 ;
        RECT 137.195 -214.365 137.525 -214.035 ;
        RECT 137.195 -215.725 137.525 -215.395 ;
        RECT 137.195 -217.085 137.525 -216.755 ;
        RECT 137.195 -218.445 137.525 -218.115 ;
        RECT 137.195 -224.09 137.525 -222.96 ;
        RECT 137.2 -224.205 137.52 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.555 132.52 138.885 133.65 ;
        RECT 138.555 128.355 138.885 128.685 ;
        RECT 138.555 126.995 138.885 127.325 ;
        RECT 138.555 125.635 138.885 125.965 ;
        RECT 138.555 124.275 138.885 124.605 ;
        RECT 138.56 123.6 138.88 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.555 -0.845 138.885 -0.515 ;
        RECT 138.555 -2.205 138.885 -1.875 ;
        RECT 138.555 -3.565 138.885 -3.235 ;
        RECT 138.56 -3.565 138.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.915 132.52 140.245 133.65 ;
        RECT 139.915 128.355 140.245 128.685 ;
        RECT 139.915 126.995 140.245 127.325 ;
        RECT 139.915 125.635 140.245 125.965 ;
        RECT 139.915 124.275 140.245 124.605 ;
        RECT 139.92 123.6 140.24 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.915 -0.845 140.245 -0.515 ;
        RECT 139.915 -2.205 140.245 -1.875 ;
        RECT 139.915 -3.565 140.245 -3.235 ;
        RECT 139.92 -3.565 140.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.275 132.52 141.605 133.65 ;
        RECT 141.275 128.355 141.605 128.685 ;
        RECT 141.275 126.995 141.605 127.325 ;
        RECT 141.275 125.635 141.605 125.965 ;
        RECT 141.275 124.275 141.605 124.605 ;
        RECT 141.28 123.6 141.6 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.275 -0.845 141.605 -0.515 ;
        RECT 141.275 -2.205 141.605 -1.875 ;
        RECT 141.275 -3.565 141.605 -3.235 ;
        RECT 141.28 -3.565 141.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.275 -119.165 141.605 -118.835 ;
        RECT 141.275 -120.525 141.605 -120.195 ;
        RECT 141.275 -121.885 141.605 -121.555 ;
        RECT 141.275 -123.245 141.605 -122.915 ;
        RECT 141.275 -124.605 141.605 -124.275 ;
        RECT 141.275 -125.965 141.605 -125.635 ;
        RECT 141.275 -127.325 141.605 -126.995 ;
        RECT 141.275 -128.685 141.605 -128.355 ;
        RECT 141.275 -130.045 141.605 -129.715 ;
        RECT 141.275 -131.405 141.605 -131.075 ;
        RECT 141.275 -132.765 141.605 -132.435 ;
        RECT 141.275 -134.125 141.605 -133.795 ;
        RECT 141.275 -135.485 141.605 -135.155 ;
        RECT 141.275 -136.845 141.605 -136.515 ;
        RECT 141.275 -138.205 141.605 -137.875 ;
        RECT 141.275 -139.565 141.605 -139.235 ;
        RECT 141.275 -140.925 141.605 -140.595 ;
        RECT 141.275 -142.285 141.605 -141.955 ;
        RECT 141.275 -143.645 141.605 -143.315 ;
        RECT 141.275 -145.005 141.605 -144.675 ;
        RECT 141.275 -146.365 141.605 -146.035 ;
        RECT 141.275 -147.725 141.605 -147.395 ;
        RECT 141.275 -149.085 141.605 -148.755 ;
        RECT 141.275 -150.445 141.605 -150.115 ;
        RECT 141.275 -151.805 141.605 -151.475 ;
        RECT 141.275 -153.165 141.605 -152.835 ;
        RECT 141.275 -154.525 141.605 -154.195 ;
        RECT 141.275 -155.885 141.605 -155.555 ;
        RECT 141.275 -157.245 141.605 -156.915 ;
        RECT 141.275 -158.605 141.605 -158.275 ;
        RECT 141.275 -159.965 141.605 -159.635 ;
        RECT 141.275 -161.325 141.605 -160.995 ;
        RECT 141.275 -162.685 141.605 -162.355 ;
        RECT 141.275 -164.045 141.605 -163.715 ;
        RECT 141.275 -165.405 141.605 -165.075 ;
        RECT 141.275 -166.765 141.605 -166.435 ;
        RECT 141.275 -168.125 141.605 -167.795 ;
        RECT 141.275 -169.485 141.605 -169.155 ;
        RECT 141.275 -170.845 141.605 -170.515 ;
        RECT 141.275 -172.205 141.605 -171.875 ;
        RECT 141.275 -173.565 141.605 -173.235 ;
        RECT 141.275 -174.925 141.605 -174.595 ;
        RECT 141.275 -176.285 141.605 -175.955 ;
        RECT 141.275 -177.645 141.605 -177.315 ;
        RECT 141.275 -179.005 141.605 -178.675 ;
        RECT 141.275 -180.365 141.605 -180.035 ;
        RECT 141.275 -181.725 141.605 -181.395 ;
        RECT 141.275 -183.085 141.605 -182.755 ;
        RECT 141.275 -184.445 141.605 -184.115 ;
        RECT 141.275 -185.805 141.605 -185.475 ;
        RECT 141.275 -187.165 141.605 -186.835 ;
        RECT 141.275 -188.525 141.605 -188.195 ;
        RECT 141.275 -189.885 141.605 -189.555 ;
        RECT 141.275 -191.245 141.605 -190.915 ;
        RECT 141.275 -192.605 141.605 -192.275 ;
        RECT 141.275 -193.965 141.605 -193.635 ;
        RECT 141.275 -195.325 141.605 -194.995 ;
        RECT 141.275 -196.685 141.605 -196.355 ;
        RECT 141.275 -198.045 141.605 -197.715 ;
        RECT 141.275 -199.405 141.605 -199.075 ;
        RECT 141.275 -200.765 141.605 -200.435 ;
        RECT 141.275 -202.125 141.605 -201.795 ;
        RECT 141.275 -203.485 141.605 -203.155 ;
        RECT 141.275 -204.845 141.605 -204.515 ;
        RECT 141.275 -206.205 141.605 -205.875 ;
        RECT 141.275 -207.565 141.605 -207.235 ;
        RECT 141.275 -208.925 141.605 -208.595 ;
        RECT 141.275 -210.285 141.605 -209.955 ;
        RECT 141.275 -211.645 141.605 -211.315 ;
        RECT 141.275 -213.005 141.605 -212.675 ;
        RECT 141.275 -214.365 141.605 -214.035 ;
        RECT 141.275 -215.725 141.605 -215.395 ;
        RECT 141.275 -217.085 141.605 -216.755 ;
        RECT 141.275 -218.445 141.605 -218.115 ;
        RECT 141.275 -224.09 141.605 -222.96 ;
        RECT 141.28 -224.205 141.6 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.635 132.52 142.965 133.65 ;
        RECT 142.635 128.355 142.965 128.685 ;
        RECT 142.635 126.995 142.965 127.325 ;
        RECT 142.635 125.635 142.965 125.965 ;
        RECT 142.635 124.275 142.965 124.605 ;
        RECT 142.64 123.6 142.96 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.635 -123.245 142.965 -122.915 ;
        RECT 142.635 -124.605 142.965 -124.275 ;
        RECT 142.635 -125.965 142.965 -125.635 ;
        RECT 142.635 -127.325 142.965 -126.995 ;
        RECT 142.635 -128.685 142.965 -128.355 ;
        RECT 142.635 -130.045 142.965 -129.715 ;
        RECT 142.635 -131.405 142.965 -131.075 ;
        RECT 142.635 -132.765 142.965 -132.435 ;
        RECT 142.635 -134.125 142.965 -133.795 ;
        RECT 142.635 -135.485 142.965 -135.155 ;
        RECT 142.635 -136.845 142.965 -136.515 ;
        RECT 142.635 -138.205 142.965 -137.875 ;
        RECT 142.635 -139.565 142.965 -139.235 ;
        RECT 142.635 -140.925 142.965 -140.595 ;
        RECT 142.635 -142.285 142.965 -141.955 ;
        RECT 142.635 -143.645 142.965 -143.315 ;
        RECT 142.635 -145.005 142.965 -144.675 ;
        RECT 142.635 -146.365 142.965 -146.035 ;
        RECT 142.635 -147.725 142.965 -147.395 ;
        RECT 142.635 -149.085 142.965 -148.755 ;
        RECT 142.635 -150.445 142.965 -150.115 ;
        RECT 142.635 -151.805 142.965 -151.475 ;
        RECT 142.635 -153.165 142.965 -152.835 ;
        RECT 142.635 -154.525 142.965 -154.195 ;
        RECT 142.635 -155.885 142.965 -155.555 ;
        RECT 142.635 -157.245 142.965 -156.915 ;
        RECT 142.635 -158.605 142.965 -158.275 ;
        RECT 142.635 -159.965 142.965 -159.635 ;
        RECT 142.635 -161.325 142.965 -160.995 ;
        RECT 142.635 -162.685 142.965 -162.355 ;
        RECT 142.635 -164.045 142.965 -163.715 ;
        RECT 142.635 -165.405 142.965 -165.075 ;
        RECT 142.635 -166.765 142.965 -166.435 ;
        RECT 142.635 -168.125 142.965 -167.795 ;
        RECT 142.635 -169.485 142.965 -169.155 ;
        RECT 142.635 -170.845 142.965 -170.515 ;
        RECT 142.635 -172.205 142.965 -171.875 ;
        RECT 142.635 -173.565 142.965 -173.235 ;
        RECT 142.635 -174.925 142.965 -174.595 ;
        RECT 142.635 -176.285 142.965 -175.955 ;
        RECT 142.635 -177.645 142.965 -177.315 ;
        RECT 142.635 -179.005 142.965 -178.675 ;
        RECT 142.635 -180.365 142.965 -180.035 ;
        RECT 142.635 -181.725 142.965 -181.395 ;
        RECT 142.635 -183.085 142.965 -182.755 ;
        RECT 142.635 -184.445 142.965 -184.115 ;
        RECT 142.635 -185.805 142.965 -185.475 ;
        RECT 142.635 -187.165 142.965 -186.835 ;
        RECT 142.635 -188.525 142.965 -188.195 ;
        RECT 142.635 -189.885 142.965 -189.555 ;
        RECT 142.635 -191.245 142.965 -190.915 ;
        RECT 142.635 -192.605 142.965 -192.275 ;
        RECT 142.635 -193.965 142.965 -193.635 ;
        RECT 142.635 -195.325 142.965 -194.995 ;
        RECT 142.635 -196.685 142.965 -196.355 ;
        RECT 142.635 -198.045 142.965 -197.715 ;
        RECT 142.635 -199.405 142.965 -199.075 ;
        RECT 142.635 -200.765 142.965 -200.435 ;
        RECT 142.635 -202.125 142.965 -201.795 ;
        RECT 142.635 -203.485 142.965 -203.155 ;
        RECT 142.635 -204.845 142.965 -204.515 ;
        RECT 142.635 -206.205 142.965 -205.875 ;
        RECT 142.635 -207.565 142.965 -207.235 ;
        RECT 142.635 -208.925 142.965 -208.595 ;
        RECT 142.635 -210.285 142.965 -209.955 ;
        RECT 142.635 -211.645 142.965 -211.315 ;
        RECT 142.635 -213.005 142.965 -212.675 ;
        RECT 142.635 -214.365 142.965 -214.035 ;
        RECT 142.635 -215.725 142.965 -215.395 ;
        RECT 142.635 -217.085 142.965 -216.755 ;
        RECT 142.635 -218.445 142.965 -218.115 ;
        RECT 142.635 -224.09 142.965 -222.96 ;
        RECT 142.64 -224.205 142.96 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.96 -121.535 143.29 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.995 132.52 144.325 133.65 ;
        RECT 143.995 128.355 144.325 128.685 ;
        RECT 143.995 126.995 144.325 127.325 ;
        RECT 143.995 125.635 144.325 125.965 ;
        RECT 143.995 124.275 144.325 124.605 ;
        RECT 144 123.6 144.32 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.355 132.52 145.685 133.65 ;
        RECT 145.355 128.355 145.685 128.685 ;
        RECT 145.355 126.995 145.685 127.325 ;
        RECT 145.355 125.635 145.685 125.965 ;
        RECT 145.355 124.275 145.685 124.605 ;
        RECT 145.36 123.6 145.68 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.355 -0.845 145.685 -0.515 ;
        RECT 145.355 -2.205 145.685 -1.875 ;
        RECT 145.355 -3.565 145.685 -3.235 ;
        RECT 145.36 -3.565 145.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.715 132.52 147.045 133.65 ;
        RECT 146.715 128.355 147.045 128.685 ;
        RECT 146.715 126.995 147.045 127.325 ;
        RECT 146.715 125.635 147.045 125.965 ;
        RECT 146.715 124.275 147.045 124.605 ;
        RECT 146.72 123.6 147.04 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.715 -0.845 147.045 -0.515 ;
        RECT 146.715 -2.205 147.045 -1.875 ;
        RECT 146.715 -3.565 147.045 -3.235 ;
        RECT 146.72 -3.565 147.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.715 -119.165 147.045 -118.835 ;
        RECT 146.715 -120.525 147.045 -120.195 ;
        RECT 146.715 -121.885 147.045 -121.555 ;
        RECT 146.715 -123.245 147.045 -122.915 ;
        RECT 146.715 -124.605 147.045 -124.275 ;
        RECT 146.715 -125.965 147.045 -125.635 ;
        RECT 146.715 -127.325 147.045 -126.995 ;
        RECT 146.715 -128.685 147.045 -128.355 ;
        RECT 146.715 -130.045 147.045 -129.715 ;
        RECT 146.715 -131.405 147.045 -131.075 ;
        RECT 146.715 -132.765 147.045 -132.435 ;
        RECT 146.715 -134.125 147.045 -133.795 ;
        RECT 146.715 -135.485 147.045 -135.155 ;
        RECT 146.715 -136.845 147.045 -136.515 ;
        RECT 146.715 -138.205 147.045 -137.875 ;
        RECT 146.715 -139.565 147.045 -139.235 ;
        RECT 146.715 -140.925 147.045 -140.595 ;
        RECT 146.715 -142.285 147.045 -141.955 ;
        RECT 146.715 -143.645 147.045 -143.315 ;
        RECT 146.715 -145.005 147.045 -144.675 ;
        RECT 146.715 -146.365 147.045 -146.035 ;
        RECT 146.715 -147.725 147.045 -147.395 ;
        RECT 146.715 -149.085 147.045 -148.755 ;
        RECT 146.715 -150.445 147.045 -150.115 ;
        RECT 146.715 -151.805 147.045 -151.475 ;
        RECT 146.715 -153.165 147.045 -152.835 ;
        RECT 146.715 -154.525 147.045 -154.195 ;
        RECT 146.715 -155.885 147.045 -155.555 ;
        RECT 146.715 -157.245 147.045 -156.915 ;
        RECT 146.715 -158.605 147.045 -158.275 ;
        RECT 146.715 -159.965 147.045 -159.635 ;
        RECT 146.715 -161.325 147.045 -160.995 ;
        RECT 146.715 -162.685 147.045 -162.355 ;
        RECT 146.715 -164.045 147.045 -163.715 ;
        RECT 146.715 -165.405 147.045 -165.075 ;
        RECT 146.715 -166.765 147.045 -166.435 ;
        RECT 146.715 -168.125 147.045 -167.795 ;
        RECT 146.715 -169.485 147.045 -169.155 ;
        RECT 146.715 -170.845 147.045 -170.515 ;
        RECT 146.715 -172.205 147.045 -171.875 ;
        RECT 146.715 -173.565 147.045 -173.235 ;
        RECT 146.715 -174.925 147.045 -174.595 ;
        RECT 146.715 -176.285 147.045 -175.955 ;
        RECT 146.715 -177.645 147.045 -177.315 ;
        RECT 146.715 -179.005 147.045 -178.675 ;
        RECT 146.715 -180.365 147.045 -180.035 ;
        RECT 146.715 -181.725 147.045 -181.395 ;
        RECT 146.715 -183.085 147.045 -182.755 ;
        RECT 146.715 -184.445 147.045 -184.115 ;
        RECT 146.715 -185.805 147.045 -185.475 ;
        RECT 146.715 -187.165 147.045 -186.835 ;
        RECT 146.715 -188.525 147.045 -188.195 ;
        RECT 146.715 -189.885 147.045 -189.555 ;
        RECT 146.715 -191.245 147.045 -190.915 ;
        RECT 146.715 -192.605 147.045 -192.275 ;
        RECT 146.715 -193.965 147.045 -193.635 ;
        RECT 146.715 -195.325 147.045 -194.995 ;
        RECT 146.715 -196.685 147.045 -196.355 ;
        RECT 146.715 -198.045 147.045 -197.715 ;
        RECT 146.715 -199.405 147.045 -199.075 ;
        RECT 146.715 -200.765 147.045 -200.435 ;
        RECT 146.715 -202.125 147.045 -201.795 ;
        RECT 146.715 -203.485 147.045 -203.155 ;
        RECT 146.715 -204.845 147.045 -204.515 ;
        RECT 146.715 -206.205 147.045 -205.875 ;
        RECT 146.715 -207.565 147.045 -207.235 ;
        RECT 146.715 -208.925 147.045 -208.595 ;
        RECT 146.715 -210.285 147.045 -209.955 ;
        RECT 146.715 -211.645 147.045 -211.315 ;
        RECT 146.715 -213.005 147.045 -212.675 ;
        RECT 146.715 -214.365 147.045 -214.035 ;
        RECT 146.715 -215.725 147.045 -215.395 ;
        RECT 146.715 -217.085 147.045 -216.755 ;
        RECT 146.715 -218.445 147.045 -218.115 ;
        RECT 146.715 -224.09 147.045 -222.96 ;
        RECT 146.72 -224.205 147.04 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.075 132.52 148.405 133.65 ;
        RECT 148.075 128.355 148.405 128.685 ;
        RECT 148.075 126.995 148.405 127.325 ;
        RECT 148.075 125.635 148.405 125.965 ;
        RECT 148.075 124.275 148.405 124.605 ;
        RECT 148.08 123.6 148.4 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.075 -0.845 148.405 -0.515 ;
        RECT 148.075 -2.205 148.405 -1.875 ;
        RECT 148.075 -3.565 148.405 -3.235 ;
        RECT 148.08 -3.565 148.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.075 -119.165 148.405 -118.835 ;
        RECT 148.075 -120.525 148.405 -120.195 ;
        RECT 148.075 -121.885 148.405 -121.555 ;
        RECT 148.075 -123.245 148.405 -122.915 ;
        RECT 148.075 -124.605 148.405 -124.275 ;
        RECT 148.075 -125.965 148.405 -125.635 ;
        RECT 148.075 -127.325 148.405 -126.995 ;
        RECT 148.075 -128.685 148.405 -128.355 ;
        RECT 148.075 -130.045 148.405 -129.715 ;
        RECT 148.075 -131.405 148.405 -131.075 ;
        RECT 148.075 -132.765 148.405 -132.435 ;
        RECT 148.075 -134.125 148.405 -133.795 ;
        RECT 148.075 -135.485 148.405 -135.155 ;
        RECT 148.075 -136.845 148.405 -136.515 ;
        RECT 148.075 -138.205 148.405 -137.875 ;
        RECT 148.075 -139.565 148.405 -139.235 ;
        RECT 148.075 -140.925 148.405 -140.595 ;
        RECT 148.075 -142.285 148.405 -141.955 ;
        RECT 148.075 -143.645 148.405 -143.315 ;
        RECT 148.075 -145.005 148.405 -144.675 ;
        RECT 148.075 -146.365 148.405 -146.035 ;
        RECT 148.075 -147.725 148.405 -147.395 ;
        RECT 148.075 -149.085 148.405 -148.755 ;
        RECT 148.075 -150.445 148.405 -150.115 ;
        RECT 148.075 -151.805 148.405 -151.475 ;
        RECT 148.075 -153.165 148.405 -152.835 ;
        RECT 148.075 -154.525 148.405 -154.195 ;
        RECT 148.075 -155.885 148.405 -155.555 ;
        RECT 148.075 -157.245 148.405 -156.915 ;
        RECT 148.075 -158.605 148.405 -158.275 ;
        RECT 148.075 -159.965 148.405 -159.635 ;
        RECT 148.075 -161.325 148.405 -160.995 ;
        RECT 148.075 -162.685 148.405 -162.355 ;
        RECT 148.075 -164.045 148.405 -163.715 ;
        RECT 148.075 -165.405 148.405 -165.075 ;
        RECT 148.075 -166.765 148.405 -166.435 ;
        RECT 148.075 -168.125 148.405 -167.795 ;
        RECT 148.075 -169.485 148.405 -169.155 ;
        RECT 148.075 -170.845 148.405 -170.515 ;
        RECT 148.075 -172.205 148.405 -171.875 ;
        RECT 148.075 -173.565 148.405 -173.235 ;
        RECT 148.075 -174.925 148.405 -174.595 ;
        RECT 148.075 -176.285 148.405 -175.955 ;
        RECT 148.075 -177.645 148.405 -177.315 ;
        RECT 148.075 -179.005 148.405 -178.675 ;
        RECT 148.075 -180.365 148.405 -180.035 ;
        RECT 148.075 -181.725 148.405 -181.395 ;
        RECT 148.075 -183.085 148.405 -182.755 ;
        RECT 148.075 -184.445 148.405 -184.115 ;
        RECT 148.075 -185.805 148.405 -185.475 ;
        RECT 148.075 -187.165 148.405 -186.835 ;
        RECT 148.075 -188.525 148.405 -188.195 ;
        RECT 148.075 -189.885 148.405 -189.555 ;
        RECT 148.075 -191.245 148.405 -190.915 ;
        RECT 148.075 -192.605 148.405 -192.275 ;
        RECT 148.075 -193.965 148.405 -193.635 ;
        RECT 148.075 -195.325 148.405 -194.995 ;
        RECT 148.075 -196.685 148.405 -196.355 ;
        RECT 148.075 -198.045 148.405 -197.715 ;
        RECT 148.075 -199.405 148.405 -199.075 ;
        RECT 148.075 -200.765 148.405 -200.435 ;
        RECT 148.075 -202.125 148.405 -201.795 ;
        RECT 148.075 -203.485 148.405 -203.155 ;
        RECT 148.075 -204.845 148.405 -204.515 ;
        RECT 148.075 -206.205 148.405 -205.875 ;
        RECT 148.075 -207.565 148.405 -207.235 ;
        RECT 148.075 -208.925 148.405 -208.595 ;
        RECT 148.075 -210.285 148.405 -209.955 ;
        RECT 148.075 -211.645 148.405 -211.315 ;
        RECT 148.075 -213.005 148.405 -212.675 ;
        RECT 148.075 -214.365 148.405 -214.035 ;
        RECT 148.075 -215.725 148.405 -215.395 ;
        RECT 148.075 -217.085 148.405 -216.755 ;
        RECT 148.075 -218.445 148.405 -218.115 ;
        RECT 148.075 -224.09 148.405 -222.96 ;
        RECT 148.08 -224.205 148.4 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.06 -121.535 149.39 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.435 132.52 149.765 133.65 ;
        RECT 149.435 128.355 149.765 128.685 ;
        RECT 149.435 126.995 149.765 127.325 ;
        RECT 149.435 125.635 149.765 125.965 ;
        RECT 149.435 124.275 149.765 124.605 ;
        RECT 149.44 123.6 149.76 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.435 -123.245 149.765 -122.915 ;
        RECT 149.435 -124.605 149.765 -124.275 ;
        RECT 149.435 -125.965 149.765 -125.635 ;
        RECT 149.435 -127.325 149.765 -126.995 ;
        RECT 149.435 -128.685 149.765 -128.355 ;
        RECT 149.435 -130.045 149.765 -129.715 ;
        RECT 149.435 -131.405 149.765 -131.075 ;
        RECT 149.435 -132.765 149.765 -132.435 ;
        RECT 149.435 -134.125 149.765 -133.795 ;
        RECT 149.435 -135.485 149.765 -135.155 ;
        RECT 149.435 -136.845 149.765 -136.515 ;
        RECT 149.435 -138.205 149.765 -137.875 ;
        RECT 149.435 -139.565 149.765 -139.235 ;
        RECT 149.435 -140.925 149.765 -140.595 ;
        RECT 149.435 -142.285 149.765 -141.955 ;
        RECT 149.435 -143.645 149.765 -143.315 ;
        RECT 149.435 -145.005 149.765 -144.675 ;
        RECT 149.435 -146.365 149.765 -146.035 ;
        RECT 149.435 -147.725 149.765 -147.395 ;
        RECT 149.435 -149.085 149.765 -148.755 ;
        RECT 149.435 -150.445 149.765 -150.115 ;
        RECT 149.435 -151.805 149.765 -151.475 ;
        RECT 149.435 -153.165 149.765 -152.835 ;
        RECT 149.435 -154.525 149.765 -154.195 ;
        RECT 149.435 -155.885 149.765 -155.555 ;
        RECT 149.435 -157.245 149.765 -156.915 ;
        RECT 149.435 -158.605 149.765 -158.275 ;
        RECT 149.435 -159.965 149.765 -159.635 ;
        RECT 149.435 -161.325 149.765 -160.995 ;
        RECT 149.435 -162.685 149.765 -162.355 ;
        RECT 149.435 -164.045 149.765 -163.715 ;
        RECT 149.435 -165.405 149.765 -165.075 ;
        RECT 149.435 -166.765 149.765 -166.435 ;
        RECT 149.435 -168.125 149.765 -167.795 ;
        RECT 149.435 -169.485 149.765 -169.155 ;
        RECT 149.435 -170.845 149.765 -170.515 ;
        RECT 149.435 -172.205 149.765 -171.875 ;
        RECT 149.435 -173.565 149.765 -173.235 ;
        RECT 149.435 -174.925 149.765 -174.595 ;
        RECT 149.435 -176.285 149.765 -175.955 ;
        RECT 149.435 -177.645 149.765 -177.315 ;
        RECT 149.435 -179.005 149.765 -178.675 ;
        RECT 149.435 -180.365 149.765 -180.035 ;
        RECT 149.435 -181.725 149.765 -181.395 ;
        RECT 149.435 -183.085 149.765 -182.755 ;
        RECT 149.435 -184.445 149.765 -184.115 ;
        RECT 149.435 -185.805 149.765 -185.475 ;
        RECT 149.435 -187.165 149.765 -186.835 ;
        RECT 149.435 -188.525 149.765 -188.195 ;
        RECT 149.435 -189.885 149.765 -189.555 ;
        RECT 149.435 -191.245 149.765 -190.915 ;
        RECT 149.435 -192.605 149.765 -192.275 ;
        RECT 149.435 -193.965 149.765 -193.635 ;
        RECT 149.435 -195.325 149.765 -194.995 ;
        RECT 149.435 -196.685 149.765 -196.355 ;
        RECT 149.435 -198.045 149.765 -197.715 ;
        RECT 149.435 -199.405 149.765 -199.075 ;
        RECT 149.435 -200.765 149.765 -200.435 ;
        RECT 149.435 -202.125 149.765 -201.795 ;
        RECT 149.435 -203.485 149.765 -203.155 ;
        RECT 149.435 -204.845 149.765 -204.515 ;
        RECT 149.435 -206.205 149.765 -205.875 ;
        RECT 149.435 -207.565 149.765 -207.235 ;
        RECT 149.435 -208.925 149.765 -208.595 ;
        RECT 149.435 -210.285 149.765 -209.955 ;
        RECT 149.435 -211.645 149.765 -211.315 ;
        RECT 149.435 -213.005 149.765 -212.675 ;
        RECT 149.435 -214.365 149.765 -214.035 ;
        RECT 149.435 -215.725 149.765 -215.395 ;
        RECT 149.435 -217.085 149.765 -216.755 ;
        RECT 149.435 -218.445 149.765 -218.115 ;
        RECT 149.435 -224.09 149.765 -222.96 ;
        RECT 149.44 -224.205 149.76 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.795 132.52 151.125 133.65 ;
        RECT 150.795 128.355 151.125 128.685 ;
        RECT 150.795 126.995 151.125 127.325 ;
        RECT 150.795 125.635 151.125 125.965 ;
        RECT 150.795 124.275 151.125 124.605 ;
        RECT 150.8 123.6 151.12 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.795 -0.845 151.125 -0.515 ;
        RECT 150.795 -2.205 151.125 -1.875 ;
        RECT 150.795 -3.565 151.125 -3.235 ;
        RECT 150.8 -3.565 151.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.155 132.52 152.485 133.65 ;
        RECT 152.155 128.355 152.485 128.685 ;
        RECT 152.155 126.995 152.485 127.325 ;
        RECT 152.155 125.635 152.485 125.965 ;
        RECT 152.155 124.275 152.485 124.605 ;
        RECT 152.16 123.6 152.48 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.155 -0.845 152.485 -0.515 ;
        RECT 152.155 -2.205 152.485 -1.875 ;
        RECT 152.155 -3.565 152.485 -3.235 ;
        RECT 152.16 -3.565 152.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.515 132.52 153.845 133.65 ;
        RECT 153.515 128.355 153.845 128.685 ;
        RECT 153.515 126.995 153.845 127.325 ;
        RECT 153.515 125.635 153.845 125.965 ;
        RECT 153.515 124.275 153.845 124.605 ;
        RECT 153.52 123.6 153.84 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.515 -0.845 153.845 -0.515 ;
        RECT 153.515 -2.205 153.845 -1.875 ;
        RECT 153.515 -3.565 153.845 -3.235 ;
        RECT 153.52 -3.565 153.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.875 132.52 155.205 133.65 ;
        RECT 154.875 128.355 155.205 128.685 ;
        RECT 154.875 126.995 155.205 127.325 ;
        RECT 154.875 125.635 155.205 125.965 ;
        RECT 154.875 124.275 155.205 124.605 ;
        RECT 154.88 123.6 155.2 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.875 -123.245 155.205 -122.915 ;
        RECT 154.875 -124.605 155.205 -124.275 ;
        RECT 154.875 -125.965 155.205 -125.635 ;
        RECT 154.875 -127.325 155.205 -126.995 ;
        RECT 154.875 -128.685 155.205 -128.355 ;
        RECT 154.875 -130.045 155.205 -129.715 ;
        RECT 154.875 -131.405 155.205 -131.075 ;
        RECT 154.875 -132.765 155.205 -132.435 ;
        RECT 154.875 -134.125 155.205 -133.795 ;
        RECT 154.875 -135.485 155.205 -135.155 ;
        RECT 154.875 -136.845 155.205 -136.515 ;
        RECT 154.875 -138.205 155.205 -137.875 ;
        RECT 154.875 -139.565 155.205 -139.235 ;
        RECT 154.875 -140.925 155.205 -140.595 ;
        RECT 154.875 -142.285 155.205 -141.955 ;
        RECT 154.875 -143.645 155.205 -143.315 ;
        RECT 154.875 -145.005 155.205 -144.675 ;
        RECT 154.875 -146.365 155.205 -146.035 ;
        RECT 154.875 -147.725 155.205 -147.395 ;
        RECT 154.875 -149.085 155.205 -148.755 ;
        RECT 154.875 -150.445 155.205 -150.115 ;
        RECT 154.875 -151.805 155.205 -151.475 ;
        RECT 154.875 -153.165 155.205 -152.835 ;
        RECT 154.875 -154.525 155.205 -154.195 ;
        RECT 154.875 -155.885 155.205 -155.555 ;
        RECT 154.875 -157.245 155.205 -156.915 ;
        RECT 154.875 -158.605 155.205 -158.275 ;
        RECT 154.875 -159.965 155.205 -159.635 ;
        RECT 154.875 -161.325 155.205 -160.995 ;
        RECT 154.875 -162.685 155.205 -162.355 ;
        RECT 154.875 -164.045 155.205 -163.715 ;
        RECT 154.875 -165.405 155.205 -165.075 ;
        RECT 154.875 -166.765 155.205 -166.435 ;
        RECT 154.875 -168.125 155.205 -167.795 ;
        RECT 154.875 -169.485 155.205 -169.155 ;
        RECT 154.875 -170.845 155.205 -170.515 ;
        RECT 154.875 -172.205 155.205 -171.875 ;
        RECT 154.875 -173.565 155.205 -173.235 ;
        RECT 154.875 -174.925 155.205 -174.595 ;
        RECT 154.875 -176.285 155.205 -175.955 ;
        RECT 154.875 -177.645 155.205 -177.315 ;
        RECT 154.875 -179.005 155.205 -178.675 ;
        RECT 154.875 -180.365 155.205 -180.035 ;
        RECT 154.875 -181.725 155.205 -181.395 ;
        RECT 154.875 -183.085 155.205 -182.755 ;
        RECT 154.875 -184.445 155.205 -184.115 ;
        RECT 154.875 -185.805 155.205 -185.475 ;
        RECT 154.875 -187.165 155.205 -186.835 ;
        RECT 154.875 -188.525 155.205 -188.195 ;
        RECT 154.875 -189.885 155.205 -189.555 ;
        RECT 154.875 -191.245 155.205 -190.915 ;
        RECT 154.875 -192.605 155.205 -192.275 ;
        RECT 154.875 -193.965 155.205 -193.635 ;
        RECT 154.875 -195.325 155.205 -194.995 ;
        RECT 154.875 -196.685 155.205 -196.355 ;
        RECT 154.875 -198.045 155.205 -197.715 ;
        RECT 154.875 -199.405 155.205 -199.075 ;
        RECT 154.875 -200.765 155.205 -200.435 ;
        RECT 154.875 -202.125 155.205 -201.795 ;
        RECT 154.875 -203.485 155.205 -203.155 ;
        RECT 154.875 -204.845 155.205 -204.515 ;
        RECT 154.875 -206.205 155.205 -205.875 ;
        RECT 154.875 -207.565 155.205 -207.235 ;
        RECT 154.875 -208.925 155.205 -208.595 ;
        RECT 154.875 -210.285 155.205 -209.955 ;
        RECT 154.875 -211.645 155.205 -211.315 ;
        RECT 154.875 -213.005 155.205 -212.675 ;
        RECT 154.875 -214.365 155.205 -214.035 ;
        RECT 154.875 -215.725 155.205 -215.395 ;
        RECT 154.875 -217.085 155.205 -216.755 ;
        RECT 154.875 -218.445 155.205 -218.115 ;
        RECT 154.875 -224.09 155.205 -222.96 ;
        RECT 154.88 -224.205 155.2 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.16 -121.535 155.49 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.235 132.52 156.565 133.65 ;
        RECT 156.235 128.355 156.565 128.685 ;
        RECT 156.235 126.995 156.565 127.325 ;
        RECT 156.235 125.635 156.565 125.965 ;
        RECT 156.235 124.275 156.565 124.605 ;
        RECT 156.24 123.6 156.56 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 157.595 132.52 157.925 133.65 ;
        RECT 157.595 128.355 157.925 128.685 ;
        RECT 157.595 126.995 157.925 127.325 ;
        RECT 157.595 125.635 157.925 125.965 ;
        RECT 157.595 124.275 157.925 124.605 ;
        RECT 157.6 123.6 157.92 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 157.595 -0.845 157.925 -0.515 ;
        RECT 157.595 -2.205 157.925 -1.875 ;
        RECT 157.595 -3.565 157.925 -3.235 ;
        RECT 157.6 -3.565 157.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.955 132.52 159.285 133.65 ;
        RECT 158.955 128.355 159.285 128.685 ;
        RECT 158.955 126.995 159.285 127.325 ;
        RECT 158.955 125.635 159.285 125.965 ;
        RECT 158.955 124.275 159.285 124.605 ;
        RECT 158.96 123.6 159.28 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.955 -0.845 159.285 -0.515 ;
        RECT 158.955 -2.205 159.285 -1.875 ;
        RECT 158.955 -3.565 159.285 -3.235 ;
        RECT 158.96 -3.565 159.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.955 -119.165 159.285 -118.835 ;
        RECT 158.955 -120.525 159.285 -120.195 ;
        RECT 158.955 -121.885 159.285 -121.555 ;
        RECT 158.955 -123.245 159.285 -122.915 ;
        RECT 158.955 -124.605 159.285 -124.275 ;
        RECT 158.955 -125.965 159.285 -125.635 ;
        RECT 158.955 -127.325 159.285 -126.995 ;
        RECT 158.955 -128.685 159.285 -128.355 ;
        RECT 158.955 -130.045 159.285 -129.715 ;
        RECT 158.955 -131.405 159.285 -131.075 ;
        RECT 158.955 -132.765 159.285 -132.435 ;
        RECT 158.955 -134.125 159.285 -133.795 ;
        RECT 158.955 -135.485 159.285 -135.155 ;
        RECT 158.955 -136.845 159.285 -136.515 ;
        RECT 158.955 -138.205 159.285 -137.875 ;
        RECT 158.955 -139.565 159.285 -139.235 ;
        RECT 158.955 -140.925 159.285 -140.595 ;
        RECT 158.955 -142.285 159.285 -141.955 ;
        RECT 158.955 -143.645 159.285 -143.315 ;
        RECT 158.955 -145.005 159.285 -144.675 ;
        RECT 158.955 -146.365 159.285 -146.035 ;
        RECT 158.955 -147.725 159.285 -147.395 ;
        RECT 158.955 -149.085 159.285 -148.755 ;
        RECT 158.955 -150.445 159.285 -150.115 ;
        RECT 158.955 -151.805 159.285 -151.475 ;
        RECT 158.955 -153.165 159.285 -152.835 ;
        RECT 158.955 -154.525 159.285 -154.195 ;
        RECT 158.955 -155.885 159.285 -155.555 ;
        RECT 158.955 -157.245 159.285 -156.915 ;
        RECT 158.955 -158.605 159.285 -158.275 ;
        RECT 158.955 -159.965 159.285 -159.635 ;
        RECT 158.955 -161.325 159.285 -160.995 ;
        RECT 158.955 -162.685 159.285 -162.355 ;
        RECT 158.955 -164.045 159.285 -163.715 ;
        RECT 158.955 -165.405 159.285 -165.075 ;
        RECT 158.955 -166.765 159.285 -166.435 ;
        RECT 158.955 -168.125 159.285 -167.795 ;
        RECT 158.955 -169.485 159.285 -169.155 ;
        RECT 158.955 -170.845 159.285 -170.515 ;
        RECT 158.955 -172.205 159.285 -171.875 ;
        RECT 158.955 -173.565 159.285 -173.235 ;
        RECT 158.955 -174.925 159.285 -174.595 ;
        RECT 158.955 -176.285 159.285 -175.955 ;
        RECT 158.955 -177.645 159.285 -177.315 ;
        RECT 158.955 -179.005 159.285 -178.675 ;
        RECT 158.955 -180.365 159.285 -180.035 ;
        RECT 158.955 -181.725 159.285 -181.395 ;
        RECT 158.955 -183.085 159.285 -182.755 ;
        RECT 158.955 -184.445 159.285 -184.115 ;
        RECT 158.955 -185.805 159.285 -185.475 ;
        RECT 158.955 -187.165 159.285 -186.835 ;
        RECT 158.955 -188.525 159.285 -188.195 ;
        RECT 158.955 -189.885 159.285 -189.555 ;
        RECT 158.955 -191.245 159.285 -190.915 ;
        RECT 158.955 -192.605 159.285 -192.275 ;
        RECT 158.955 -193.965 159.285 -193.635 ;
        RECT 158.955 -195.325 159.285 -194.995 ;
        RECT 158.955 -196.685 159.285 -196.355 ;
        RECT 158.955 -198.045 159.285 -197.715 ;
        RECT 158.955 -199.405 159.285 -199.075 ;
        RECT 158.955 -200.765 159.285 -200.435 ;
        RECT 158.955 -202.125 159.285 -201.795 ;
        RECT 158.955 -203.485 159.285 -203.155 ;
        RECT 158.955 -204.845 159.285 -204.515 ;
        RECT 158.955 -206.205 159.285 -205.875 ;
        RECT 158.955 -207.565 159.285 -207.235 ;
        RECT 158.955 -208.925 159.285 -208.595 ;
        RECT 158.955 -210.285 159.285 -209.955 ;
        RECT 158.955 -211.645 159.285 -211.315 ;
        RECT 158.955 -213.005 159.285 -212.675 ;
        RECT 158.955 -214.365 159.285 -214.035 ;
        RECT 158.955 -215.725 159.285 -215.395 ;
        RECT 158.955 -217.085 159.285 -216.755 ;
        RECT 158.955 -218.445 159.285 -218.115 ;
        RECT 158.955 -224.09 159.285 -222.96 ;
        RECT 158.96 -224.205 159.28 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.315 132.52 160.645 133.65 ;
        RECT 160.315 128.355 160.645 128.685 ;
        RECT 160.315 126.995 160.645 127.325 ;
        RECT 160.315 125.635 160.645 125.965 ;
        RECT 160.315 124.275 160.645 124.605 ;
        RECT 160.32 123.6 160.64 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.315 -0.845 160.645 -0.515 ;
        RECT 160.315 -2.205 160.645 -1.875 ;
        RECT 160.315 -3.565 160.645 -3.235 ;
        RECT 160.32 -3.565 160.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.315 -119.165 160.645 -118.835 ;
        RECT 160.315 -120.525 160.645 -120.195 ;
        RECT 160.315 -121.885 160.645 -121.555 ;
        RECT 160.315 -123.245 160.645 -122.915 ;
        RECT 160.315 -124.605 160.645 -124.275 ;
        RECT 160.315 -125.965 160.645 -125.635 ;
        RECT 160.315 -127.325 160.645 -126.995 ;
        RECT 160.315 -128.685 160.645 -128.355 ;
        RECT 160.315 -130.045 160.645 -129.715 ;
        RECT 160.315 -131.405 160.645 -131.075 ;
        RECT 160.315 -132.765 160.645 -132.435 ;
        RECT 160.315 -134.125 160.645 -133.795 ;
        RECT 160.315 -135.485 160.645 -135.155 ;
        RECT 160.315 -136.845 160.645 -136.515 ;
        RECT 160.315 -138.205 160.645 -137.875 ;
        RECT 160.315 -139.565 160.645 -139.235 ;
        RECT 160.315 -140.925 160.645 -140.595 ;
        RECT 160.315 -142.285 160.645 -141.955 ;
        RECT 160.315 -143.645 160.645 -143.315 ;
        RECT 160.315 -145.005 160.645 -144.675 ;
        RECT 160.315 -146.365 160.645 -146.035 ;
        RECT 160.315 -147.725 160.645 -147.395 ;
        RECT 160.315 -149.085 160.645 -148.755 ;
        RECT 160.315 -150.445 160.645 -150.115 ;
        RECT 160.315 -151.805 160.645 -151.475 ;
        RECT 160.315 -153.165 160.645 -152.835 ;
        RECT 160.315 -154.525 160.645 -154.195 ;
        RECT 160.315 -155.885 160.645 -155.555 ;
        RECT 160.315 -157.245 160.645 -156.915 ;
        RECT 160.315 -158.605 160.645 -158.275 ;
        RECT 160.315 -159.965 160.645 -159.635 ;
        RECT 160.315 -161.325 160.645 -160.995 ;
        RECT 160.315 -162.685 160.645 -162.355 ;
        RECT 160.315 -164.045 160.645 -163.715 ;
        RECT 160.315 -165.405 160.645 -165.075 ;
        RECT 160.315 -166.765 160.645 -166.435 ;
        RECT 160.315 -168.125 160.645 -167.795 ;
        RECT 160.315 -169.485 160.645 -169.155 ;
        RECT 160.315 -170.845 160.645 -170.515 ;
        RECT 160.315 -172.205 160.645 -171.875 ;
        RECT 160.315 -173.565 160.645 -173.235 ;
        RECT 160.315 -174.925 160.645 -174.595 ;
        RECT 160.315 -176.285 160.645 -175.955 ;
        RECT 160.315 -177.645 160.645 -177.315 ;
        RECT 160.315 -179.005 160.645 -178.675 ;
        RECT 160.315 -180.365 160.645 -180.035 ;
        RECT 160.315 -181.725 160.645 -181.395 ;
        RECT 160.315 -183.085 160.645 -182.755 ;
        RECT 160.315 -184.445 160.645 -184.115 ;
        RECT 160.315 -185.805 160.645 -185.475 ;
        RECT 160.315 -187.165 160.645 -186.835 ;
        RECT 160.315 -188.525 160.645 -188.195 ;
        RECT 160.315 -189.885 160.645 -189.555 ;
        RECT 160.315 -191.245 160.645 -190.915 ;
        RECT 160.315 -192.605 160.645 -192.275 ;
        RECT 160.315 -193.965 160.645 -193.635 ;
        RECT 160.315 -195.325 160.645 -194.995 ;
        RECT 160.315 -196.685 160.645 -196.355 ;
        RECT 160.315 -198.045 160.645 -197.715 ;
        RECT 160.315 -199.405 160.645 -199.075 ;
        RECT 160.315 -200.765 160.645 -200.435 ;
        RECT 160.315 -202.125 160.645 -201.795 ;
        RECT 160.315 -203.485 160.645 -203.155 ;
        RECT 160.315 -204.845 160.645 -204.515 ;
        RECT 160.315 -206.205 160.645 -205.875 ;
        RECT 160.315 -207.565 160.645 -207.235 ;
        RECT 160.315 -208.925 160.645 -208.595 ;
        RECT 160.315 -210.285 160.645 -209.955 ;
        RECT 160.315 -211.645 160.645 -211.315 ;
        RECT 160.315 -213.005 160.645 -212.675 ;
        RECT 160.315 -214.365 160.645 -214.035 ;
        RECT 160.315 -215.725 160.645 -215.395 ;
        RECT 160.315 -217.085 160.645 -216.755 ;
        RECT 160.315 -218.445 160.645 -218.115 ;
        RECT 160.315 -224.09 160.645 -222.96 ;
        RECT 160.32 -224.205 160.64 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.26 -121.535 161.59 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.675 132.52 162.005 133.65 ;
        RECT 161.675 128.355 162.005 128.685 ;
        RECT 161.675 126.995 162.005 127.325 ;
        RECT 161.675 125.635 162.005 125.965 ;
        RECT 161.675 124.275 162.005 124.605 ;
        RECT 161.68 123.6 162 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.675 -123.245 162.005 -122.915 ;
        RECT 161.675 -124.605 162.005 -124.275 ;
        RECT 161.675 -125.965 162.005 -125.635 ;
        RECT 161.675 -127.325 162.005 -126.995 ;
        RECT 161.675 -128.685 162.005 -128.355 ;
        RECT 161.675 -130.045 162.005 -129.715 ;
        RECT 161.675 -131.405 162.005 -131.075 ;
        RECT 161.675 -132.765 162.005 -132.435 ;
        RECT 161.675 -134.125 162.005 -133.795 ;
        RECT 161.675 -135.485 162.005 -135.155 ;
        RECT 161.675 -136.845 162.005 -136.515 ;
        RECT 161.675 -138.205 162.005 -137.875 ;
        RECT 161.675 -139.565 162.005 -139.235 ;
        RECT 161.675 -140.925 162.005 -140.595 ;
        RECT 161.675 -142.285 162.005 -141.955 ;
        RECT 161.675 -143.645 162.005 -143.315 ;
        RECT 161.675 -145.005 162.005 -144.675 ;
        RECT 161.675 -146.365 162.005 -146.035 ;
        RECT 161.675 -147.725 162.005 -147.395 ;
        RECT 161.675 -149.085 162.005 -148.755 ;
        RECT 161.675 -150.445 162.005 -150.115 ;
        RECT 161.675 -151.805 162.005 -151.475 ;
        RECT 161.675 -153.165 162.005 -152.835 ;
        RECT 161.675 -154.525 162.005 -154.195 ;
        RECT 161.675 -155.885 162.005 -155.555 ;
        RECT 161.675 -157.245 162.005 -156.915 ;
        RECT 161.675 -158.605 162.005 -158.275 ;
        RECT 161.675 -159.965 162.005 -159.635 ;
        RECT 161.675 -161.325 162.005 -160.995 ;
        RECT 161.675 -162.685 162.005 -162.355 ;
        RECT 161.675 -164.045 162.005 -163.715 ;
        RECT 161.675 -165.405 162.005 -165.075 ;
        RECT 161.675 -166.765 162.005 -166.435 ;
        RECT 161.675 -168.125 162.005 -167.795 ;
        RECT 161.675 -169.485 162.005 -169.155 ;
        RECT 161.675 -170.845 162.005 -170.515 ;
        RECT 161.675 -172.205 162.005 -171.875 ;
        RECT 161.675 -173.565 162.005 -173.235 ;
        RECT 161.675 -174.925 162.005 -174.595 ;
        RECT 161.675 -176.285 162.005 -175.955 ;
        RECT 161.675 -177.645 162.005 -177.315 ;
        RECT 161.675 -179.005 162.005 -178.675 ;
        RECT 161.675 -180.365 162.005 -180.035 ;
        RECT 161.675 -181.725 162.005 -181.395 ;
        RECT 161.675 -183.085 162.005 -182.755 ;
        RECT 161.675 -184.445 162.005 -184.115 ;
        RECT 161.675 -185.805 162.005 -185.475 ;
        RECT 161.675 -187.165 162.005 -186.835 ;
        RECT 161.675 -188.525 162.005 -188.195 ;
        RECT 161.675 -189.885 162.005 -189.555 ;
        RECT 161.675 -191.245 162.005 -190.915 ;
        RECT 161.675 -192.605 162.005 -192.275 ;
        RECT 161.675 -193.965 162.005 -193.635 ;
        RECT 161.675 -195.325 162.005 -194.995 ;
        RECT 161.675 -196.685 162.005 -196.355 ;
        RECT 161.675 -198.045 162.005 -197.715 ;
        RECT 161.675 -199.405 162.005 -199.075 ;
        RECT 161.675 -200.765 162.005 -200.435 ;
        RECT 161.675 -202.125 162.005 -201.795 ;
        RECT 161.675 -203.485 162.005 -203.155 ;
        RECT 161.675 -204.845 162.005 -204.515 ;
        RECT 161.675 -206.205 162.005 -205.875 ;
        RECT 161.675 -207.565 162.005 -207.235 ;
        RECT 161.675 -208.925 162.005 -208.595 ;
        RECT 161.675 -210.285 162.005 -209.955 ;
        RECT 161.675 -211.645 162.005 -211.315 ;
        RECT 161.675 -213.005 162.005 -212.675 ;
        RECT 161.675 -214.365 162.005 -214.035 ;
        RECT 161.675 -215.725 162.005 -215.395 ;
        RECT 161.675 -217.085 162.005 -216.755 ;
        RECT 161.675 -218.445 162.005 -218.115 ;
        RECT 161.675 -224.09 162.005 -222.96 ;
        RECT 161.68 -224.205 162 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.035 132.52 163.365 133.65 ;
        RECT 163.035 128.355 163.365 128.685 ;
        RECT 163.035 126.995 163.365 127.325 ;
        RECT 163.035 125.635 163.365 125.965 ;
        RECT 163.035 124.275 163.365 124.605 ;
        RECT 163.04 123.6 163.36 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.035 -0.845 163.365 -0.515 ;
        RECT 163.035 -2.205 163.365 -1.875 ;
        RECT 163.035 -3.565 163.365 -3.235 ;
        RECT 163.04 -3.565 163.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.395 132.52 164.725 133.65 ;
        RECT 164.395 128.355 164.725 128.685 ;
        RECT 164.395 126.995 164.725 127.325 ;
        RECT 164.395 125.635 164.725 125.965 ;
        RECT 164.395 124.275 164.725 124.605 ;
        RECT 164.4 123.6 164.72 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.395 -0.845 164.725 -0.515 ;
        RECT 164.395 -2.205 164.725 -1.875 ;
        RECT 164.395 -3.565 164.725 -3.235 ;
        RECT 164.4 -3.565 164.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.755 132.52 166.085 133.65 ;
        RECT 165.755 128.355 166.085 128.685 ;
        RECT 165.755 126.995 166.085 127.325 ;
        RECT 165.755 125.635 166.085 125.965 ;
        RECT 165.755 124.275 166.085 124.605 ;
        RECT 165.76 123.6 166.08 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.755 -0.845 166.085 -0.515 ;
        RECT 165.755 -2.205 166.085 -1.875 ;
        RECT 165.755 -3.565 166.085 -3.235 ;
        RECT 165.76 -3.565 166.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.755 -224.09 166.085 -222.96 ;
        RECT 165.76 -224.205 166.08 -118.16 ;
        RECT 165.755 -119.165 166.085 -118.835 ;
        RECT 165.755 -120.525 166.085 -120.195 ;
        RECT 165.755 -121.885 166.085 -121.555 ;
        RECT 165.755 -123.245 166.085 -122.915 ;
        RECT 165.755 -124.605 166.085 -124.275 ;
        RECT 165.755 -125.965 166.085 -125.635 ;
        RECT 165.755 -127.325 166.085 -126.995 ;
        RECT 165.755 -128.685 166.085 -128.355 ;
        RECT 165.755 -130.045 166.085 -129.715 ;
        RECT 165.755 -131.405 166.085 -131.075 ;
        RECT 165.755 -132.765 166.085 -132.435 ;
        RECT 165.755 -134.125 166.085 -133.795 ;
        RECT 165.755 -135.485 166.085 -135.155 ;
        RECT 165.755 -136.845 166.085 -136.515 ;
        RECT 165.755 -138.205 166.085 -137.875 ;
        RECT 165.755 -139.565 166.085 -139.235 ;
        RECT 165.755 -140.925 166.085 -140.595 ;
        RECT 165.755 -142.285 166.085 -141.955 ;
        RECT 165.755 -143.645 166.085 -143.315 ;
        RECT 165.755 -145.005 166.085 -144.675 ;
        RECT 165.755 -146.365 166.085 -146.035 ;
        RECT 165.755 -147.725 166.085 -147.395 ;
        RECT 165.755 -149.085 166.085 -148.755 ;
        RECT 165.755 -150.445 166.085 -150.115 ;
        RECT 165.755 -151.805 166.085 -151.475 ;
        RECT 165.755 -153.165 166.085 -152.835 ;
        RECT 165.755 -154.525 166.085 -154.195 ;
        RECT 165.755 -155.885 166.085 -155.555 ;
        RECT 165.755 -157.245 166.085 -156.915 ;
        RECT 165.755 -158.605 166.085 -158.275 ;
        RECT 165.755 -159.965 166.085 -159.635 ;
        RECT 165.755 -161.325 166.085 -160.995 ;
        RECT 165.755 -162.685 166.085 -162.355 ;
        RECT 165.755 -164.045 166.085 -163.715 ;
        RECT 165.755 -165.405 166.085 -165.075 ;
        RECT 165.755 -166.765 166.085 -166.435 ;
        RECT 165.755 -168.125 166.085 -167.795 ;
        RECT 165.755 -169.485 166.085 -169.155 ;
        RECT 165.755 -170.845 166.085 -170.515 ;
        RECT 165.755 -172.205 166.085 -171.875 ;
        RECT 165.755 -173.565 166.085 -173.235 ;
        RECT 165.755 -174.925 166.085 -174.595 ;
        RECT 165.755 -176.285 166.085 -175.955 ;
        RECT 165.755 -177.645 166.085 -177.315 ;
        RECT 165.755 -179.005 166.085 -178.675 ;
        RECT 165.755 -180.365 166.085 -180.035 ;
        RECT 165.755 -181.725 166.085 -181.395 ;
        RECT 165.755 -183.085 166.085 -182.755 ;
        RECT 165.755 -184.445 166.085 -184.115 ;
        RECT 165.755 -185.805 166.085 -185.475 ;
        RECT 165.755 -187.165 166.085 -186.835 ;
        RECT 165.755 -188.525 166.085 -188.195 ;
        RECT 165.755 -189.885 166.085 -189.555 ;
        RECT 165.755 -191.245 166.085 -190.915 ;
        RECT 165.755 -192.605 166.085 -192.275 ;
        RECT 165.755 -193.965 166.085 -193.635 ;
        RECT 165.755 -195.325 166.085 -194.995 ;
        RECT 165.755 -196.685 166.085 -196.355 ;
        RECT 165.755 -198.045 166.085 -197.715 ;
        RECT 165.755 -199.405 166.085 -199.075 ;
        RECT 165.755 -200.765 166.085 -200.435 ;
        RECT 165.755 -202.125 166.085 -201.795 ;
        RECT 165.755 -203.485 166.085 -203.155 ;
        RECT 165.755 -204.845 166.085 -204.515 ;
        RECT 165.755 -206.205 166.085 -205.875 ;
        RECT 165.755 -207.565 166.085 -207.235 ;
        RECT 165.755 -208.925 166.085 -208.595 ;
        RECT 165.755 -210.285 166.085 -209.955 ;
        RECT 165.755 -211.645 166.085 -211.315 ;
        RECT 165.755 -213.005 166.085 -212.675 ;
        RECT 165.755 -214.365 166.085 -214.035 ;
        RECT 165.755 -215.725 166.085 -215.395 ;
        RECT 165.755 -217.085 166.085 -216.755 ;
        RECT 165.755 -218.445 166.085 -218.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.835 132.52 102.165 133.65 ;
        RECT 101.835 128.355 102.165 128.685 ;
        RECT 101.835 126.995 102.165 127.325 ;
        RECT 101.835 125.635 102.165 125.965 ;
        RECT 101.835 124.275 102.165 124.605 ;
        RECT 101.84 123.6 102.16 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.835 -0.845 102.165 -0.515 ;
        RECT 101.835 -2.205 102.165 -1.875 ;
        RECT 101.835 -3.565 102.165 -3.235 ;
        RECT 101.84 -3.565 102.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.195 132.52 103.525 133.65 ;
        RECT 103.195 128.355 103.525 128.685 ;
        RECT 103.195 126.995 103.525 127.325 ;
        RECT 103.195 125.635 103.525 125.965 ;
        RECT 103.195 124.275 103.525 124.605 ;
        RECT 103.2 123.6 103.52 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.195 -0.845 103.525 -0.515 ;
        RECT 103.195 -2.205 103.525 -1.875 ;
        RECT 103.195 -3.565 103.525 -3.235 ;
        RECT 103.2 -3.565 103.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.555 132.52 104.885 133.65 ;
        RECT 104.555 128.355 104.885 128.685 ;
        RECT 104.555 126.995 104.885 127.325 ;
        RECT 104.555 125.635 104.885 125.965 ;
        RECT 104.555 124.275 104.885 124.605 ;
        RECT 104.56 123.6 104.88 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.555 -0.845 104.885 -0.515 ;
        RECT 104.555 -2.205 104.885 -1.875 ;
        RECT 104.555 -3.565 104.885 -3.235 ;
        RECT 104.56 -3.565 104.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.915 132.52 106.245 133.65 ;
        RECT 105.915 128.355 106.245 128.685 ;
        RECT 105.915 126.995 106.245 127.325 ;
        RECT 105.915 125.635 106.245 125.965 ;
        RECT 105.915 124.275 106.245 124.605 ;
        RECT 105.92 123.6 106.24 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.915 -123.245 106.245 -122.915 ;
        RECT 105.915 -124.605 106.245 -124.275 ;
        RECT 105.915 -125.965 106.245 -125.635 ;
        RECT 105.915 -127.325 106.245 -126.995 ;
        RECT 105.915 -128.685 106.245 -128.355 ;
        RECT 105.915 -130.045 106.245 -129.715 ;
        RECT 105.915 -131.405 106.245 -131.075 ;
        RECT 105.915 -132.765 106.245 -132.435 ;
        RECT 105.915 -134.125 106.245 -133.795 ;
        RECT 105.915 -135.485 106.245 -135.155 ;
        RECT 105.915 -136.845 106.245 -136.515 ;
        RECT 105.915 -138.205 106.245 -137.875 ;
        RECT 105.915 -139.565 106.245 -139.235 ;
        RECT 105.915 -140.925 106.245 -140.595 ;
        RECT 105.915 -142.285 106.245 -141.955 ;
        RECT 105.915 -143.645 106.245 -143.315 ;
        RECT 105.915 -145.005 106.245 -144.675 ;
        RECT 105.915 -146.365 106.245 -146.035 ;
        RECT 105.915 -147.725 106.245 -147.395 ;
        RECT 105.915 -149.085 106.245 -148.755 ;
        RECT 105.915 -150.445 106.245 -150.115 ;
        RECT 105.915 -151.805 106.245 -151.475 ;
        RECT 105.915 -153.165 106.245 -152.835 ;
        RECT 105.915 -154.525 106.245 -154.195 ;
        RECT 105.915 -155.885 106.245 -155.555 ;
        RECT 105.915 -157.245 106.245 -156.915 ;
        RECT 105.915 -158.605 106.245 -158.275 ;
        RECT 105.915 -159.965 106.245 -159.635 ;
        RECT 105.915 -161.325 106.245 -160.995 ;
        RECT 105.915 -162.685 106.245 -162.355 ;
        RECT 105.915 -164.045 106.245 -163.715 ;
        RECT 105.915 -165.405 106.245 -165.075 ;
        RECT 105.915 -166.765 106.245 -166.435 ;
        RECT 105.915 -168.125 106.245 -167.795 ;
        RECT 105.915 -169.485 106.245 -169.155 ;
        RECT 105.915 -170.845 106.245 -170.515 ;
        RECT 105.915 -172.205 106.245 -171.875 ;
        RECT 105.915 -173.565 106.245 -173.235 ;
        RECT 105.915 -174.925 106.245 -174.595 ;
        RECT 105.915 -176.285 106.245 -175.955 ;
        RECT 105.915 -177.645 106.245 -177.315 ;
        RECT 105.915 -179.005 106.245 -178.675 ;
        RECT 105.915 -180.365 106.245 -180.035 ;
        RECT 105.915 -181.725 106.245 -181.395 ;
        RECT 105.915 -183.085 106.245 -182.755 ;
        RECT 105.915 -184.445 106.245 -184.115 ;
        RECT 105.915 -185.805 106.245 -185.475 ;
        RECT 105.915 -187.165 106.245 -186.835 ;
        RECT 105.915 -188.525 106.245 -188.195 ;
        RECT 105.915 -189.885 106.245 -189.555 ;
        RECT 105.915 -191.245 106.245 -190.915 ;
        RECT 105.915 -192.605 106.245 -192.275 ;
        RECT 105.915 -193.965 106.245 -193.635 ;
        RECT 105.915 -195.325 106.245 -194.995 ;
        RECT 105.915 -196.685 106.245 -196.355 ;
        RECT 105.915 -198.045 106.245 -197.715 ;
        RECT 105.915 -199.405 106.245 -199.075 ;
        RECT 105.915 -200.765 106.245 -200.435 ;
        RECT 105.915 -202.125 106.245 -201.795 ;
        RECT 105.915 -203.485 106.245 -203.155 ;
        RECT 105.915 -204.845 106.245 -204.515 ;
        RECT 105.915 -206.205 106.245 -205.875 ;
        RECT 105.915 -207.565 106.245 -207.235 ;
        RECT 105.915 -208.925 106.245 -208.595 ;
        RECT 105.915 -210.285 106.245 -209.955 ;
        RECT 105.915 -211.645 106.245 -211.315 ;
        RECT 105.915 -213.005 106.245 -212.675 ;
        RECT 105.915 -214.365 106.245 -214.035 ;
        RECT 105.915 -215.725 106.245 -215.395 ;
        RECT 105.915 -217.085 106.245 -216.755 ;
        RECT 105.915 -218.445 106.245 -218.115 ;
        RECT 105.915 -224.09 106.245 -222.96 ;
        RECT 105.92 -224.205 106.24 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.36 -121.535 106.69 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.275 132.52 107.605 133.65 ;
        RECT 107.275 128.355 107.605 128.685 ;
        RECT 107.275 126.995 107.605 127.325 ;
        RECT 107.275 125.635 107.605 125.965 ;
        RECT 107.275 124.275 107.605 124.605 ;
        RECT 107.28 123.6 107.6 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.635 132.52 108.965 133.65 ;
        RECT 108.635 128.355 108.965 128.685 ;
        RECT 108.635 126.995 108.965 127.325 ;
        RECT 108.635 125.635 108.965 125.965 ;
        RECT 108.635 124.275 108.965 124.605 ;
        RECT 108.64 123.6 108.96 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.635 -0.845 108.965 -0.515 ;
        RECT 108.635 -2.205 108.965 -1.875 ;
        RECT 108.635 -3.565 108.965 -3.235 ;
        RECT 108.64 -3.565 108.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.995 132.52 110.325 133.65 ;
        RECT 109.995 128.355 110.325 128.685 ;
        RECT 109.995 126.995 110.325 127.325 ;
        RECT 109.995 125.635 110.325 125.965 ;
        RECT 109.995 124.275 110.325 124.605 ;
        RECT 110 123.6 110.32 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.995 -0.845 110.325 -0.515 ;
        RECT 109.995 -2.205 110.325 -1.875 ;
        RECT 109.995 -3.565 110.325 -3.235 ;
        RECT 110 -3.565 110.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.355 132.52 111.685 133.65 ;
        RECT 111.355 128.355 111.685 128.685 ;
        RECT 111.355 126.995 111.685 127.325 ;
        RECT 111.355 125.635 111.685 125.965 ;
        RECT 111.355 124.275 111.685 124.605 ;
        RECT 111.36 123.6 111.68 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.355 -0.845 111.685 -0.515 ;
        RECT 111.355 -2.205 111.685 -1.875 ;
        RECT 111.355 -3.565 111.685 -3.235 ;
        RECT 111.36 -3.565 111.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.355 -119.165 111.685 -118.835 ;
        RECT 111.355 -120.525 111.685 -120.195 ;
        RECT 111.355 -121.885 111.685 -121.555 ;
        RECT 111.355 -123.245 111.685 -122.915 ;
        RECT 111.355 -124.605 111.685 -124.275 ;
        RECT 111.355 -125.965 111.685 -125.635 ;
        RECT 111.355 -127.325 111.685 -126.995 ;
        RECT 111.355 -128.685 111.685 -128.355 ;
        RECT 111.355 -130.045 111.685 -129.715 ;
        RECT 111.355 -131.405 111.685 -131.075 ;
        RECT 111.355 -132.765 111.685 -132.435 ;
        RECT 111.355 -134.125 111.685 -133.795 ;
        RECT 111.355 -135.485 111.685 -135.155 ;
        RECT 111.355 -136.845 111.685 -136.515 ;
        RECT 111.355 -138.205 111.685 -137.875 ;
        RECT 111.355 -139.565 111.685 -139.235 ;
        RECT 111.355 -140.925 111.685 -140.595 ;
        RECT 111.355 -142.285 111.685 -141.955 ;
        RECT 111.355 -143.645 111.685 -143.315 ;
        RECT 111.355 -145.005 111.685 -144.675 ;
        RECT 111.355 -146.365 111.685 -146.035 ;
        RECT 111.355 -147.725 111.685 -147.395 ;
        RECT 111.355 -149.085 111.685 -148.755 ;
        RECT 111.355 -150.445 111.685 -150.115 ;
        RECT 111.355 -151.805 111.685 -151.475 ;
        RECT 111.355 -153.165 111.685 -152.835 ;
        RECT 111.355 -154.525 111.685 -154.195 ;
        RECT 111.355 -155.885 111.685 -155.555 ;
        RECT 111.355 -157.245 111.685 -156.915 ;
        RECT 111.355 -158.605 111.685 -158.275 ;
        RECT 111.355 -159.965 111.685 -159.635 ;
        RECT 111.355 -161.325 111.685 -160.995 ;
        RECT 111.355 -162.685 111.685 -162.355 ;
        RECT 111.355 -164.045 111.685 -163.715 ;
        RECT 111.355 -165.405 111.685 -165.075 ;
        RECT 111.355 -166.765 111.685 -166.435 ;
        RECT 111.355 -168.125 111.685 -167.795 ;
        RECT 111.355 -169.485 111.685 -169.155 ;
        RECT 111.355 -170.845 111.685 -170.515 ;
        RECT 111.355 -172.205 111.685 -171.875 ;
        RECT 111.355 -173.565 111.685 -173.235 ;
        RECT 111.355 -174.925 111.685 -174.595 ;
        RECT 111.355 -176.285 111.685 -175.955 ;
        RECT 111.355 -177.645 111.685 -177.315 ;
        RECT 111.355 -179.005 111.685 -178.675 ;
        RECT 111.355 -180.365 111.685 -180.035 ;
        RECT 111.355 -181.725 111.685 -181.395 ;
        RECT 111.355 -183.085 111.685 -182.755 ;
        RECT 111.355 -184.445 111.685 -184.115 ;
        RECT 111.355 -185.805 111.685 -185.475 ;
        RECT 111.355 -187.165 111.685 -186.835 ;
        RECT 111.355 -188.525 111.685 -188.195 ;
        RECT 111.355 -189.885 111.685 -189.555 ;
        RECT 111.355 -191.245 111.685 -190.915 ;
        RECT 111.355 -192.605 111.685 -192.275 ;
        RECT 111.355 -193.965 111.685 -193.635 ;
        RECT 111.355 -195.325 111.685 -194.995 ;
        RECT 111.355 -196.685 111.685 -196.355 ;
        RECT 111.355 -198.045 111.685 -197.715 ;
        RECT 111.355 -199.405 111.685 -199.075 ;
        RECT 111.355 -200.765 111.685 -200.435 ;
        RECT 111.355 -202.125 111.685 -201.795 ;
        RECT 111.355 -203.485 111.685 -203.155 ;
        RECT 111.355 -204.845 111.685 -204.515 ;
        RECT 111.355 -206.205 111.685 -205.875 ;
        RECT 111.355 -207.565 111.685 -207.235 ;
        RECT 111.355 -208.925 111.685 -208.595 ;
        RECT 111.355 -210.285 111.685 -209.955 ;
        RECT 111.355 -211.645 111.685 -211.315 ;
        RECT 111.355 -213.005 111.685 -212.675 ;
        RECT 111.355 -214.365 111.685 -214.035 ;
        RECT 111.355 -215.725 111.685 -215.395 ;
        RECT 111.355 -217.085 111.685 -216.755 ;
        RECT 111.355 -218.445 111.685 -218.115 ;
        RECT 111.355 -224.09 111.685 -222.96 ;
        RECT 111.36 -224.205 111.68 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.46 -121.535 112.79 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.715 132.52 113.045 133.65 ;
        RECT 112.715 128.355 113.045 128.685 ;
        RECT 112.715 126.995 113.045 127.325 ;
        RECT 112.715 125.635 113.045 125.965 ;
        RECT 112.715 124.275 113.045 124.605 ;
        RECT 112.72 123.6 113.04 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.715 -123.245 113.045 -122.915 ;
        RECT 112.715 -124.605 113.045 -124.275 ;
        RECT 112.715 -125.965 113.045 -125.635 ;
        RECT 112.715 -127.325 113.045 -126.995 ;
        RECT 112.715 -128.685 113.045 -128.355 ;
        RECT 112.715 -130.045 113.045 -129.715 ;
        RECT 112.715 -131.405 113.045 -131.075 ;
        RECT 112.715 -132.765 113.045 -132.435 ;
        RECT 112.715 -134.125 113.045 -133.795 ;
        RECT 112.715 -135.485 113.045 -135.155 ;
        RECT 112.715 -136.845 113.045 -136.515 ;
        RECT 112.715 -138.205 113.045 -137.875 ;
        RECT 112.715 -139.565 113.045 -139.235 ;
        RECT 112.715 -140.925 113.045 -140.595 ;
        RECT 112.715 -142.285 113.045 -141.955 ;
        RECT 112.715 -143.645 113.045 -143.315 ;
        RECT 112.715 -145.005 113.045 -144.675 ;
        RECT 112.715 -146.365 113.045 -146.035 ;
        RECT 112.715 -147.725 113.045 -147.395 ;
        RECT 112.715 -149.085 113.045 -148.755 ;
        RECT 112.715 -150.445 113.045 -150.115 ;
        RECT 112.715 -151.805 113.045 -151.475 ;
        RECT 112.715 -153.165 113.045 -152.835 ;
        RECT 112.715 -154.525 113.045 -154.195 ;
        RECT 112.715 -155.885 113.045 -155.555 ;
        RECT 112.715 -157.245 113.045 -156.915 ;
        RECT 112.715 -158.605 113.045 -158.275 ;
        RECT 112.715 -159.965 113.045 -159.635 ;
        RECT 112.715 -161.325 113.045 -160.995 ;
        RECT 112.715 -162.685 113.045 -162.355 ;
        RECT 112.715 -164.045 113.045 -163.715 ;
        RECT 112.715 -165.405 113.045 -165.075 ;
        RECT 112.715 -166.765 113.045 -166.435 ;
        RECT 112.715 -168.125 113.045 -167.795 ;
        RECT 112.715 -169.485 113.045 -169.155 ;
        RECT 112.715 -170.845 113.045 -170.515 ;
        RECT 112.715 -172.205 113.045 -171.875 ;
        RECT 112.715 -173.565 113.045 -173.235 ;
        RECT 112.715 -174.925 113.045 -174.595 ;
        RECT 112.715 -176.285 113.045 -175.955 ;
        RECT 112.715 -177.645 113.045 -177.315 ;
        RECT 112.715 -179.005 113.045 -178.675 ;
        RECT 112.715 -180.365 113.045 -180.035 ;
        RECT 112.715 -181.725 113.045 -181.395 ;
        RECT 112.715 -183.085 113.045 -182.755 ;
        RECT 112.715 -184.445 113.045 -184.115 ;
        RECT 112.715 -185.805 113.045 -185.475 ;
        RECT 112.715 -187.165 113.045 -186.835 ;
        RECT 112.715 -188.525 113.045 -188.195 ;
        RECT 112.715 -189.885 113.045 -189.555 ;
        RECT 112.715 -191.245 113.045 -190.915 ;
        RECT 112.715 -192.605 113.045 -192.275 ;
        RECT 112.715 -193.965 113.045 -193.635 ;
        RECT 112.715 -195.325 113.045 -194.995 ;
        RECT 112.715 -196.685 113.045 -196.355 ;
        RECT 112.715 -198.045 113.045 -197.715 ;
        RECT 112.715 -199.405 113.045 -199.075 ;
        RECT 112.715 -200.765 113.045 -200.435 ;
        RECT 112.715 -202.125 113.045 -201.795 ;
        RECT 112.715 -203.485 113.045 -203.155 ;
        RECT 112.715 -204.845 113.045 -204.515 ;
        RECT 112.715 -206.205 113.045 -205.875 ;
        RECT 112.715 -207.565 113.045 -207.235 ;
        RECT 112.715 -208.925 113.045 -208.595 ;
        RECT 112.715 -210.285 113.045 -209.955 ;
        RECT 112.715 -211.645 113.045 -211.315 ;
        RECT 112.715 -213.005 113.045 -212.675 ;
        RECT 112.715 -214.365 113.045 -214.035 ;
        RECT 112.715 -215.725 113.045 -215.395 ;
        RECT 112.715 -217.085 113.045 -216.755 ;
        RECT 112.715 -218.445 113.045 -218.115 ;
        RECT 112.715 -224.09 113.045 -222.96 ;
        RECT 112.72 -224.205 113.04 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.075 132.52 114.405 133.65 ;
        RECT 114.075 128.355 114.405 128.685 ;
        RECT 114.075 126.995 114.405 127.325 ;
        RECT 114.075 125.635 114.405 125.965 ;
        RECT 114.075 124.275 114.405 124.605 ;
        RECT 114.08 123.6 114.4 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.075 -0.845 114.405 -0.515 ;
        RECT 114.075 -2.205 114.405 -1.875 ;
        RECT 114.075 -3.565 114.405 -3.235 ;
        RECT 114.08 -3.565 114.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.435 132.52 115.765 133.65 ;
        RECT 115.435 128.355 115.765 128.685 ;
        RECT 115.435 126.995 115.765 127.325 ;
        RECT 115.435 125.635 115.765 125.965 ;
        RECT 115.435 124.275 115.765 124.605 ;
        RECT 115.44 123.6 115.76 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.435 -0.845 115.765 -0.515 ;
        RECT 115.435 -2.205 115.765 -1.875 ;
        RECT 115.435 -3.565 115.765 -3.235 ;
        RECT 115.44 -3.565 115.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.795 132.52 117.125 133.65 ;
        RECT 116.795 128.355 117.125 128.685 ;
        RECT 116.795 126.995 117.125 127.325 ;
        RECT 116.795 125.635 117.125 125.965 ;
        RECT 116.795 124.275 117.125 124.605 ;
        RECT 116.8 123.6 117.12 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.795 -0.845 117.125 -0.515 ;
        RECT 116.795 -2.205 117.125 -1.875 ;
        RECT 116.795 -3.565 117.125 -3.235 ;
        RECT 116.8 -3.565 117.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.795 -119.165 117.125 -118.835 ;
        RECT 116.795 -120.525 117.125 -120.195 ;
        RECT 116.795 -121.885 117.125 -121.555 ;
        RECT 116.795 -123.245 117.125 -122.915 ;
        RECT 116.795 -124.605 117.125 -124.275 ;
        RECT 116.795 -125.965 117.125 -125.635 ;
        RECT 116.795 -127.325 117.125 -126.995 ;
        RECT 116.795 -128.685 117.125 -128.355 ;
        RECT 116.795 -130.045 117.125 -129.715 ;
        RECT 116.795 -131.405 117.125 -131.075 ;
        RECT 116.795 -132.765 117.125 -132.435 ;
        RECT 116.795 -134.125 117.125 -133.795 ;
        RECT 116.795 -135.485 117.125 -135.155 ;
        RECT 116.795 -136.845 117.125 -136.515 ;
        RECT 116.795 -138.205 117.125 -137.875 ;
        RECT 116.795 -139.565 117.125 -139.235 ;
        RECT 116.795 -140.925 117.125 -140.595 ;
        RECT 116.795 -142.285 117.125 -141.955 ;
        RECT 116.795 -143.645 117.125 -143.315 ;
        RECT 116.795 -145.005 117.125 -144.675 ;
        RECT 116.795 -146.365 117.125 -146.035 ;
        RECT 116.795 -147.725 117.125 -147.395 ;
        RECT 116.795 -149.085 117.125 -148.755 ;
        RECT 116.795 -150.445 117.125 -150.115 ;
        RECT 116.795 -151.805 117.125 -151.475 ;
        RECT 116.795 -153.165 117.125 -152.835 ;
        RECT 116.795 -154.525 117.125 -154.195 ;
        RECT 116.795 -155.885 117.125 -155.555 ;
        RECT 116.795 -157.245 117.125 -156.915 ;
        RECT 116.795 -158.605 117.125 -158.275 ;
        RECT 116.795 -159.965 117.125 -159.635 ;
        RECT 116.795 -161.325 117.125 -160.995 ;
        RECT 116.795 -162.685 117.125 -162.355 ;
        RECT 116.795 -164.045 117.125 -163.715 ;
        RECT 116.795 -165.405 117.125 -165.075 ;
        RECT 116.795 -166.765 117.125 -166.435 ;
        RECT 116.795 -168.125 117.125 -167.795 ;
        RECT 116.795 -169.485 117.125 -169.155 ;
        RECT 116.795 -170.845 117.125 -170.515 ;
        RECT 116.795 -172.205 117.125 -171.875 ;
        RECT 116.795 -173.565 117.125 -173.235 ;
        RECT 116.795 -174.925 117.125 -174.595 ;
        RECT 116.795 -176.285 117.125 -175.955 ;
        RECT 116.795 -177.645 117.125 -177.315 ;
        RECT 116.795 -179.005 117.125 -178.675 ;
        RECT 116.795 -180.365 117.125 -180.035 ;
        RECT 116.795 -181.725 117.125 -181.395 ;
        RECT 116.795 -183.085 117.125 -182.755 ;
        RECT 116.795 -184.445 117.125 -184.115 ;
        RECT 116.795 -185.805 117.125 -185.475 ;
        RECT 116.795 -187.165 117.125 -186.835 ;
        RECT 116.795 -188.525 117.125 -188.195 ;
        RECT 116.795 -189.885 117.125 -189.555 ;
        RECT 116.795 -191.245 117.125 -190.915 ;
        RECT 116.795 -192.605 117.125 -192.275 ;
        RECT 116.795 -193.965 117.125 -193.635 ;
        RECT 116.795 -195.325 117.125 -194.995 ;
        RECT 116.795 -196.685 117.125 -196.355 ;
        RECT 116.795 -198.045 117.125 -197.715 ;
        RECT 116.795 -199.405 117.125 -199.075 ;
        RECT 116.795 -200.765 117.125 -200.435 ;
        RECT 116.795 -202.125 117.125 -201.795 ;
        RECT 116.795 -203.485 117.125 -203.155 ;
        RECT 116.795 -204.845 117.125 -204.515 ;
        RECT 116.795 -206.205 117.125 -205.875 ;
        RECT 116.795 -207.565 117.125 -207.235 ;
        RECT 116.795 -208.925 117.125 -208.595 ;
        RECT 116.795 -210.285 117.125 -209.955 ;
        RECT 116.795 -211.645 117.125 -211.315 ;
        RECT 116.795 -213.005 117.125 -212.675 ;
        RECT 116.795 -214.365 117.125 -214.035 ;
        RECT 116.795 -215.725 117.125 -215.395 ;
        RECT 116.795 -217.085 117.125 -216.755 ;
        RECT 116.795 -218.445 117.125 -218.115 ;
        RECT 116.795 -224.09 117.125 -222.96 ;
        RECT 116.8 -224.205 117.12 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.155 132.52 118.485 133.65 ;
        RECT 118.155 128.355 118.485 128.685 ;
        RECT 118.155 126.995 118.485 127.325 ;
        RECT 118.155 125.635 118.485 125.965 ;
        RECT 118.155 124.275 118.485 124.605 ;
        RECT 118.16 123.6 118.48 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.155 -123.245 118.485 -122.915 ;
        RECT 118.155 -124.605 118.485 -124.275 ;
        RECT 118.155 -125.965 118.485 -125.635 ;
        RECT 118.155 -127.325 118.485 -126.995 ;
        RECT 118.155 -128.685 118.485 -128.355 ;
        RECT 118.155 -130.045 118.485 -129.715 ;
        RECT 118.155 -131.405 118.485 -131.075 ;
        RECT 118.155 -132.765 118.485 -132.435 ;
        RECT 118.155 -134.125 118.485 -133.795 ;
        RECT 118.155 -135.485 118.485 -135.155 ;
        RECT 118.155 -136.845 118.485 -136.515 ;
        RECT 118.155 -138.205 118.485 -137.875 ;
        RECT 118.155 -139.565 118.485 -139.235 ;
        RECT 118.155 -140.925 118.485 -140.595 ;
        RECT 118.155 -142.285 118.485 -141.955 ;
        RECT 118.155 -143.645 118.485 -143.315 ;
        RECT 118.155 -145.005 118.485 -144.675 ;
        RECT 118.155 -146.365 118.485 -146.035 ;
        RECT 118.155 -147.725 118.485 -147.395 ;
        RECT 118.155 -149.085 118.485 -148.755 ;
        RECT 118.155 -150.445 118.485 -150.115 ;
        RECT 118.155 -151.805 118.485 -151.475 ;
        RECT 118.155 -153.165 118.485 -152.835 ;
        RECT 118.155 -154.525 118.485 -154.195 ;
        RECT 118.155 -155.885 118.485 -155.555 ;
        RECT 118.155 -157.245 118.485 -156.915 ;
        RECT 118.155 -158.605 118.485 -158.275 ;
        RECT 118.155 -159.965 118.485 -159.635 ;
        RECT 118.155 -161.325 118.485 -160.995 ;
        RECT 118.155 -162.685 118.485 -162.355 ;
        RECT 118.155 -164.045 118.485 -163.715 ;
        RECT 118.155 -165.405 118.485 -165.075 ;
        RECT 118.155 -166.765 118.485 -166.435 ;
        RECT 118.155 -168.125 118.485 -167.795 ;
        RECT 118.155 -169.485 118.485 -169.155 ;
        RECT 118.155 -170.845 118.485 -170.515 ;
        RECT 118.155 -172.205 118.485 -171.875 ;
        RECT 118.155 -173.565 118.485 -173.235 ;
        RECT 118.155 -174.925 118.485 -174.595 ;
        RECT 118.155 -176.285 118.485 -175.955 ;
        RECT 118.155 -177.645 118.485 -177.315 ;
        RECT 118.155 -179.005 118.485 -178.675 ;
        RECT 118.155 -180.365 118.485 -180.035 ;
        RECT 118.155 -181.725 118.485 -181.395 ;
        RECT 118.155 -183.085 118.485 -182.755 ;
        RECT 118.155 -184.445 118.485 -184.115 ;
        RECT 118.155 -185.805 118.485 -185.475 ;
        RECT 118.155 -187.165 118.485 -186.835 ;
        RECT 118.155 -188.525 118.485 -188.195 ;
        RECT 118.155 -189.885 118.485 -189.555 ;
        RECT 118.155 -191.245 118.485 -190.915 ;
        RECT 118.155 -192.605 118.485 -192.275 ;
        RECT 118.155 -193.965 118.485 -193.635 ;
        RECT 118.155 -195.325 118.485 -194.995 ;
        RECT 118.155 -196.685 118.485 -196.355 ;
        RECT 118.155 -198.045 118.485 -197.715 ;
        RECT 118.155 -199.405 118.485 -199.075 ;
        RECT 118.155 -200.765 118.485 -200.435 ;
        RECT 118.155 -202.125 118.485 -201.795 ;
        RECT 118.155 -203.485 118.485 -203.155 ;
        RECT 118.155 -204.845 118.485 -204.515 ;
        RECT 118.155 -206.205 118.485 -205.875 ;
        RECT 118.155 -207.565 118.485 -207.235 ;
        RECT 118.155 -208.925 118.485 -208.595 ;
        RECT 118.155 -210.285 118.485 -209.955 ;
        RECT 118.155 -211.645 118.485 -211.315 ;
        RECT 118.155 -213.005 118.485 -212.675 ;
        RECT 118.155 -214.365 118.485 -214.035 ;
        RECT 118.155 -215.725 118.485 -215.395 ;
        RECT 118.155 -217.085 118.485 -216.755 ;
        RECT 118.155 -218.445 118.485 -218.115 ;
        RECT 118.155 -224.09 118.485 -222.96 ;
        RECT 118.16 -224.205 118.48 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.56 -121.535 118.89 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.515 132.52 119.845 133.65 ;
        RECT 119.515 128.355 119.845 128.685 ;
        RECT 119.515 126.995 119.845 127.325 ;
        RECT 119.515 125.635 119.845 125.965 ;
        RECT 119.515 124.275 119.845 124.605 ;
        RECT 119.52 123.6 119.84 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.875 132.52 121.205 133.65 ;
        RECT 120.875 128.355 121.205 128.685 ;
        RECT 120.875 126.995 121.205 127.325 ;
        RECT 120.875 125.635 121.205 125.965 ;
        RECT 120.875 124.275 121.205 124.605 ;
        RECT 120.88 123.6 121.2 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.875 -0.845 121.205 -0.515 ;
        RECT 120.875 -2.205 121.205 -1.875 ;
        RECT 120.875 -3.565 121.205 -3.235 ;
        RECT 120.88 -3.565 121.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.235 132.52 122.565 133.65 ;
        RECT 122.235 128.355 122.565 128.685 ;
        RECT 122.235 126.995 122.565 127.325 ;
        RECT 122.235 125.635 122.565 125.965 ;
        RECT 122.235 124.275 122.565 124.605 ;
        RECT 122.24 123.6 122.56 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.235 -0.845 122.565 -0.515 ;
        RECT 122.235 -2.205 122.565 -1.875 ;
        RECT 122.235 -3.565 122.565 -3.235 ;
        RECT 122.24 -3.565 122.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.595 132.52 123.925 133.65 ;
        RECT 123.595 128.355 123.925 128.685 ;
        RECT 123.595 126.995 123.925 127.325 ;
        RECT 123.595 125.635 123.925 125.965 ;
        RECT 123.595 124.275 123.925 124.605 ;
        RECT 123.6 123.6 123.92 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.595 -0.845 123.925 -0.515 ;
        RECT 123.595 -2.205 123.925 -1.875 ;
        RECT 123.595 -3.565 123.925 -3.235 ;
        RECT 123.6 -3.565 123.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.595 -119.165 123.925 -118.835 ;
        RECT 123.595 -120.525 123.925 -120.195 ;
        RECT 123.595 -121.885 123.925 -121.555 ;
        RECT 123.595 -123.245 123.925 -122.915 ;
        RECT 123.595 -124.605 123.925 -124.275 ;
        RECT 123.595 -125.965 123.925 -125.635 ;
        RECT 123.595 -127.325 123.925 -126.995 ;
        RECT 123.595 -128.685 123.925 -128.355 ;
        RECT 123.595 -130.045 123.925 -129.715 ;
        RECT 123.595 -131.405 123.925 -131.075 ;
        RECT 123.595 -132.765 123.925 -132.435 ;
        RECT 123.595 -134.125 123.925 -133.795 ;
        RECT 123.595 -135.485 123.925 -135.155 ;
        RECT 123.595 -136.845 123.925 -136.515 ;
        RECT 123.595 -138.205 123.925 -137.875 ;
        RECT 123.595 -139.565 123.925 -139.235 ;
        RECT 123.595 -140.925 123.925 -140.595 ;
        RECT 123.595 -142.285 123.925 -141.955 ;
        RECT 123.595 -143.645 123.925 -143.315 ;
        RECT 123.595 -145.005 123.925 -144.675 ;
        RECT 123.595 -146.365 123.925 -146.035 ;
        RECT 123.595 -147.725 123.925 -147.395 ;
        RECT 123.595 -149.085 123.925 -148.755 ;
        RECT 123.595 -150.445 123.925 -150.115 ;
        RECT 123.595 -151.805 123.925 -151.475 ;
        RECT 123.595 -153.165 123.925 -152.835 ;
        RECT 123.595 -154.525 123.925 -154.195 ;
        RECT 123.595 -155.885 123.925 -155.555 ;
        RECT 123.595 -157.245 123.925 -156.915 ;
        RECT 123.595 -158.605 123.925 -158.275 ;
        RECT 123.595 -159.965 123.925 -159.635 ;
        RECT 123.595 -161.325 123.925 -160.995 ;
        RECT 123.595 -162.685 123.925 -162.355 ;
        RECT 123.595 -164.045 123.925 -163.715 ;
        RECT 123.595 -165.405 123.925 -165.075 ;
        RECT 123.595 -166.765 123.925 -166.435 ;
        RECT 123.595 -168.125 123.925 -167.795 ;
        RECT 123.595 -169.485 123.925 -169.155 ;
        RECT 123.595 -170.845 123.925 -170.515 ;
        RECT 123.595 -172.205 123.925 -171.875 ;
        RECT 123.595 -173.565 123.925 -173.235 ;
        RECT 123.595 -174.925 123.925 -174.595 ;
        RECT 123.595 -176.285 123.925 -175.955 ;
        RECT 123.595 -177.645 123.925 -177.315 ;
        RECT 123.595 -179.005 123.925 -178.675 ;
        RECT 123.595 -180.365 123.925 -180.035 ;
        RECT 123.595 -181.725 123.925 -181.395 ;
        RECT 123.595 -183.085 123.925 -182.755 ;
        RECT 123.595 -184.445 123.925 -184.115 ;
        RECT 123.595 -185.805 123.925 -185.475 ;
        RECT 123.595 -187.165 123.925 -186.835 ;
        RECT 123.595 -188.525 123.925 -188.195 ;
        RECT 123.595 -189.885 123.925 -189.555 ;
        RECT 123.595 -191.245 123.925 -190.915 ;
        RECT 123.595 -192.605 123.925 -192.275 ;
        RECT 123.595 -193.965 123.925 -193.635 ;
        RECT 123.595 -195.325 123.925 -194.995 ;
        RECT 123.595 -196.685 123.925 -196.355 ;
        RECT 123.595 -198.045 123.925 -197.715 ;
        RECT 123.595 -199.405 123.925 -199.075 ;
        RECT 123.595 -200.765 123.925 -200.435 ;
        RECT 123.595 -202.125 123.925 -201.795 ;
        RECT 123.595 -203.485 123.925 -203.155 ;
        RECT 123.595 -204.845 123.925 -204.515 ;
        RECT 123.595 -206.205 123.925 -205.875 ;
        RECT 123.595 -207.565 123.925 -207.235 ;
        RECT 123.595 -208.925 123.925 -208.595 ;
        RECT 123.595 -210.285 123.925 -209.955 ;
        RECT 123.595 -211.645 123.925 -211.315 ;
        RECT 123.595 -213.005 123.925 -212.675 ;
        RECT 123.595 -214.365 123.925 -214.035 ;
        RECT 123.595 -215.725 123.925 -215.395 ;
        RECT 123.595 -217.085 123.925 -216.755 ;
        RECT 123.595 -218.445 123.925 -218.115 ;
        RECT 123.595 -224.09 123.925 -222.96 ;
        RECT 123.6 -224.205 123.92 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.66 -121.535 124.99 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.955 132.52 125.285 133.65 ;
        RECT 124.955 128.355 125.285 128.685 ;
        RECT 124.955 126.995 125.285 127.325 ;
        RECT 124.955 125.635 125.285 125.965 ;
        RECT 124.955 124.275 125.285 124.605 ;
        RECT 124.96 123.6 125.28 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.955 -123.245 125.285 -122.915 ;
        RECT 124.955 -124.605 125.285 -124.275 ;
        RECT 124.955 -125.965 125.285 -125.635 ;
        RECT 124.955 -127.325 125.285 -126.995 ;
        RECT 124.955 -128.685 125.285 -128.355 ;
        RECT 124.955 -130.045 125.285 -129.715 ;
        RECT 124.955 -131.405 125.285 -131.075 ;
        RECT 124.955 -132.765 125.285 -132.435 ;
        RECT 124.955 -134.125 125.285 -133.795 ;
        RECT 124.955 -135.485 125.285 -135.155 ;
        RECT 124.955 -136.845 125.285 -136.515 ;
        RECT 124.955 -138.205 125.285 -137.875 ;
        RECT 124.955 -139.565 125.285 -139.235 ;
        RECT 124.955 -140.925 125.285 -140.595 ;
        RECT 124.955 -142.285 125.285 -141.955 ;
        RECT 124.955 -143.645 125.285 -143.315 ;
        RECT 124.955 -145.005 125.285 -144.675 ;
        RECT 124.955 -146.365 125.285 -146.035 ;
        RECT 124.955 -147.725 125.285 -147.395 ;
        RECT 124.955 -149.085 125.285 -148.755 ;
        RECT 124.955 -150.445 125.285 -150.115 ;
        RECT 124.955 -151.805 125.285 -151.475 ;
        RECT 124.955 -153.165 125.285 -152.835 ;
        RECT 124.955 -154.525 125.285 -154.195 ;
        RECT 124.955 -155.885 125.285 -155.555 ;
        RECT 124.955 -157.245 125.285 -156.915 ;
        RECT 124.955 -158.605 125.285 -158.275 ;
        RECT 124.955 -159.965 125.285 -159.635 ;
        RECT 124.955 -161.325 125.285 -160.995 ;
        RECT 124.955 -162.685 125.285 -162.355 ;
        RECT 124.955 -164.045 125.285 -163.715 ;
        RECT 124.955 -165.405 125.285 -165.075 ;
        RECT 124.955 -166.765 125.285 -166.435 ;
        RECT 124.955 -168.125 125.285 -167.795 ;
        RECT 124.955 -169.485 125.285 -169.155 ;
        RECT 124.955 -170.845 125.285 -170.515 ;
        RECT 124.955 -172.205 125.285 -171.875 ;
        RECT 124.955 -173.565 125.285 -173.235 ;
        RECT 124.955 -174.925 125.285 -174.595 ;
        RECT 124.955 -176.285 125.285 -175.955 ;
        RECT 124.955 -177.645 125.285 -177.315 ;
        RECT 124.955 -179.005 125.285 -178.675 ;
        RECT 124.955 -180.365 125.285 -180.035 ;
        RECT 124.955 -181.725 125.285 -181.395 ;
        RECT 124.955 -183.085 125.285 -182.755 ;
        RECT 124.955 -184.445 125.285 -184.115 ;
        RECT 124.955 -185.805 125.285 -185.475 ;
        RECT 124.955 -187.165 125.285 -186.835 ;
        RECT 124.955 -188.525 125.285 -188.195 ;
        RECT 124.955 -189.885 125.285 -189.555 ;
        RECT 124.955 -191.245 125.285 -190.915 ;
        RECT 124.955 -192.605 125.285 -192.275 ;
        RECT 124.955 -193.965 125.285 -193.635 ;
        RECT 124.955 -195.325 125.285 -194.995 ;
        RECT 124.955 -196.685 125.285 -196.355 ;
        RECT 124.955 -198.045 125.285 -197.715 ;
        RECT 124.955 -199.405 125.285 -199.075 ;
        RECT 124.955 -200.765 125.285 -200.435 ;
        RECT 124.955 -202.125 125.285 -201.795 ;
        RECT 124.955 -203.485 125.285 -203.155 ;
        RECT 124.955 -204.845 125.285 -204.515 ;
        RECT 124.955 -206.205 125.285 -205.875 ;
        RECT 124.955 -207.565 125.285 -207.235 ;
        RECT 124.955 -208.925 125.285 -208.595 ;
        RECT 124.955 -210.285 125.285 -209.955 ;
        RECT 124.955 -211.645 125.285 -211.315 ;
        RECT 124.955 -213.005 125.285 -212.675 ;
        RECT 124.955 -214.365 125.285 -214.035 ;
        RECT 124.955 -215.725 125.285 -215.395 ;
        RECT 124.955 -217.085 125.285 -216.755 ;
        RECT 124.955 -218.445 125.285 -218.115 ;
        RECT 124.955 -224.09 125.285 -222.96 ;
        RECT 124.96 -224.205 125.28 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.315 132.52 126.645 133.65 ;
        RECT 126.315 128.355 126.645 128.685 ;
        RECT 126.315 126.995 126.645 127.325 ;
        RECT 126.315 125.635 126.645 125.965 ;
        RECT 126.315 124.275 126.645 124.605 ;
        RECT 126.32 123.6 126.64 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.315 -0.845 126.645 -0.515 ;
        RECT 126.315 -2.205 126.645 -1.875 ;
        RECT 126.315 -3.565 126.645 -3.235 ;
        RECT 126.32 -3.565 126.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.675 132.52 128.005 133.65 ;
        RECT 127.675 128.355 128.005 128.685 ;
        RECT 127.675 126.995 128.005 127.325 ;
        RECT 127.675 125.635 128.005 125.965 ;
        RECT 127.675 124.275 128.005 124.605 ;
        RECT 127.68 123.6 128 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.675 -0.845 128.005 -0.515 ;
        RECT 127.675 -2.205 128.005 -1.875 ;
        RECT 127.675 -3.565 128.005 -3.235 ;
        RECT 127.68 -3.565 128 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.035 132.52 129.365 133.65 ;
        RECT 129.035 128.355 129.365 128.685 ;
        RECT 129.035 126.995 129.365 127.325 ;
        RECT 129.035 125.635 129.365 125.965 ;
        RECT 129.035 124.275 129.365 124.605 ;
        RECT 129.04 123.6 129.36 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.035 -0.845 129.365 -0.515 ;
        RECT 129.035 -2.205 129.365 -1.875 ;
        RECT 129.035 -3.565 129.365 -3.235 ;
        RECT 129.04 -3.565 129.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.035 -119.165 129.365 -118.835 ;
        RECT 129.035 -120.525 129.365 -120.195 ;
        RECT 129.035 -121.885 129.365 -121.555 ;
        RECT 129.035 -123.245 129.365 -122.915 ;
        RECT 129.035 -124.605 129.365 -124.275 ;
        RECT 129.035 -125.965 129.365 -125.635 ;
        RECT 129.035 -127.325 129.365 -126.995 ;
        RECT 129.035 -128.685 129.365 -128.355 ;
        RECT 129.035 -130.045 129.365 -129.715 ;
        RECT 129.035 -131.405 129.365 -131.075 ;
        RECT 129.035 -132.765 129.365 -132.435 ;
        RECT 129.035 -134.125 129.365 -133.795 ;
        RECT 129.035 -135.485 129.365 -135.155 ;
        RECT 129.035 -136.845 129.365 -136.515 ;
        RECT 129.035 -138.205 129.365 -137.875 ;
        RECT 129.035 -139.565 129.365 -139.235 ;
        RECT 129.035 -140.925 129.365 -140.595 ;
        RECT 129.035 -142.285 129.365 -141.955 ;
        RECT 129.035 -143.645 129.365 -143.315 ;
        RECT 129.035 -145.005 129.365 -144.675 ;
        RECT 129.035 -146.365 129.365 -146.035 ;
        RECT 129.035 -147.725 129.365 -147.395 ;
        RECT 129.035 -149.085 129.365 -148.755 ;
        RECT 129.035 -150.445 129.365 -150.115 ;
        RECT 129.035 -151.805 129.365 -151.475 ;
        RECT 129.035 -153.165 129.365 -152.835 ;
        RECT 129.035 -154.525 129.365 -154.195 ;
        RECT 129.035 -155.885 129.365 -155.555 ;
        RECT 129.035 -157.245 129.365 -156.915 ;
        RECT 129.035 -158.605 129.365 -158.275 ;
        RECT 129.035 -159.965 129.365 -159.635 ;
        RECT 129.035 -161.325 129.365 -160.995 ;
        RECT 129.035 -162.685 129.365 -162.355 ;
        RECT 129.035 -164.045 129.365 -163.715 ;
        RECT 129.035 -165.405 129.365 -165.075 ;
        RECT 129.035 -166.765 129.365 -166.435 ;
        RECT 129.035 -168.125 129.365 -167.795 ;
        RECT 129.035 -169.485 129.365 -169.155 ;
        RECT 129.035 -170.845 129.365 -170.515 ;
        RECT 129.035 -172.205 129.365 -171.875 ;
        RECT 129.035 -173.565 129.365 -173.235 ;
        RECT 129.035 -174.925 129.365 -174.595 ;
        RECT 129.035 -176.285 129.365 -175.955 ;
        RECT 129.035 -177.645 129.365 -177.315 ;
        RECT 129.035 -179.005 129.365 -178.675 ;
        RECT 129.035 -180.365 129.365 -180.035 ;
        RECT 129.035 -181.725 129.365 -181.395 ;
        RECT 129.035 -183.085 129.365 -182.755 ;
        RECT 129.035 -184.445 129.365 -184.115 ;
        RECT 129.035 -185.805 129.365 -185.475 ;
        RECT 129.035 -187.165 129.365 -186.835 ;
        RECT 129.035 -188.525 129.365 -188.195 ;
        RECT 129.035 -189.885 129.365 -189.555 ;
        RECT 129.035 -191.245 129.365 -190.915 ;
        RECT 129.035 -192.605 129.365 -192.275 ;
        RECT 129.035 -193.965 129.365 -193.635 ;
        RECT 129.035 -195.325 129.365 -194.995 ;
        RECT 129.035 -196.685 129.365 -196.355 ;
        RECT 129.035 -198.045 129.365 -197.715 ;
        RECT 129.035 -199.405 129.365 -199.075 ;
        RECT 129.035 -200.765 129.365 -200.435 ;
        RECT 129.035 -202.125 129.365 -201.795 ;
        RECT 129.035 -203.485 129.365 -203.155 ;
        RECT 129.035 -204.845 129.365 -204.515 ;
        RECT 129.035 -206.205 129.365 -205.875 ;
        RECT 129.035 -207.565 129.365 -207.235 ;
        RECT 129.035 -208.925 129.365 -208.595 ;
        RECT 129.035 -210.285 129.365 -209.955 ;
        RECT 129.035 -211.645 129.365 -211.315 ;
        RECT 129.035 -213.005 129.365 -212.675 ;
        RECT 129.035 -214.365 129.365 -214.035 ;
        RECT 129.035 -215.725 129.365 -215.395 ;
        RECT 129.035 -217.085 129.365 -216.755 ;
        RECT 129.035 -218.445 129.365 -218.115 ;
        RECT 129.035 -224.09 129.365 -222.96 ;
        RECT 129.04 -224.205 129.36 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.395 132.52 130.725 133.65 ;
        RECT 130.395 128.355 130.725 128.685 ;
        RECT 130.395 126.995 130.725 127.325 ;
        RECT 130.395 125.635 130.725 125.965 ;
        RECT 130.395 124.275 130.725 124.605 ;
        RECT 130.4 123.6 130.72 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.395 -123.245 130.725 -122.915 ;
        RECT 130.395 -124.605 130.725 -124.275 ;
        RECT 130.395 -125.965 130.725 -125.635 ;
        RECT 130.395 -127.325 130.725 -126.995 ;
        RECT 130.395 -128.685 130.725 -128.355 ;
        RECT 130.395 -130.045 130.725 -129.715 ;
        RECT 130.395 -131.405 130.725 -131.075 ;
        RECT 130.395 -132.765 130.725 -132.435 ;
        RECT 130.395 -134.125 130.725 -133.795 ;
        RECT 130.395 -135.485 130.725 -135.155 ;
        RECT 130.395 -136.845 130.725 -136.515 ;
        RECT 130.395 -138.205 130.725 -137.875 ;
        RECT 130.395 -139.565 130.725 -139.235 ;
        RECT 130.395 -140.925 130.725 -140.595 ;
        RECT 130.395 -142.285 130.725 -141.955 ;
        RECT 130.395 -143.645 130.725 -143.315 ;
        RECT 130.395 -145.005 130.725 -144.675 ;
        RECT 130.395 -146.365 130.725 -146.035 ;
        RECT 130.395 -147.725 130.725 -147.395 ;
        RECT 130.395 -149.085 130.725 -148.755 ;
        RECT 130.395 -150.445 130.725 -150.115 ;
        RECT 130.395 -151.805 130.725 -151.475 ;
        RECT 130.395 -153.165 130.725 -152.835 ;
        RECT 130.395 -154.525 130.725 -154.195 ;
        RECT 130.395 -155.885 130.725 -155.555 ;
        RECT 130.395 -157.245 130.725 -156.915 ;
        RECT 130.395 -158.605 130.725 -158.275 ;
        RECT 130.395 -159.965 130.725 -159.635 ;
        RECT 130.395 -161.325 130.725 -160.995 ;
        RECT 130.395 -162.685 130.725 -162.355 ;
        RECT 130.395 -164.045 130.725 -163.715 ;
        RECT 130.395 -165.405 130.725 -165.075 ;
        RECT 130.395 -166.765 130.725 -166.435 ;
        RECT 130.395 -168.125 130.725 -167.795 ;
        RECT 130.395 -169.485 130.725 -169.155 ;
        RECT 130.395 -170.845 130.725 -170.515 ;
        RECT 130.395 -172.205 130.725 -171.875 ;
        RECT 130.395 -173.565 130.725 -173.235 ;
        RECT 130.395 -174.925 130.725 -174.595 ;
        RECT 130.395 -176.285 130.725 -175.955 ;
        RECT 130.395 -177.645 130.725 -177.315 ;
        RECT 130.395 -179.005 130.725 -178.675 ;
        RECT 130.395 -180.365 130.725 -180.035 ;
        RECT 130.395 -181.725 130.725 -181.395 ;
        RECT 130.395 -183.085 130.725 -182.755 ;
        RECT 130.395 -184.445 130.725 -184.115 ;
        RECT 130.395 -185.805 130.725 -185.475 ;
        RECT 130.395 -187.165 130.725 -186.835 ;
        RECT 130.395 -188.525 130.725 -188.195 ;
        RECT 130.395 -189.885 130.725 -189.555 ;
        RECT 130.395 -191.245 130.725 -190.915 ;
        RECT 130.395 -192.605 130.725 -192.275 ;
        RECT 130.395 -193.965 130.725 -193.635 ;
        RECT 130.395 -195.325 130.725 -194.995 ;
        RECT 130.395 -196.685 130.725 -196.355 ;
        RECT 130.395 -198.045 130.725 -197.715 ;
        RECT 130.395 -199.405 130.725 -199.075 ;
        RECT 130.395 -200.765 130.725 -200.435 ;
        RECT 130.395 -202.125 130.725 -201.795 ;
        RECT 130.395 -203.485 130.725 -203.155 ;
        RECT 130.395 -204.845 130.725 -204.515 ;
        RECT 130.395 -206.205 130.725 -205.875 ;
        RECT 130.395 -207.565 130.725 -207.235 ;
        RECT 130.395 -208.925 130.725 -208.595 ;
        RECT 130.395 -210.285 130.725 -209.955 ;
        RECT 130.395 -211.645 130.725 -211.315 ;
        RECT 130.395 -213.005 130.725 -212.675 ;
        RECT 130.395 -214.365 130.725 -214.035 ;
        RECT 130.395 -215.725 130.725 -215.395 ;
        RECT 130.395 -217.085 130.725 -216.755 ;
        RECT 130.395 -218.445 130.725 -218.115 ;
        RECT 130.395 -224.09 130.725 -222.96 ;
        RECT 130.4 -224.205 130.72 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.76 -121.535 131.09 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.755 132.52 132.085 133.65 ;
        RECT 131.755 128.355 132.085 128.685 ;
        RECT 131.755 126.995 132.085 127.325 ;
        RECT 131.755 125.635 132.085 125.965 ;
        RECT 131.755 124.275 132.085 124.605 ;
        RECT 131.76 123.6 132.08 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.115 132.52 133.445 133.65 ;
        RECT 133.115 128.355 133.445 128.685 ;
        RECT 133.115 126.995 133.445 127.325 ;
        RECT 133.115 125.635 133.445 125.965 ;
        RECT 133.115 124.275 133.445 124.605 ;
        RECT 133.12 123.6 133.44 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.115 -0.845 133.445 -0.515 ;
        RECT 133.115 -2.205 133.445 -1.875 ;
        RECT 133.115 -3.565 133.445 -3.235 ;
        RECT 133.12 -3.565 133.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.475 132.52 134.805 133.65 ;
        RECT 134.475 128.355 134.805 128.685 ;
        RECT 134.475 126.995 134.805 127.325 ;
        RECT 134.475 125.635 134.805 125.965 ;
        RECT 134.475 124.275 134.805 124.605 ;
        RECT 134.48 123.6 134.8 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.475 -0.845 134.805 -0.515 ;
        RECT 134.475 -2.205 134.805 -1.875 ;
        RECT 134.475 -3.565 134.805 -3.235 ;
        RECT 134.48 -3.565 134.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.475 -119.165 134.805 -118.835 ;
        RECT 134.475 -120.525 134.805 -120.195 ;
        RECT 134.475 -121.885 134.805 -121.555 ;
        RECT 134.475 -123.245 134.805 -122.915 ;
        RECT 134.475 -124.605 134.805 -124.275 ;
        RECT 134.475 -125.965 134.805 -125.635 ;
        RECT 134.475 -127.325 134.805 -126.995 ;
        RECT 134.475 -128.685 134.805 -128.355 ;
        RECT 134.475 -130.045 134.805 -129.715 ;
        RECT 134.475 -131.405 134.805 -131.075 ;
        RECT 134.475 -132.765 134.805 -132.435 ;
        RECT 134.475 -134.125 134.805 -133.795 ;
        RECT 134.475 -135.485 134.805 -135.155 ;
        RECT 134.475 -136.845 134.805 -136.515 ;
        RECT 134.475 -138.205 134.805 -137.875 ;
        RECT 134.475 -139.565 134.805 -139.235 ;
        RECT 134.475 -140.925 134.805 -140.595 ;
        RECT 134.475 -142.285 134.805 -141.955 ;
        RECT 134.475 -143.645 134.805 -143.315 ;
        RECT 134.475 -145.005 134.805 -144.675 ;
        RECT 134.475 -146.365 134.805 -146.035 ;
        RECT 134.475 -147.725 134.805 -147.395 ;
        RECT 134.475 -149.085 134.805 -148.755 ;
        RECT 134.475 -150.445 134.805 -150.115 ;
        RECT 134.475 -151.805 134.805 -151.475 ;
        RECT 134.475 -153.165 134.805 -152.835 ;
        RECT 134.475 -154.525 134.805 -154.195 ;
        RECT 134.475 -155.885 134.805 -155.555 ;
        RECT 134.475 -157.245 134.805 -156.915 ;
        RECT 134.475 -158.605 134.805 -158.275 ;
        RECT 134.475 -159.965 134.805 -159.635 ;
        RECT 134.475 -161.325 134.805 -160.995 ;
        RECT 134.475 -162.685 134.805 -162.355 ;
        RECT 134.475 -164.045 134.805 -163.715 ;
        RECT 134.475 -165.405 134.805 -165.075 ;
        RECT 134.475 -166.765 134.805 -166.435 ;
        RECT 134.475 -168.125 134.805 -167.795 ;
        RECT 134.475 -169.485 134.805 -169.155 ;
        RECT 134.475 -170.845 134.805 -170.515 ;
        RECT 134.475 -172.205 134.805 -171.875 ;
        RECT 134.475 -173.565 134.805 -173.235 ;
        RECT 134.475 -174.925 134.805 -174.595 ;
        RECT 134.475 -176.285 134.805 -175.955 ;
        RECT 134.475 -177.645 134.805 -177.315 ;
        RECT 134.475 -179.005 134.805 -178.675 ;
        RECT 134.475 -180.365 134.805 -180.035 ;
        RECT 134.475 -181.725 134.805 -181.395 ;
        RECT 134.475 -183.085 134.805 -182.755 ;
        RECT 134.475 -184.445 134.805 -184.115 ;
        RECT 134.475 -185.805 134.805 -185.475 ;
        RECT 134.475 -187.165 134.805 -186.835 ;
        RECT 134.475 -188.525 134.805 -188.195 ;
        RECT 134.475 -189.885 134.805 -189.555 ;
        RECT 134.475 -191.245 134.805 -190.915 ;
        RECT 134.475 -192.605 134.805 -192.275 ;
        RECT 134.475 -193.965 134.805 -193.635 ;
        RECT 134.475 -195.325 134.805 -194.995 ;
        RECT 134.475 -196.685 134.805 -196.355 ;
        RECT 134.475 -198.045 134.805 -197.715 ;
        RECT 134.475 -199.405 134.805 -199.075 ;
        RECT 134.475 -200.765 134.805 -200.435 ;
        RECT 134.475 -202.125 134.805 -201.795 ;
        RECT 134.475 -203.485 134.805 -203.155 ;
        RECT 134.475 -204.845 134.805 -204.515 ;
        RECT 134.475 -206.205 134.805 -205.875 ;
        RECT 134.475 -207.565 134.805 -207.235 ;
        RECT 134.475 -208.925 134.805 -208.595 ;
        RECT 134.475 -210.285 134.805 -209.955 ;
        RECT 134.475 -211.645 134.805 -211.315 ;
        RECT 134.475 -213.005 134.805 -212.675 ;
        RECT 134.475 -214.365 134.805 -214.035 ;
        RECT 134.475 -215.725 134.805 -215.395 ;
        RECT 134.475 -217.085 134.805 -216.755 ;
        RECT 134.475 -218.445 134.805 -218.115 ;
        RECT 134.475 -224.09 134.805 -222.96 ;
        RECT 134.48 -224.205 134.8 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.835 132.52 136.165 133.65 ;
        RECT 135.835 128.355 136.165 128.685 ;
        RECT 135.835 126.995 136.165 127.325 ;
        RECT 135.835 125.635 136.165 125.965 ;
        RECT 135.835 124.275 136.165 124.605 ;
        RECT 135.84 123.6 136.16 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.835 -0.845 136.165 -0.515 ;
        RECT 135.835 -2.205 136.165 -1.875 ;
        RECT 135.835 -3.565 136.165 -3.235 ;
        RECT 135.84 -3.565 136.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.835 -195.325 136.165 -194.995 ;
        RECT 135.835 -196.685 136.165 -196.355 ;
        RECT 135.835 -198.045 136.165 -197.715 ;
        RECT 135.835 -199.405 136.165 -199.075 ;
        RECT 135.835 -200.765 136.165 -200.435 ;
        RECT 135.835 -202.125 136.165 -201.795 ;
        RECT 135.835 -203.485 136.165 -203.155 ;
        RECT 135.835 -204.845 136.165 -204.515 ;
        RECT 135.835 -206.205 136.165 -205.875 ;
        RECT 135.835 -207.565 136.165 -207.235 ;
        RECT 135.835 -208.925 136.165 -208.595 ;
        RECT 135.835 -210.285 136.165 -209.955 ;
        RECT 135.835 -211.645 136.165 -211.315 ;
        RECT 135.835 -213.005 136.165 -212.675 ;
        RECT 135.835 -214.365 136.165 -214.035 ;
        RECT 135.835 -215.725 136.165 -215.395 ;
        RECT 135.835 -217.085 136.165 -216.755 ;
        RECT 135.835 -218.445 136.165 -218.115 ;
        RECT 135.835 -224.09 136.165 -222.96 ;
        RECT 135.84 -224.205 136.16 -118.16 ;
        RECT 135.835 -119.165 136.165 -118.835 ;
        RECT 135.835 -120.525 136.165 -120.195 ;
        RECT 135.835 -121.885 136.165 -121.555 ;
        RECT 135.835 -123.245 136.165 -122.915 ;
        RECT 135.835 -124.605 136.165 -124.275 ;
        RECT 135.835 -125.965 136.165 -125.635 ;
        RECT 135.835 -127.325 136.165 -126.995 ;
        RECT 135.835 -128.685 136.165 -128.355 ;
        RECT 135.835 -130.045 136.165 -129.715 ;
        RECT 135.835 -131.405 136.165 -131.075 ;
        RECT 135.835 -132.765 136.165 -132.435 ;
        RECT 135.835 -134.125 136.165 -133.795 ;
        RECT 135.835 -135.485 136.165 -135.155 ;
        RECT 135.835 -136.845 136.165 -136.515 ;
        RECT 135.835 -138.205 136.165 -137.875 ;
        RECT 135.835 -139.565 136.165 -139.235 ;
        RECT 135.835 -140.925 136.165 -140.595 ;
        RECT 135.835 -142.285 136.165 -141.955 ;
        RECT 135.835 -143.645 136.165 -143.315 ;
        RECT 135.835 -145.005 136.165 -144.675 ;
        RECT 135.835 -146.365 136.165 -146.035 ;
        RECT 135.835 -147.725 136.165 -147.395 ;
        RECT 135.835 -149.085 136.165 -148.755 ;
        RECT 135.835 -150.445 136.165 -150.115 ;
        RECT 135.835 -151.805 136.165 -151.475 ;
        RECT 135.835 -153.165 136.165 -152.835 ;
        RECT 135.835 -154.525 136.165 -154.195 ;
        RECT 135.835 -155.885 136.165 -155.555 ;
        RECT 135.835 -157.245 136.165 -156.915 ;
        RECT 135.835 -158.605 136.165 -158.275 ;
        RECT 135.835 -159.965 136.165 -159.635 ;
        RECT 135.835 -161.325 136.165 -160.995 ;
        RECT 135.835 -162.685 136.165 -162.355 ;
        RECT 135.835 -164.045 136.165 -163.715 ;
        RECT 135.835 -165.405 136.165 -165.075 ;
        RECT 135.835 -166.765 136.165 -166.435 ;
        RECT 135.835 -168.125 136.165 -167.795 ;
        RECT 135.835 -169.485 136.165 -169.155 ;
        RECT 135.835 -170.845 136.165 -170.515 ;
        RECT 135.835 -172.205 136.165 -171.875 ;
        RECT 135.835 -173.565 136.165 -173.235 ;
        RECT 135.835 -174.925 136.165 -174.595 ;
        RECT 135.835 -176.285 136.165 -175.955 ;
        RECT 135.835 -177.645 136.165 -177.315 ;
        RECT 135.835 -179.005 136.165 -178.675 ;
        RECT 135.835 -180.365 136.165 -180.035 ;
        RECT 135.835 -181.725 136.165 -181.395 ;
        RECT 135.835 -183.085 136.165 -182.755 ;
        RECT 135.835 -184.445 136.165 -184.115 ;
        RECT 135.835 -185.805 136.165 -185.475 ;
        RECT 135.835 -187.165 136.165 -186.835 ;
        RECT 135.835 -188.525 136.165 -188.195 ;
        RECT 135.835 -189.885 136.165 -189.555 ;
        RECT 135.835 -191.245 136.165 -190.915 ;
        RECT 135.835 -192.605 136.165 -192.275 ;
        RECT 135.835 -193.965 136.165 -193.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.86 -121.535 76.19 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.995 132.52 76.325 133.65 ;
        RECT 75.995 128.355 76.325 128.685 ;
        RECT 75.995 126.995 76.325 127.325 ;
        RECT 75.995 125.635 76.325 125.965 ;
        RECT 75.995 124.275 76.325 124.605 ;
        RECT 76 123.6 76.32 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.995 -123.245 76.325 -122.915 ;
        RECT 75.995 -124.605 76.325 -124.275 ;
        RECT 75.995 -125.965 76.325 -125.635 ;
        RECT 75.995 -127.325 76.325 -126.995 ;
        RECT 75.995 -128.685 76.325 -128.355 ;
        RECT 75.995 -130.045 76.325 -129.715 ;
        RECT 75.995 -131.405 76.325 -131.075 ;
        RECT 75.995 -132.765 76.325 -132.435 ;
        RECT 75.995 -134.125 76.325 -133.795 ;
        RECT 75.995 -135.485 76.325 -135.155 ;
        RECT 75.995 -136.845 76.325 -136.515 ;
        RECT 75.995 -138.205 76.325 -137.875 ;
        RECT 75.995 -139.565 76.325 -139.235 ;
        RECT 75.995 -140.925 76.325 -140.595 ;
        RECT 75.995 -142.285 76.325 -141.955 ;
        RECT 75.995 -143.645 76.325 -143.315 ;
        RECT 75.995 -145.005 76.325 -144.675 ;
        RECT 75.995 -146.365 76.325 -146.035 ;
        RECT 75.995 -147.725 76.325 -147.395 ;
        RECT 75.995 -149.085 76.325 -148.755 ;
        RECT 75.995 -150.445 76.325 -150.115 ;
        RECT 75.995 -151.805 76.325 -151.475 ;
        RECT 75.995 -153.165 76.325 -152.835 ;
        RECT 75.995 -154.525 76.325 -154.195 ;
        RECT 75.995 -155.885 76.325 -155.555 ;
        RECT 75.995 -157.245 76.325 -156.915 ;
        RECT 75.995 -158.605 76.325 -158.275 ;
        RECT 75.995 -159.965 76.325 -159.635 ;
        RECT 75.995 -161.325 76.325 -160.995 ;
        RECT 75.995 -162.685 76.325 -162.355 ;
        RECT 75.995 -164.045 76.325 -163.715 ;
        RECT 75.995 -165.405 76.325 -165.075 ;
        RECT 75.995 -166.765 76.325 -166.435 ;
        RECT 75.995 -168.125 76.325 -167.795 ;
        RECT 75.995 -169.485 76.325 -169.155 ;
        RECT 75.995 -170.845 76.325 -170.515 ;
        RECT 75.995 -172.205 76.325 -171.875 ;
        RECT 75.995 -173.565 76.325 -173.235 ;
        RECT 75.995 -174.925 76.325 -174.595 ;
        RECT 75.995 -176.285 76.325 -175.955 ;
        RECT 75.995 -177.645 76.325 -177.315 ;
        RECT 75.995 -179.005 76.325 -178.675 ;
        RECT 75.995 -180.365 76.325 -180.035 ;
        RECT 75.995 -181.725 76.325 -181.395 ;
        RECT 75.995 -183.085 76.325 -182.755 ;
        RECT 75.995 -184.445 76.325 -184.115 ;
        RECT 75.995 -185.805 76.325 -185.475 ;
        RECT 75.995 -187.165 76.325 -186.835 ;
        RECT 75.995 -188.525 76.325 -188.195 ;
        RECT 75.995 -189.885 76.325 -189.555 ;
        RECT 75.995 -191.245 76.325 -190.915 ;
        RECT 75.995 -192.605 76.325 -192.275 ;
        RECT 75.995 -193.965 76.325 -193.635 ;
        RECT 75.995 -195.325 76.325 -194.995 ;
        RECT 75.995 -196.685 76.325 -196.355 ;
        RECT 75.995 -198.045 76.325 -197.715 ;
        RECT 75.995 -199.405 76.325 -199.075 ;
        RECT 75.995 -200.765 76.325 -200.435 ;
        RECT 75.995 -202.125 76.325 -201.795 ;
        RECT 75.995 -203.485 76.325 -203.155 ;
        RECT 75.995 -204.845 76.325 -204.515 ;
        RECT 75.995 -206.205 76.325 -205.875 ;
        RECT 75.995 -207.565 76.325 -207.235 ;
        RECT 75.995 -208.925 76.325 -208.595 ;
        RECT 75.995 -210.285 76.325 -209.955 ;
        RECT 75.995 -211.645 76.325 -211.315 ;
        RECT 75.995 -213.005 76.325 -212.675 ;
        RECT 75.995 -214.365 76.325 -214.035 ;
        RECT 75.995 -215.725 76.325 -215.395 ;
        RECT 75.995 -217.085 76.325 -216.755 ;
        RECT 75.995 -218.445 76.325 -218.115 ;
        RECT 75.995 -224.09 76.325 -222.96 ;
        RECT 76 -224.205 76.32 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.355 132.52 77.685 133.65 ;
        RECT 77.355 128.355 77.685 128.685 ;
        RECT 77.355 126.995 77.685 127.325 ;
        RECT 77.355 125.635 77.685 125.965 ;
        RECT 77.355 124.275 77.685 124.605 ;
        RECT 77.36 123.6 77.68 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.355 -0.845 77.685 -0.515 ;
        RECT 77.355 -2.205 77.685 -1.875 ;
        RECT 77.355 -3.565 77.685 -3.235 ;
        RECT 77.36 -3.565 77.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.715 132.52 79.045 133.65 ;
        RECT 78.715 128.355 79.045 128.685 ;
        RECT 78.715 126.995 79.045 127.325 ;
        RECT 78.715 125.635 79.045 125.965 ;
        RECT 78.715 124.275 79.045 124.605 ;
        RECT 78.72 123.6 79.04 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.715 -0.845 79.045 -0.515 ;
        RECT 78.715 -2.205 79.045 -1.875 ;
        RECT 78.715 -3.565 79.045 -3.235 ;
        RECT 78.72 -3.565 79.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.075 132.52 80.405 133.65 ;
        RECT 80.075 128.355 80.405 128.685 ;
        RECT 80.075 126.995 80.405 127.325 ;
        RECT 80.075 125.635 80.405 125.965 ;
        RECT 80.075 124.275 80.405 124.605 ;
        RECT 80.08 123.6 80.4 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.075 -0.845 80.405 -0.515 ;
        RECT 80.075 -2.205 80.405 -1.875 ;
        RECT 80.075 -3.565 80.405 -3.235 ;
        RECT 80.08 -3.565 80.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.075 -119.165 80.405 -118.835 ;
        RECT 80.075 -120.525 80.405 -120.195 ;
        RECT 80.075 -121.885 80.405 -121.555 ;
        RECT 80.075 -123.245 80.405 -122.915 ;
        RECT 80.075 -124.605 80.405 -124.275 ;
        RECT 80.075 -125.965 80.405 -125.635 ;
        RECT 80.075 -127.325 80.405 -126.995 ;
        RECT 80.075 -128.685 80.405 -128.355 ;
        RECT 80.075 -130.045 80.405 -129.715 ;
        RECT 80.075 -131.405 80.405 -131.075 ;
        RECT 80.075 -132.765 80.405 -132.435 ;
        RECT 80.075 -134.125 80.405 -133.795 ;
        RECT 80.075 -135.485 80.405 -135.155 ;
        RECT 80.075 -136.845 80.405 -136.515 ;
        RECT 80.075 -138.205 80.405 -137.875 ;
        RECT 80.075 -139.565 80.405 -139.235 ;
        RECT 80.075 -140.925 80.405 -140.595 ;
        RECT 80.075 -142.285 80.405 -141.955 ;
        RECT 80.075 -143.645 80.405 -143.315 ;
        RECT 80.075 -145.005 80.405 -144.675 ;
        RECT 80.075 -146.365 80.405 -146.035 ;
        RECT 80.075 -147.725 80.405 -147.395 ;
        RECT 80.075 -149.085 80.405 -148.755 ;
        RECT 80.075 -150.445 80.405 -150.115 ;
        RECT 80.075 -151.805 80.405 -151.475 ;
        RECT 80.075 -153.165 80.405 -152.835 ;
        RECT 80.075 -154.525 80.405 -154.195 ;
        RECT 80.075 -155.885 80.405 -155.555 ;
        RECT 80.075 -157.245 80.405 -156.915 ;
        RECT 80.075 -158.605 80.405 -158.275 ;
        RECT 80.075 -159.965 80.405 -159.635 ;
        RECT 80.075 -161.325 80.405 -160.995 ;
        RECT 80.075 -162.685 80.405 -162.355 ;
        RECT 80.075 -164.045 80.405 -163.715 ;
        RECT 80.075 -165.405 80.405 -165.075 ;
        RECT 80.075 -166.765 80.405 -166.435 ;
        RECT 80.075 -168.125 80.405 -167.795 ;
        RECT 80.075 -169.485 80.405 -169.155 ;
        RECT 80.075 -170.845 80.405 -170.515 ;
        RECT 80.075 -172.205 80.405 -171.875 ;
        RECT 80.075 -173.565 80.405 -173.235 ;
        RECT 80.075 -174.925 80.405 -174.595 ;
        RECT 80.075 -176.285 80.405 -175.955 ;
        RECT 80.075 -177.645 80.405 -177.315 ;
        RECT 80.075 -179.005 80.405 -178.675 ;
        RECT 80.075 -180.365 80.405 -180.035 ;
        RECT 80.075 -181.725 80.405 -181.395 ;
        RECT 80.075 -183.085 80.405 -182.755 ;
        RECT 80.075 -184.445 80.405 -184.115 ;
        RECT 80.075 -185.805 80.405 -185.475 ;
        RECT 80.075 -187.165 80.405 -186.835 ;
        RECT 80.075 -188.525 80.405 -188.195 ;
        RECT 80.075 -189.885 80.405 -189.555 ;
        RECT 80.075 -191.245 80.405 -190.915 ;
        RECT 80.075 -192.605 80.405 -192.275 ;
        RECT 80.075 -193.965 80.405 -193.635 ;
        RECT 80.075 -195.325 80.405 -194.995 ;
        RECT 80.075 -196.685 80.405 -196.355 ;
        RECT 80.075 -198.045 80.405 -197.715 ;
        RECT 80.075 -199.405 80.405 -199.075 ;
        RECT 80.075 -200.765 80.405 -200.435 ;
        RECT 80.075 -202.125 80.405 -201.795 ;
        RECT 80.075 -203.485 80.405 -203.155 ;
        RECT 80.075 -204.845 80.405 -204.515 ;
        RECT 80.075 -206.205 80.405 -205.875 ;
        RECT 80.075 -207.565 80.405 -207.235 ;
        RECT 80.075 -208.925 80.405 -208.595 ;
        RECT 80.075 -210.285 80.405 -209.955 ;
        RECT 80.075 -211.645 80.405 -211.315 ;
        RECT 80.075 -213.005 80.405 -212.675 ;
        RECT 80.075 -214.365 80.405 -214.035 ;
        RECT 80.075 -215.725 80.405 -215.395 ;
        RECT 80.075 -217.085 80.405 -216.755 ;
        RECT 80.075 -218.445 80.405 -218.115 ;
        RECT 80.075 -224.09 80.405 -222.96 ;
        RECT 80.08 -224.205 80.4 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.435 132.52 81.765 133.65 ;
        RECT 81.435 128.355 81.765 128.685 ;
        RECT 81.435 126.995 81.765 127.325 ;
        RECT 81.435 125.635 81.765 125.965 ;
        RECT 81.435 124.275 81.765 124.605 ;
        RECT 81.44 123.6 81.76 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.435 -123.245 81.765 -122.915 ;
        RECT 81.435 -124.605 81.765 -124.275 ;
        RECT 81.435 -125.965 81.765 -125.635 ;
        RECT 81.435 -127.325 81.765 -126.995 ;
        RECT 81.435 -128.685 81.765 -128.355 ;
        RECT 81.435 -130.045 81.765 -129.715 ;
        RECT 81.435 -131.405 81.765 -131.075 ;
        RECT 81.435 -132.765 81.765 -132.435 ;
        RECT 81.435 -134.125 81.765 -133.795 ;
        RECT 81.435 -135.485 81.765 -135.155 ;
        RECT 81.435 -136.845 81.765 -136.515 ;
        RECT 81.435 -138.205 81.765 -137.875 ;
        RECT 81.435 -139.565 81.765 -139.235 ;
        RECT 81.435 -140.925 81.765 -140.595 ;
        RECT 81.435 -142.285 81.765 -141.955 ;
        RECT 81.435 -143.645 81.765 -143.315 ;
        RECT 81.435 -145.005 81.765 -144.675 ;
        RECT 81.435 -146.365 81.765 -146.035 ;
        RECT 81.435 -147.725 81.765 -147.395 ;
        RECT 81.435 -149.085 81.765 -148.755 ;
        RECT 81.435 -150.445 81.765 -150.115 ;
        RECT 81.435 -151.805 81.765 -151.475 ;
        RECT 81.435 -153.165 81.765 -152.835 ;
        RECT 81.435 -154.525 81.765 -154.195 ;
        RECT 81.435 -155.885 81.765 -155.555 ;
        RECT 81.435 -157.245 81.765 -156.915 ;
        RECT 81.435 -158.605 81.765 -158.275 ;
        RECT 81.435 -159.965 81.765 -159.635 ;
        RECT 81.435 -161.325 81.765 -160.995 ;
        RECT 81.435 -162.685 81.765 -162.355 ;
        RECT 81.435 -164.045 81.765 -163.715 ;
        RECT 81.435 -165.405 81.765 -165.075 ;
        RECT 81.435 -166.765 81.765 -166.435 ;
        RECT 81.435 -168.125 81.765 -167.795 ;
        RECT 81.435 -169.485 81.765 -169.155 ;
        RECT 81.435 -170.845 81.765 -170.515 ;
        RECT 81.435 -172.205 81.765 -171.875 ;
        RECT 81.435 -173.565 81.765 -173.235 ;
        RECT 81.435 -174.925 81.765 -174.595 ;
        RECT 81.435 -176.285 81.765 -175.955 ;
        RECT 81.435 -177.645 81.765 -177.315 ;
        RECT 81.435 -179.005 81.765 -178.675 ;
        RECT 81.435 -180.365 81.765 -180.035 ;
        RECT 81.435 -181.725 81.765 -181.395 ;
        RECT 81.435 -183.085 81.765 -182.755 ;
        RECT 81.435 -184.445 81.765 -184.115 ;
        RECT 81.435 -185.805 81.765 -185.475 ;
        RECT 81.435 -187.165 81.765 -186.835 ;
        RECT 81.435 -188.525 81.765 -188.195 ;
        RECT 81.435 -189.885 81.765 -189.555 ;
        RECT 81.435 -191.245 81.765 -190.915 ;
        RECT 81.435 -192.605 81.765 -192.275 ;
        RECT 81.435 -193.965 81.765 -193.635 ;
        RECT 81.435 -195.325 81.765 -194.995 ;
        RECT 81.435 -196.685 81.765 -196.355 ;
        RECT 81.435 -198.045 81.765 -197.715 ;
        RECT 81.435 -199.405 81.765 -199.075 ;
        RECT 81.435 -200.765 81.765 -200.435 ;
        RECT 81.435 -202.125 81.765 -201.795 ;
        RECT 81.435 -203.485 81.765 -203.155 ;
        RECT 81.435 -204.845 81.765 -204.515 ;
        RECT 81.435 -206.205 81.765 -205.875 ;
        RECT 81.435 -207.565 81.765 -207.235 ;
        RECT 81.435 -208.925 81.765 -208.595 ;
        RECT 81.435 -210.285 81.765 -209.955 ;
        RECT 81.435 -211.645 81.765 -211.315 ;
        RECT 81.435 -213.005 81.765 -212.675 ;
        RECT 81.435 -214.365 81.765 -214.035 ;
        RECT 81.435 -215.725 81.765 -215.395 ;
        RECT 81.435 -217.085 81.765 -216.755 ;
        RECT 81.435 -218.445 81.765 -218.115 ;
        RECT 81.435 -224.09 81.765 -222.96 ;
        RECT 81.44 -224.205 81.76 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.96 -121.535 82.29 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.795 132.52 83.125 133.65 ;
        RECT 82.795 128.355 83.125 128.685 ;
        RECT 82.795 126.995 83.125 127.325 ;
        RECT 82.795 125.635 83.125 125.965 ;
        RECT 82.795 124.275 83.125 124.605 ;
        RECT 82.8 123.6 83.12 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.155 132.52 84.485 133.65 ;
        RECT 84.155 128.355 84.485 128.685 ;
        RECT 84.155 126.995 84.485 127.325 ;
        RECT 84.155 125.635 84.485 125.965 ;
        RECT 84.155 124.275 84.485 124.605 ;
        RECT 84.16 123.6 84.48 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.155 -0.845 84.485 -0.515 ;
        RECT 84.155 -2.205 84.485 -1.875 ;
        RECT 84.155 -3.565 84.485 -3.235 ;
        RECT 84.16 -3.565 84.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.155 -119.165 84.485 -118.835 ;
        RECT 84.155 -120.525 84.485 -120.195 ;
        RECT 84.155 -121.885 84.485 -121.555 ;
        RECT 84.155 -123.245 84.485 -122.915 ;
        RECT 84.155 -124.605 84.485 -124.275 ;
        RECT 84.155 -125.965 84.485 -125.635 ;
        RECT 84.155 -127.325 84.485 -126.995 ;
        RECT 84.155 -128.685 84.485 -128.355 ;
        RECT 84.155 -130.045 84.485 -129.715 ;
        RECT 84.155 -131.405 84.485 -131.075 ;
        RECT 84.155 -132.765 84.485 -132.435 ;
        RECT 84.155 -134.125 84.485 -133.795 ;
        RECT 84.155 -135.485 84.485 -135.155 ;
        RECT 84.155 -136.845 84.485 -136.515 ;
        RECT 84.155 -138.205 84.485 -137.875 ;
        RECT 84.155 -139.565 84.485 -139.235 ;
        RECT 84.155 -140.925 84.485 -140.595 ;
        RECT 84.155 -142.285 84.485 -141.955 ;
        RECT 84.155 -143.645 84.485 -143.315 ;
        RECT 84.155 -145.005 84.485 -144.675 ;
        RECT 84.155 -146.365 84.485 -146.035 ;
        RECT 84.155 -147.725 84.485 -147.395 ;
        RECT 84.155 -149.085 84.485 -148.755 ;
        RECT 84.155 -150.445 84.485 -150.115 ;
        RECT 84.155 -151.805 84.485 -151.475 ;
        RECT 84.155 -153.165 84.485 -152.835 ;
        RECT 84.155 -154.525 84.485 -154.195 ;
        RECT 84.155 -155.885 84.485 -155.555 ;
        RECT 84.155 -157.245 84.485 -156.915 ;
        RECT 84.155 -158.605 84.485 -158.275 ;
        RECT 84.155 -159.965 84.485 -159.635 ;
        RECT 84.155 -161.325 84.485 -160.995 ;
        RECT 84.155 -162.685 84.485 -162.355 ;
        RECT 84.155 -164.045 84.485 -163.715 ;
        RECT 84.155 -165.405 84.485 -165.075 ;
        RECT 84.155 -166.765 84.485 -166.435 ;
        RECT 84.155 -168.125 84.485 -167.795 ;
        RECT 84.155 -169.485 84.485 -169.155 ;
        RECT 84.155 -170.845 84.485 -170.515 ;
        RECT 84.155 -172.205 84.485 -171.875 ;
        RECT 84.155 -173.565 84.485 -173.235 ;
        RECT 84.155 -174.925 84.485 -174.595 ;
        RECT 84.155 -176.285 84.485 -175.955 ;
        RECT 84.155 -177.645 84.485 -177.315 ;
        RECT 84.155 -179.005 84.485 -178.675 ;
        RECT 84.155 -180.365 84.485 -180.035 ;
        RECT 84.155 -181.725 84.485 -181.395 ;
        RECT 84.155 -183.085 84.485 -182.755 ;
        RECT 84.155 -184.445 84.485 -184.115 ;
        RECT 84.155 -185.805 84.485 -185.475 ;
        RECT 84.155 -187.165 84.485 -186.835 ;
        RECT 84.155 -188.525 84.485 -188.195 ;
        RECT 84.155 -189.885 84.485 -189.555 ;
        RECT 84.155 -191.245 84.485 -190.915 ;
        RECT 84.155 -192.605 84.485 -192.275 ;
        RECT 84.155 -193.965 84.485 -193.635 ;
        RECT 84.155 -195.325 84.485 -194.995 ;
        RECT 84.155 -196.685 84.485 -196.355 ;
        RECT 84.155 -198.045 84.485 -197.715 ;
        RECT 84.155 -199.405 84.485 -199.075 ;
        RECT 84.155 -200.765 84.485 -200.435 ;
        RECT 84.155 -202.125 84.485 -201.795 ;
        RECT 84.155 -203.485 84.485 -203.155 ;
        RECT 84.155 -204.845 84.485 -204.515 ;
        RECT 84.155 -206.205 84.485 -205.875 ;
        RECT 84.155 -207.565 84.485 -207.235 ;
        RECT 84.155 -208.925 84.485 -208.595 ;
        RECT 84.155 -210.285 84.485 -209.955 ;
        RECT 84.155 -211.645 84.485 -211.315 ;
        RECT 84.155 -213.005 84.485 -212.675 ;
        RECT 84.155 -214.365 84.485 -214.035 ;
        RECT 84.155 -215.725 84.485 -215.395 ;
        RECT 84.155 -217.085 84.485 -216.755 ;
        RECT 84.155 -218.445 84.485 -218.115 ;
        RECT 84.155 -224.09 84.485 -222.96 ;
        RECT 84.16 -224.205 84.48 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.515 132.52 85.845 133.65 ;
        RECT 85.515 128.355 85.845 128.685 ;
        RECT 85.515 126.995 85.845 127.325 ;
        RECT 85.515 125.635 85.845 125.965 ;
        RECT 85.515 124.275 85.845 124.605 ;
        RECT 85.52 123.6 85.84 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.515 -0.845 85.845 -0.515 ;
        RECT 85.515 -2.205 85.845 -1.875 ;
        RECT 85.515 -3.565 85.845 -3.235 ;
        RECT 85.52 -3.565 85.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.875 132.52 87.205 133.65 ;
        RECT 86.875 128.355 87.205 128.685 ;
        RECT 86.875 126.995 87.205 127.325 ;
        RECT 86.875 125.635 87.205 125.965 ;
        RECT 86.875 124.275 87.205 124.605 ;
        RECT 86.88 123.6 87.2 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.875 -0.845 87.205 -0.515 ;
        RECT 86.875 -2.205 87.205 -1.875 ;
        RECT 86.875 -3.565 87.205 -3.235 ;
        RECT 86.88 -3.565 87.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.875 -119.165 87.205 -118.835 ;
        RECT 86.875 -120.525 87.205 -120.195 ;
        RECT 86.875 -121.885 87.205 -121.555 ;
        RECT 86.875 -123.245 87.205 -122.915 ;
        RECT 86.875 -124.605 87.205 -124.275 ;
        RECT 86.875 -125.965 87.205 -125.635 ;
        RECT 86.875 -127.325 87.205 -126.995 ;
        RECT 86.875 -128.685 87.205 -128.355 ;
        RECT 86.875 -130.045 87.205 -129.715 ;
        RECT 86.875 -131.405 87.205 -131.075 ;
        RECT 86.875 -132.765 87.205 -132.435 ;
        RECT 86.875 -134.125 87.205 -133.795 ;
        RECT 86.875 -135.485 87.205 -135.155 ;
        RECT 86.875 -136.845 87.205 -136.515 ;
        RECT 86.875 -138.205 87.205 -137.875 ;
        RECT 86.875 -139.565 87.205 -139.235 ;
        RECT 86.875 -140.925 87.205 -140.595 ;
        RECT 86.875 -142.285 87.205 -141.955 ;
        RECT 86.875 -143.645 87.205 -143.315 ;
        RECT 86.875 -145.005 87.205 -144.675 ;
        RECT 86.875 -146.365 87.205 -146.035 ;
        RECT 86.875 -147.725 87.205 -147.395 ;
        RECT 86.875 -149.085 87.205 -148.755 ;
        RECT 86.875 -150.445 87.205 -150.115 ;
        RECT 86.875 -151.805 87.205 -151.475 ;
        RECT 86.875 -153.165 87.205 -152.835 ;
        RECT 86.875 -154.525 87.205 -154.195 ;
        RECT 86.875 -155.885 87.205 -155.555 ;
        RECT 86.875 -157.245 87.205 -156.915 ;
        RECT 86.875 -158.605 87.205 -158.275 ;
        RECT 86.875 -159.965 87.205 -159.635 ;
        RECT 86.875 -161.325 87.205 -160.995 ;
        RECT 86.875 -162.685 87.205 -162.355 ;
        RECT 86.875 -164.045 87.205 -163.715 ;
        RECT 86.875 -165.405 87.205 -165.075 ;
        RECT 86.875 -166.765 87.205 -166.435 ;
        RECT 86.875 -168.125 87.205 -167.795 ;
        RECT 86.875 -169.485 87.205 -169.155 ;
        RECT 86.875 -170.845 87.205 -170.515 ;
        RECT 86.875 -172.205 87.205 -171.875 ;
        RECT 86.875 -173.565 87.205 -173.235 ;
        RECT 86.875 -174.925 87.205 -174.595 ;
        RECT 86.875 -176.285 87.205 -175.955 ;
        RECT 86.875 -177.645 87.205 -177.315 ;
        RECT 86.875 -179.005 87.205 -178.675 ;
        RECT 86.875 -180.365 87.205 -180.035 ;
        RECT 86.875 -181.725 87.205 -181.395 ;
        RECT 86.875 -183.085 87.205 -182.755 ;
        RECT 86.875 -184.445 87.205 -184.115 ;
        RECT 86.875 -185.805 87.205 -185.475 ;
        RECT 86.875 -187.165 87.205 -186.835 ;
        RECT 86.875 -188.525 87.205 -188.195 ;
        RECT 86.875 -189.885 87.205 -189.555 ;
        RECT 86.875 -191.245 87.205 -190.915 ;
        RECT 86.875 -192.605 87.205 -192.275 ;
        RECT 86.875 -193.965 87.205 -193.635 ;
        RECT 86.875 -195.325 87.205 -194.995 ;
        RECT 86.875 -196.685 87.205 -196.355 ;
        RECT 86.875 -198.045 87.205 -197.715 ;
        RECT 86.875 -199.405 87.205 -199.075 ;
        RECT 86.875 -200.765 87.205 -200.435 ;
        RECT 86.875 -202.125 87.205 -201.795 ;
        RECT 86.875 -203.485 87.205 -203.155 ;
        RECT 86.875 -204.845 87.205 -204.515 ;
        RECT 86.875 -206.205 87.205 -205.875 ;
        RECT 86.875 -207.565 87.205 -207.235 ;
        RECT 86.875 -208.925 87.205 -208.595 ;
        RECT 86.875 -210.285 87.205 -209.955 ;
        RECT 86.875 -211.645 87.205 -211.315 ;
        RECT 86.875 -213.005 87.205 -212.675 ;
        RECT 86.875 -214.365 87.205 -214.035 ;
        RECT 86.875 -215.725 87.205 -215.395 ;
        RECT 86.875 -217.085 87.205 -216.755 ;
        RECT 86.875 -218.445 87.205 -218.115 ;
        RECT 86.875 -224.09 87.205 -222.96 ;
        RECT 86.88 -224.205 87.2 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.06 -121.535 88.39 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.235 132.52 88.565 133.65 ;
        RECT 88.235 128.355 88.565 128.685 ;
        RECT 88.235 126.995 88.565 127.325 ;
        RECT 88.235 125.635 88.565 125.965 ;
        RECT 88.235 124.275 88.565 124.605 ;
        RECT 88.24 123.6 88.56 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.235 -123.245 88.565 -122.915 ;
        RECT 88.235 -124.605 88.565 -124.275 ;
        RECT 88.235 -125.965 88.565 -125.635 ;
        RECT 88.235 -127.325 88.565 -126.995 ;
        RECT 88.235 -128.685 88.565 -128.355 ;
        RECT 88.235 -130.045 88.565 -129.715 ;
        RECT 88.235 -131.405 88.565 -131.075 ;
        RECT 88.235 -132.765 88.565 -132.435 ;
        RECT 88.235 -134.125 88.565 -133.795 ;
        RECT 88.235 -135.485 88.565 -135.155 ;
        RECT 88.235 -136.845 88.565 -136.515 ;
        RECT 88.235 -138.205 88.565 -137.875 ;
        RECT 88.235 -139.565 88.565 -139.235 ;
        RECT 88.235 -140.925 88.565 -140.595 ;
        RECT 88.235 -142.285 88.565 -141.955 ;
        RECT 88.235 -143.645 88.565 -143.315 ;
        RECT 88.235 -145.005 88.565 -144.675 ;
        RECT 88.235 -146.365 88.565 -146.035 ;
        RECT 88.235 -147.725 88.565 -147.395 ;
        RECT 88.235 -149.085 88.565 -148.755 ;
        RECT 88.235 -150.445 88.565 -150.115 ;
        RECT 88.235 -151.805 88.565 -151.475 ;
        RECT 88.235 -153.165 88.565 -152.835 ;
        RECT 88.235 -154.525 88.565 -154.195 ;
        RECT 88.235 -155.885 88.565 -155.555 ;
        RECT 88.235 -157.245 88.565 -156.915 ;
        RECT 88.235 -158.605 88.565 -158.275 ;
        RECT 88.235 -159.965 88.565 -159.635 ;
        RECT 88.235 -161.325 88.565 -160.995 ;
        RECT 88.235 -162.685 88.565 -162.355 ;
        RECT 88.235 -164.045 88.565 -163.715 ;
        RECT 88.235 -165.405 88.565 -165.075 ;
        RECT 88.235 -166.765 88.565 -166.435 ;
        RECT 88.235 -168.125 88.565 -167.795 ;
        RECT 88.235 -169.485 88.565 -169.155 ;
        RECT 88.235 -170.845 88.565 -170.515 ;
        RECT 88.235 -172.205 88.565 -171.875 ;
        RECT 88.235 -173.565 88.565 -173.235 ;
        RECT 88.235 -174.925 88.565 -174.595 ;
        RECT 88.235 -176.285 88.565 -175.955 ;
        RECT 88.235 -177.645 88.565 -177.315 ;
        RECT 88.235 -179.005 88.565 -178.675 ;
        RECT 88.235 -180.365 88.565 -180.035 ;
        RECT 88.235 -181.725 88.565 -181.395 ;
        RECT 88.235 -183.085 88.565 -182.755 ;
        RECT 88.235 -184.445 88.565 -184.115 ;
        RECT 88.235 -185.805 88.565 -185.475 ;
        RECT 88.235 -187.165 88.565 -186.835 ;
        RECT 88.235 -188.525 88.565 -188.195 ;
        RECT 88.235 -189.885 88.565 -189.555 ;
        RECT 88.235 -191.245 88.565 -190.915 ;
        RECT 88.235 -192.605 88.565 -192.275 ;
        RECT 88.235 -193.965 88.565 -193.635 ;
        RECT 88.235 -195.325 88.565 -194.995 ;
        RECT 88.235 -196.685 88.565 -196.355 ;
        RECT 88.235 -198.045 88.565 -197.715 ;
        RECT 88.235 -199.405 88.565 -199.075 ;
        RECT 88.235 -200.765 88.565 -200.435 ;
        RECT 88.235 -202.125 88.565 -201.795 ;
        RECT 88.235 -203.485 88.565 -203.155 ;
        RECT 88.235 -204.845 88.565 -204.515 ;
        RECT 88.235 -206.205 88.565 -205.875 ;
        RECT 88.235 -207.565 88.565 -207.235 ;
        RECT 88.235 -208.925 88.565 -208.595 ;
        RECT 88.235 -210.285 88.565 -209.955 ;
        RECT 88.235 -211.645 88.565 -211.315 ;
        RECT 88.235 -213.005 88.565 -212.675 ;
        RECT 88.235 -214.365 88.565 -214.035 ;
        RECT 88.235 -215.725 88.565 -215.395 ;
        RECT 88.235 -217.085 88.565 -216.755 ;
        RECT 88.235 -218.445 88.565 -218.115 ;
        RECT 88.235 -224.09 88.565 -222.96 ;
        RECT 88.24 -224.205 88.56 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.595 132.52 89.925 133.65 ;
        RECT 89.595 128.355 89.925 128.685 ;
        RECT 89.595 126.995 89.925 127.325 ;
        RECT 89.595 125.635 89.925 125.965 ;
        RECT 89.595 124.275 89.925 124.605 ;
        RECT 89.6 123.6 89.92 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.595 -0.845 89.925 -0.515 ;
        RECT 89.595 -2.205 89.925 -1.875 ;
        RECT 89.595 -3.565 89.925 -3.235 ;
        RECT 89.6 -3.565 89.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.955 132.52 91.285 133.65 ;
        RECT 90.955 128.355 91.285 128.685 ;
        RECT 90.955 126.995 91.285 127.325 ;
        RECT 90.955 125.635 91.285 125.965 ;
        RECT 90.955 124.275 91.285 124.605 ;
        RECT 90.96 123.6 91.28 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.955 -0.845 91.285 -0.515 ;
        RECT 90.955 -2.205 91.285 -1.875 ;
        RECT 90.955 -3.565 91.285 -3.235 ;
        RECT 90.96 -3.565 91.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.315 132.52 92.645 133.65 ;
        RECT 92.315 128.355 92.645 128.685 ;
        RECT 92.315 126.995 92.645 127.325 ;
        RECT 92.315 125.635 92.645 125.965 ;
        RECT 92.315 124.275 92.645 124.605 ;
        RECT 92.32 123.6 92.64 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.315 -0.845 92.645 -0.515 ;
        RECT 92.315 -2.205 92.645 -1.875 ;
        RECT 92.315 -3.565 92.645 -3.235 ;
        RECT 92.32 -3.565 92.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.315 -119.165 92.645 -118.835 ;
        RECT 92.315 -120.525 92.645 -120.195 ;
        RECT 92.315 -121.885 92.645 -121.555 ;
        RECT 92.315 -123.245 92.645 -122.915 ;
        RECT 92.315 -124.605 92.645 -124.275 ;
        RECT 92.315 -125.965 92.645 -125.635 ;
        RECT 92.315 -127.325 92.645 -126.995 ;
        RECT 92.315 -128.685 92.645 -128.355 ;
        RECT 92.315 -130.045 92.645 -129.715 ;
        RECT 92.315 -131.405 92.645 -131.075 ;
        RECT 92.315 -132.765 92.645 -132.435 ;
        RECT 92.315 -134.125 92.645 -133.795 ;
        RECT 92.315 -135.485 92.645 -135.155 ;
        RECT 92.315 -136.845 92.645 -136.515 ;
        RECT 92.315 -138.205 92.645 -137.875 ;
        RECT 92.315 -139.565 92.645 -139.235 ;
        RECT 92.315 -140.925 92.645 -140.595 ;
        RECT 92.315 -142.285 92.645 -141.955 ;
        RECT 92.315 -143.645 92.645 -143.315 ;
        RECT 92.315 -145.005 92.645 -144.675 ;
        RECT 92.315 -146.365 92.645 -146.035 ;
        RECT 92.315 -147.725 92.645 -147.395 ;
        RECT 92.315 -149.085 92.645 -148.755 ;
        RECT 92.315 -150.445 92.645 -150.115 ;
        RECT 92.315 -151.805 92.645 -151.475 ;
        RECT 92.315 -153.165 92.645 -152.835 ;
        RECT 92.315 -154.525 92.645 -154.195 ;
        RECT 92.315 -155.885 92.645 -155.555 ;
        RECT 92.315 -157.245 92.645 -156.915 ;
        RECT 92.315 -158.605 92.645 -158.275 ;
        RECT 92.315 -159.965 92.645 -159.635 ;
        RECT 92.315 -161.325 92.645 -160.995 ;
        RECT 92.315 -162.685 92.645 -162.355 ;
        RECT 92.315 -164.045 92.645 -163.715 ;
        RECT 92.315 -165.405 92.645 -165.075 ;
        RECT 92.315 -166.765 92.645 -166.435 ;
        RECT 92.315 -168.125 92.645 -167.795 ;
        RECT 92.315 -169.485 92.645 -169.155 ;
        RECT 92.315 -170.845 92.645 -170.515 ;
        RECT 92.315 -172.205 92.645 -171.875 ;
        RECT 92.315 -173.565 92.645 -173.235 ;
        RECT 92.315 -174.925 92.645 -174.595 ;
        RECT 92.315 -176.285 92.645 -175.955 ;
        RECT 92.315 -177.645 92.645 -177.315 ;
        RECT 92.315 -179.005 92.645 -178.675 ;
        RECT 92.315 -180.365 92.645 -180.035 ;
        RECT 92.315 -181.725 92.645 -181.395 ;
        RECT 92.315 -183.085 92.645 -182.755 ;
        RECT 92.315 -184.445 92.645 -184.115 ;
        RECT 92.315 -185.805 92.645 -185.475 ;
        RECT 92.315 -187.165 92.645 -186.835 ;
        RECT 92.315 -188.525 92.645 -188.195 ;
        RECT 92.315 -189.885 92.645 -189.555 ;
        RECT 92.315 -191.245 92.645 -190.915 ;
        RECT 92.315 -192.605 92.645 -192.275 ;
        RECT 92.315 -193.965 92.645 -193.635 ;
        RECT 92.315 -195.325 92.645 -194.995 ;
        RECT 92.315 -196.685 92.645 -196.355 ;
        RECT 92.315 -198.045 92.645 -197.715 ;
        RECT 92.315 -199.405 92.645 -199.075 ;
        RECT 92.315 -200.765 92.645 -200.435 ;
        RECT 92.315 -202.125 92.645 -201.795 ;
        RECT 92.315 -203.485 92.645 -203.155 ;
        RECT 92.315 -204.845 92.645 -204.515 ;
        RECT 92.315 -206.205 92.645 -205.875 ;
        RECT 92.315 -207.565 92.645 -207.235 ;
        RECT 92.315 -208.925 92.645 -208.595 ;
        RECT 92.315 -210.285 92.645 -209.955 ;
        RECT 92.315 -211.645 92.645 -211.315 ;
        RECT 92.315 -213.005 92.645 -212.675 ;
        RECT 92.315 -214.365 92.645 -214.035 ;
        RECT 92.315 -215.725 92.645 -215.395 ;
        RECT 92.315 -217.085 92.645 -216.755 ;
        RECT 92.315 -218.445 92.645 -218.115 ;
        RECT 92.315 -224.09 92.645 -222.96 ;
        RECT 92.32 -224.205 92.64 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.675 132.52 94.005 133.65 ;
        RECT 93.675 128.355 94.005 128.685 ;
        RECT 93.675 126.995 94.005 127.325 ;
        RECT 93.675 125.635 94.005 125.965 ;
        RECT 93.675 124.275 94.005 124.605 ;
        RECT 93.68 123.6 94 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.675 -123.245 94.005 -122.915 ;
        RECT 93.675 -124.605 94.005 -124.275 ;
        RECT 93.675 -125.965 94.005 -125.635 ;
        RECT 93.675 -127.325 94.005 -126.995 ;
        RECT 93.675 -128.685 94.005 -128.355 ;
        RECT 93.675 -130.045 94.005 -129.715 ;
        RECT 93.675 -131.405 94.005 -131.075 ;
        RECT 93.675 -132.765 94.005 -132.435 ;
        RECT 93.675 -134.125 94.005 -133.795 ;
        RECT 93.675 -135.485 94.005 -135.155 ;
        RECT 93.675 -136.845 94.005 -136.515 ;
        RECT 93.675 -138.205 94.005 -137.875 ;
        RECT 93.675 -139.565 94.005 -139.235 ;
        RECT 93.675 -140.925 94.005 -140.595 ;
        RECT 93.675 -142.285 94.005 -141.955 ;
        RECT 93.675 -143.645 94.005 -143.315 ;
        RECT 93.675 -145.005 94.005 -144.675 ;
        RECT 93.675 -146.365 94.005 -146.035 ;
        RECT 93.675 -147.725 94.005 -147.395 ;
        RECT 93.675 -149.085 94.005 -148.755 ;
        RECT 93.675 -150.445 94.005 -150.115 ;
        RECT 93.675 -151.805 94.005 -151.475 ;
        RECT 93.675 -153.165 94.005 -152.835 ;
        RECT 93.675 -154.525 94.005 -154.195 ;
        RECT 93.675 -155.885 94.005 -155.555 ;
        RECT 93.675 -157.245 94.005 -156.915 ;
        RECT 93.675 -158.605 94.005 -158.275 ;
        RECT 93.675 -159.965 94.005 -159.635 ;
        RECT 93.675 -161.325 94.005 -160.995 ;
        RECT 93.675 -162.685 94.005 -162.355 ;
        RECT 93.675 -164.045 94.005 -163.715 ;
        RECT 93.675 -165.405 94.005 -165.075 ;
        RECT 93.675 -166.765 94.005 -166.435 ;
        RECT 93.675 -168.125 94.005 -167.795 ;
        RECT 93.675 -169.485 94.005 -169.155 ;
        RECT 93.675 -170.845 94.005 -170.515 ;
        RECT 93.675 -172.205 94.005 -171.875 ;
        RECT 93.675 -173.565 94.005 -173.235 ;
        RECT 93.675 -174.925 94.005 -174.595 ;
        RECT 93.675 -176.285 94.005 -175.955 ;
        RECT 93.675 -177.645 94.005 -177.315 ;
        RECT 93.675 -179.005 94.005 -178.675 ;
        RECT 93.675 -180.365 94.005 -180.035 ;
        RECT 93.675 -181.725 94.005 -181.395 ;
        RECT 93.675 -183.085 94.005 -182.755 ;
        RECT 93.675 -184.445 94.005 -184.115 ;
        RECT 93.675 -185.805 94.005 -185.475 ;
        RECT 93.675 -187.165 94.005 -186.835 ;
        RECT 93.675 -188.525 94.005 -188.195 ;
        RECT 93.675 -189.885 94.005 -189.555 ;
        RECT 93.675 -191.245 94.005 -190.915 ;
        RECT 93.675 -192.605 94.005 -192.275 ;
        RECT 93.675 -193.965 94.005 -193.635 ;
        RECT 93.675 -195.325 94.005 -194.995 ;
        RECT 93.675 -196.685 94.005 -196.355 ;
        RECT 93.675 -198.045 94.005 -197.715 ;
        RECT 93.675 -199.405 94.005 -199.075 ;
        RECT 93.675 -200.765 94.005 -200.435 ;
        RECT 93.675 -202.125 94.005 -201.795 ;
        RECT 93.675 -203.485 94.005 -203.155 ;
        RECT 93.675 -204.845 94.005 -204.515 ;
        RECT 93.675 -206.205 94.005 -205.875 ;
        RECT 93.675 -207.565 94.005 -207.235 ;
        RECT 93.675 -208.925 94.005 -208.595 ;
        RECT 93.675 -210.285 94.005 -209.955 ;
        RECT 93.675 -211.645 94.005 -211.315 ;
        RECT 93.675 -213.005 94.005 -212.675 ;
        RECT 93.675 -214.365 94.005 -214.035 ;
        RECT 93.675 -215.725 94.005 -215.395 ;
        RECT 93.675 -217.085 94.005 -216.755 ;
        RECT 93.675 -218.445 94.005 -218.115 ;
        RECT 93.675 -224.09 94.005 -222.96 ;
        RECT 93.68 -224.205 94 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.16 -121.535 94.49 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.035 132.52 95.365 133.65 ;
        RECT 95.035 128.355 95.365 128.685 ;
        RECT 95.035 126.995 95.365 127.325 ;
        RECT 95.035 125.635 95.365 125.965 ;
        RECT 95.035 124.275 95.365 124.605 ;
        RECT 95.04 123.6 95.36 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.395 132.52 96.725 133.65 ;
        RECT 96.395 128.355 96.725 128.685 ;
        RECT 96.395 126.995 96.725 127.325 ;
        RECT 96.395 125.635 96.725 125.965 ;
        RECT 96.395 124.275 96.725 124.605 ;
        RECT 96.4 123.6 96.72 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.395 -0.845 96.725 -0.515 ;
        RECT 96.395 -2.205 96.725 -1.875 ;
        RECT 96.395 -3.565 96.725 -3.235 ;
        RECT 96.4 -3.565 96.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.395 -119.165 96.725 -118.835 ;
        RECT 96.395 -120.525 96.725 -120.195 ;
        RECT 96.395 -121.885 96.725 -121.555 ;
        RECT 96.395 -123.245 96.725 -122.915 ;
        RECT 96.395 -124.605 96.725 -124.275 ;
        RECT 96.395 -125.965 96.725 -125.635 ;
        RECT 96.395 -127.325 96.725 -126.995 ;
        RECT 96.395 -128.685 96.725 -128.355 ;
        RECT 96.395 -130.045 96.725 -129.715 ;
        RECT 96.395 -131.405 96.725 -131.075 ;
        RECT 96.395 -132.765 96.725 -132.435 ;
        RECT 96.395 -134.125 96.725 -133.795 ;
        RECT 96.395 -135.485 96.725 -135.155 ;
        RECT 96.395 -136.845 96.725 -136.515 ;
        RECT 96.395 -138.205 96.725 -137.875 ;
        RECT 96.395 -139.565 96.725 -139.235 ;
        RECT 96.395 -140.925 96.725 -140.595 ;
        RECT 96.395 -142.285 96.725 -141.955 ;
        RECT 96.395 -143.645 96.725 -143.315 ;
        RECT 96.395 -145.005 96.725 -144.675 ;
        RECT 96.395 -146.365 96.725 -146.035 ;
        RECT 96.395 -147.725 96.725 -147.395 ;
        RECT 96.395 -149.085 96.725 -148.755 ;
        RECT 96.395 -150.445 96.725 -150.115 ;
        RECT 96.395 -151.805 96.725 -151.475 ;
        RECT 96.395 -153.165 96.725 -152.835 ;
        RECT 96.395 -154.525 96.725 -154.195 ;
        RECT 96.395 -155.885 96.725 -155.555 ;
        RECT 96.395 -157.245 96.725 -156.915 ;
        RECT 96.395 -158.605 96.725 -158.275 ;
        RECT 96.395 -159.965 96.725 -159.635 ;
        RECT 96.395 -161.325 96.725 -160.995 ;
        RECT 96.395 -162.685 96.725 -162.355 ;
        RECT 96.395 -164.045 96.725 -163.715 ;
        RECT 96.395 -165.405 96.725 -165.075 ;
        RECT 96.395 -166.765 96.725 -166.435 ;
        RECT 96.395 -168.125 96.725 -167.795 ;
        RECT 96.395 -169.485 96.725 -169.155 ;
        RECT 96.395 -170.845 96.725 -170.515 ;
        RECT 96.395 -172.205 96.725 -171.875 ;
        RECT 96.395 -173.565 96.725 -173.235 ;
        RECT 96.395 -174.925 96.725 -174.595 ;
        RECT 96.395 -176.285 96.725 -175.955 ;
        RECT 96.395 -177.645 96.725 -177.315 ;
        RECT 96.395 -179.005 96.725 -178.675 ;
        RECT 96.395 -180.365 96.725 -180.035 ;
        RECT 96.395 -181.725 96.725 -181.395 ;
        RECT 96.395 -183.085 96.725 -182.755 ;
        RECT 96.395 -184.445 96.725 -184.115 ;
        RECT 96.395 -185.805 96.725 -185.475 ;
        RECT 96.395 -187.165 96.725 -186.835 ;
        RECT 96.395 -188.525 96.725 -188.195 ;
        RECT 96.395 -189.885 96.725 -189.555 ;
        RECT 96.395 -191.245 96.725 -190.915 ;
        RECT 96.395 -192.605 96.725 -192.275 ;
        RECT 96.395 -193.965 96.725 -193.635 ;
        RECT 96.395 -195.325 96.725 -194.995 ;
        RECT 96.395 -196.685 96.725 -196.355 ;
        RECT 96.395 -198.045 96.725 -197.715 ;
        RECT 96.395 -199.405 96.725 -199.075 ;
        RECT 96.395 -200.765 96.725 -200.435 ;
        RECT 96.395 -202.125 96.725 -201.795 ;
        RECT 96.395 -203.485 96.725 -203.155 ;
        RECT 96.395 -204.845 96.725 -204.515 ;
        RECT 96.395 -206.205 96.725 -205.875 ;
        RECT 96.395 -207.565 96.725 -207.235 ;
        RECT 96.395 -208.925 96.725 -208.595 ;
        RECT 96.395 -210.285 96.725 -209.955 ;
        RECT 96.395 -211.645 96.725 -211.315 ;
        RECT 96.395 -213.005 96.725 -212.675 ;
        RECT 96.395 -214.365 96.725 -214.035 ;
        RECT 96.395 -215.725 96.725 -215.395 ;
        RECT 96.395 -217.085 96.725 -216.755 ;
        RECT 96.395 -218.445 96.725 -218.115 ;
        RECT 96.395 -224.09 96.725 -222.96 ;
        RECT 96.4 -224.205 96.72 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.755 132.52 98.085 133.65 ;
        RECT 97.755 128.355 98.085 128.685 ;
        RECT 97.755 126.995 98.085 127.325 ;
        RECT 97.755 125.635 98.085 125.965 ;
        RECT 97.755 124.275 98.085 124.605 ;
        RECT 97.76 123.6 98.08 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.755 -0.845 98.085 -0.515 ;
        RECT 97.755 -2.205 98.085 -1.875 ;
        RECT 97.755 -3.565 98.085 -3.235 ;
        RECT 97.76 -3.565 98.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.115 132.52 99.445 133.65 ;
        RECT 99.115 128.355 99.445 128.685 ;
        RECT 99.115 126.995 99.445 127.325 ;
        RECT 99.115 125.635 99.445 125.965 ;
        RECT 99.115 124.275 99.445 124.605 ;
        RECT 99.12 123.6 99.44 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.115 -0.845 99.445 -0.515 ;
        RECT 99.115 -2.205 99.445 -1.875 ;
        RECT 99.115 -3.565 99.445 -3.235 ;
        RECT 99.12 -3.565 99.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.115 -119.165 99.445 -118.835 ;
        RECT 99.115 -120.525 99.445 -120.195 ;
        RECT 99.115 -121.885 99.445 -121.555 ;
        RECT 99.115 -123.245 99.445 -122.915 ;
        RECT 99.115 -124.605 99.445 -124.275 ;
        RECT 99.115 -125.965 99.445 -125.635 ;
        RECT 99.115 -127.325 99.445 -126.995 ;
        RECT 99.115 -128.685 99.445 -128.355 ;
        RECT 99.115 -130.045 99.445 -129.715 ;
        RECT 99.115 -131.405 99.445 -131.075 ;
        RECT 99.115 -132.765 99.445 -132.435 ;
        RECT 99.115 -134.125 99.445 -133.795 ;
        RECT 99.115 -135.485 99.445 -135.155 ;
        RECT 99.115 -136.845 99.445 -136.515 ;
        RECT 99.115 -138.205 99.445 -137.875 ;
        RECT 99.115 -139.565 99.445 -139.235 ;
        RECT 99.115 -140.925 99.445 -140.595 ;
        RECT 99.115 -142.285 99.445 -141.955 ;
        RECT 99.115 -143.645 99.445 -143.315 ;
        RECT 99.115 -145.005 99.445 -144.675 ;
        RECT 99.115 -146.365 99.445 -146.035 ;
        RECT 99.115 -147.725 99.445 -147.395 ;
        RECT 99.115 -149.085 99.445 -148.755 ;
        RECT 99.115 -150.445 99.445 -150.115 ;
        RECT 99.115 -151.805 99.445 -151.475 ;
        RECT 99.115 -153.165 99.445 -152.835 ;
        RECT 99.115 -154.525 99.445 -154.195 ;
        RECT 99.115 -155.885 99.445 -155.555 ;
        RECT 99.115 -157.245 99.445 -156.915 ;
        RECT 99.115 -158.605 99.445 -158.275 ;
        RECT 99.115 -159.965 99.445 -159.635 ;
        RECT 99.115 -161.325 99.445 -160.995 ;
        RECT 99.115 -162.685 99.445 -162.355 ;
        RECT 99.115 -164.045 99.445 -163.715 ;
        RECT 99.115 -165.405 99.445 -165.075 ;
        RECT 99.115 -166.765 99.445 -166.435 ;
        RECT 99.115 -168.125 99.445 -167.795 ;
        RECT 99.115 -169.485 99.445 -169.155 ;
        RECT 99.115 -170.845 99.445 -170.515 ;
        RECT 99.115 -172.205 99.445 -171.875 ;
        RECT 99.115 -173.565 99.445 -173.235 ;
        RECT 99.115 -174.925 99.445 -174.595 ;
        RECT 99.115 -176.285 99.445 -175.955 ;
        RECT 99.115 -177.645 99.445 -177.315 ;
        RECT 99.115 -179.005 99.445 -178.675 ;
        RECT 99.115 -180.365 99.445 -180.035 ;
        RECT 99.115 -181.725 99.445 -181.395 ;
        RECT 99.115 -183.085 99.445 -182.755 ;
        RECT 99.115 -184.445 99.445 -184.115 ;
        RECT 99.115 -185.805 99.445 -185.475 ;
        RECT 99.115 -187.165 99.445 -186.835 ;
        RECT 99.115 -188.525 99.445 -188.195 ;
        RECT 99.115 -189.885 99.445 -189.555 ;
        RECT 99.115 -191.245 99.445 -190.915 ;
        RECT 99.115 -192.605 99.445 -192.275 ;
        RECT 99.115 -193.965 99.445 -193.635 ;
        RECT 99.115 -195.325 99.445 -194.995 ;
        RECT 99.115 -196.685 99.445 -196.355 ;
        RECT 99.115 -198.045 99.445 -197.715 ;
        RECT 99.115 -199.405 99.445 -199.075 ;
        RECT 99.115 -200.765 99.445 -200.435 ;
        RECT 99.115 -202.125 99.445 -201.795 ;
        RECT 99.115 -203.485 99.445 -203.155 ;
        RECT 99.115 -204.845 99.445 -204.515 ;
        RECT 99.115 -206.205 99.445 -205.875 ;
        RECT 99.115 -207.565 99.445 -207.235 ;
        RECT 99.115 -208.925 99.445 -208.595 ;
        RECT 99.115 -210.285 99.445 -209.955 ;
        RECT 99.115 -211.645 99.445 -211.315 ;
        RECT 99.115 -213.005 99.445 -212.675 ;
        RECT 99.115 -214.365 99.445 -214.035 ;
        RECT 99.115 -215.725 99.445 -215.395 ;
        RECT 99.115 -217.085 99.445 -216.755 ;
        RECT 99.115 -218.445 99.445 -218.115 ;
        RECT 99.115 -224.09 99.445 -222.96 ;
        RECT 99.12 -224.205 99.44 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.26 -121.535 100.59 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.475 132.52 100.805 133.65 ;
        RECT 100.475 128.355 100.805 128.685 ;
        RECT 100.475 126.995 100.805 127.325 ;
        RECT 100.475 125.635 100.805 125.965 ;
        RECT 100.475 124.275 100.805 124.605 ;
        RECT 100.48 123.6 100.8 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.475 -125.965 100.805 -125.635 ;
        RECT 100.475 -127.325 100.805 -126.995 ;
        RECT 100.475 -128.685 100.805 -128.355 ;
        RECT 100.475 -130.045 100.805 -129.715 ;
        RECT 100.475 -131.405 100.805 -131.075 ;
        RECT 100.475 -132.765 100.805 -132.435 ;
        RECT 100.475 -134.125 100.805 -133.795 ;
        RECT 100.475 -135.485 100.805 -135.155 ;
        RECT 100.475 -136.845 100.805 -136.515 ;
        RECT 100.475 -138.205 100.805 -137.875 ;
        RECT 100.475 -139.565 100.805 -139.235 ;
        RECT 100.475 -140.925 100.805 -140.595 ;
        RECT 100.475 -142.285 100.805 -141.955 ;
        RECT 100.475 -143.645 100.805 -143.315 ;
        RECT 100.475 -145.005 100.805 -144.675 ;
        RECT 100.475 -146.365 100.805 -146.035 ;
        RECT 100.475 -147.725 100.805 -147.395 ;
        RECT 100.475 -149.085 100.805 -148.755 ;
        RECT 100.475 -150.445 100.805 -150.115 ;
        RECT 100.475 -151.805 100.805 -151.475 ;
        RECT 100.475 -153.165 100.805 -152.835 ;
        RECT 100.475 -154.525 100.805 -154.195 ;
        RECT 100.475 -155.885 100.805 -155.555 ;
        RECT 100.475 -157.245 100.805 -156.915 ;
        RECT 100.475 -158.605 100.805 -158.275 ;
        RECT 100.475 -159.965 100.805 -159.635 ;
        RECT 100.475 -161.325 100.805 -160.995 ;
        RECT 100.475 -162.685 100.805 -162.355 ;
        RECT 100.475 -164.045 100.805 -163.715 ;
        RECT 100.475 -165.405 100.805 -165.075 ;
        RECT 100.475 -166.765 100.805 -166.435 ;
        RECT 100.475 -168.125 100.805 -167.795 ;
        RECT 100.475 -169.485 100.805 -169.155 ;
        RECT 100.475 -170.845 100.805 -170.515 ;
        RECT 100.475 -172.205 100.805 -171.875 ;
        RECT 100.475 -173.565 100.805 -173.235 ;
        RECT 100.475 -174.925 100.805 -174.595 ;
        RECT 100.475 -176.285 100.805 -175.955 ;
        RECT 100.475 -177.645 100.805 -177.315 ;
        RECT 100.475 -179.005 100.805 -178.675 ;
        RECT 100.475 -180.365 100.805 -180.035 ;
        RECT 100.475 -181.725 100.805 -181.395 ;
        RECT 100.475 -183.085 100.805 -182.755 ;
        RECT 100.475 -184.445 100.805 -184.115 ;
        RECT 100.475 -185.805 100.805 -185.475 ;
        RECT 100.475 -187.165 100.805 -186.835 ;
        RECT 100.475 -188.525 100.805 -188.195 ;
        RECT 100.475 -189.885 100.805 -189.555 ;
        RECT 100.475 -191.245 100.805 -190.915 ;
        RECT 100.475 -192.605 100.805 -192.275 ;
        RECT 100.475 -193.965 100.805 -193.635 ;
        RECT 100.475 -195.325 100.805 -194.995 ;
        RECT 100.475 -196.685 100.805 -196.355 ;
        RECT 100.475 -198.045 100.805 -197.715 ;
        RECT 100.475 -199.405 100.805 -199.075 ;
        RECT 100.475 -200.765 100.805 -200.435 ;
        RECT 100.475 -202.125 100.805 -201.795 ;
        RECT 100.475 -203.485 100.805 -203.155 ;
        RECT 100.475 -204.845 100.805 -204.515 ;
        RECT 100.475 -206.205 100.805 -205.875 ;
        RECT 100.475 -207.565 100.805 -207.235 ;
        RECT 100.475 -208.925 100.805 -208.595 ;
        RECT 100.475 -210.285 100.805 -209.955 ;
        RECT 100.475 -211.645 100.805 -211.315 ;
        RECT 100.475 -213.005 100.805 -212.675 ;
        RECT 100.475 -214.365 100.805 -214.035 ;
        RECT 100.475 -215.725 100.805 -215.395 ;
        RECT 100.475 -217.085 100.805 -216.755 ;
        RECT 100.475 -218.445 100.805 -218.115 ;
        RECT 100.475 -224.09 100.805 -222.96 ;
        RECT 100.48 -224.205 100.8 -122.24 ;
        RECT 100.475 -123.245 100.805 -122.915 ;
        RECT 100.475 -124.605 100.805 -124.275 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.36 -121.535 45.69 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.075 132.52 46.405 133.65 ;
        RECT 46.075 128.355 46.405 128.685 ;
        RECT 46.075 126.995 46.405 127.325 ;
        RECT 46.075 125.635 46.405 125.965 ;
        RECT 46.075 124.275 46.405 124.605 ;
        RECT 46.08 123.6 46.4 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.435 132.52 47.765 133.65 ;
        RECT 47.435 128.355 47.765 128.685 ;
        RECT 47.435 126.995 47.765 127.325 ;
        RECT 47.435 125.635 47.765 125.965 ;
        RECT 47.435 124.275 47.765 124.605 ;
        RECT 47.44 123.6 47.76 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.435 -0.845 47.765 -0.515 ;
        RECT 47.435 -2.205 47.765 -1.875 ;
        RECT 47.435 -3.565 47.765 -3.235 ;
        RECT 47.44 -3.565 47.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.795 132.52 49.125 133.65 ;
        RECT 48.795 128.355 49.125 128.685 ;
        RECT 48.795 126.995 49.125 127.325 ;
        RECT 48.795 125.635 49.125 125.965 ;
        RECT 48.795 124.275 49.125 124.605 ;
        RECT 48.8 123.6 49.12 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.795 -0.845 49.125 -0.515 ;
        RECT 48.795 -2.205 49.125 -1.875 ;
        RECT 48.795 -3.565 49.125 -3.235 ;
        RECT 48.8 -3.565 49.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.155 132.52 50.485 133.65 ;
        RECT 50.155 128.355 50.485 128.685 ;
        RECT 50.155 126.995 50.485 127.325 ;
        RECT 50.155 125.635 50.485 125.965 ;
        RECT 50.155 124.275 50.485 124.605 ;
        RECT 50.16 123.6 50.48 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.155 -0.845 50.485 -0.515 ;
        RECT 50.155 -2.205 50.485 -1.875 ;
        RECT 50.155 -3.565 50.485 -3.235 ;
        RECT 50.16 -3.565 50.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.155 -119.165 50.485 -118.835 ;
        RECT 50.155 -120.525 50.485 -120.195 ;
        RECT 50.155 -121.885 50.485 -121.555 ;
        RECT 50.155 -123.245 50.485 -122.915 ;
        RECT 50.155 -124.605 50.485 -124.275 ;
        RECT 50.155 -125.965 50.485 -125.635 ;
        RECT 50.155 -127.325 50.485 -126.995 ;
        RECT 50.155 -128.685 50.485 -128.355 ;
        RECT 50.155 -130.045 50.485 -129.715 ;
        RECT 50.155 -131.405 50.485 -131.075 ;
        RECT 50.155 -132.765 50.485 -132.435 ;
        RECT 50.155 -134.125 50.485 -133.795 ;
        RECT 50.155 -135.485 50.485 -135.155 ;
        RECT 50.155 -136.845 50.485 -136.515 ;
        RECT 50.155 -138.205 50.485 -137.875 ;
        RECT 50.155 -139.565 50.485 -139.235 ;
        RECT 50.155 -140.925 50.485 -140.595 ;
        RECT 50.155 -142.285 50.485 -141.955 ;
        RECT 50.155 -143.645 50.485 -143.315 ;
        RECT 50.155 -145.005 50.485 -144.675 ;
        RECT 50.155 -146.365 50.485 -146.035 ;
        RECT 50.155 -147.725 50.485 -147.395 ;
        RECT 50.155 -149.085 50.485 -148.755 ;
        RECT 50.155 -150.445 50.485 -150.115 ;
        RECT 50.155 -151.805 50.485 -151.475 ;
        RECT 50.155 -153.165 50.485 -152.835 ;
        RECT 50.155 -154.525 50.485 -154.195 ;
        RECT 50.155 -155.885 50.485 -155.555 ;
        RECT 50.155 -157.245 50.485 -156.915 ;
        RECT 50.155 -158.605 50.485 -158.275 ;
        RECT 50.155 -159.965 50.485 -159.635 ;
        RECT 50.155 -161.325 50.485 -160.995 ;
        RECT 50.155 -162.685 50.485 -162.355 ;
        RECT 50.155 -164.045 50.485 -163.715 ;
        RECT 50.155 -165.405 50.485 -165.075 ;
        RECT 50.155 -166.765 50.485 -166.435 ;
        RECT 50.155 -168.125 50.485 -167.795 ;
        RECT 50.155 -169.485 50.485 -169.155 ;
        RECT 50.155 -170.845 50.485 -170.515 ;
        RECT 50.155 -172.205 50.485 -171.875 ;
        RECT 50.155 -173.565 50.485 -173.235 ;
        RECT 50.155 -174.925 50.485 -174.595 ;
        RECT 50.155 -176.285 50.485 -175.955 ;
        RECT 50.155 -177.645 50.485 -177.315 ;
        RECT 50.155 -179.005 50.485 -178.675 ;
        RECT 50.155 -180.365 50.485 -180.035 ;
        RECT 50.155 -181.725 50.485 -181.395 ;
        RECT 50.155 -183.085 50.485 -182.755 ;
        RECT 50.155 -184.445 50.485 -184.115 ;
        RECT 50.155 -185.805 50.485 -185.475 ;
        RECT 50.155 -187.165 50.485 -186.835 ;
        RECT 50.155 -188.525 50.485 -188.195 ;
        RECT 50.155 -189.885 50.485 -189.555 ;
        RECT 50.155 -191.245 50.485 -190.915 ;
        RECT 50.155 -192.605 50.485 -192.275 ;
        RECT 50.155 -193.965 50.485 -193.635 ;
        RECT 50.155 -195.325 50.485 -194.995 ;
        RECT 50.155 -196.685 50.485 -196.355 ;
        RECT 50.155 -198.045 50.485 -197.715 ;
        RECT 50.155 -199.405 50.485 -199.075 ;
        RECT 50.155 -200.765 50.485 -200.435 ;
        RECT 50.155 -202.125 50.485 -201.795 ;
        RECT 50.155 -203.485 50.485 -203.155 ;
        RECT 50.155 -204.845 50.485 -204.515 ;
        RECT 50.155 -206.205 50.485 -205.875 ;
        RECT 50.155 -207.565 50.485 -207.235 ;
        RECT 50.155 -208.925 50.485 -208.595 ;
        RECT 50.155 -210.285 50.485 -209.955 ;
        RECT 50.155 -211.645 50.485 -211.315 ;
        RECT 50.155 -213.005 50.485 -212.675 ;
        RECT 50.155 -214.365 50.485 -214.035 ;
        RECT 50.155 -215.725 50.485 -215.395 ;
        RECT 50.155 -217.085 50.485 -216.755 ;
        RECT 50.155 -218.445 50.485 -218.115 ;
        RECT 50.155 -224.09 50.485 -222.96 ;
        RECT 50.16 -224.205 50.48 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.46 -121.535 51.79 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.515 132.52 51.845 133.65 ;
        RECT 51.515 128.355 51.845 128.685 ;
        RECT 51.515 126.995 51.845 127.325 ;
        RECT 51.515 125.635 51.845 125.965 ;
        RECT 51.515 124.275 51.845 124.605 ;
        RECT 51.52 123.6 51.84 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.515 -123.245 51.845 -122.915 ;
        RECT 51.515 -124.605 51.845 -124.275 ;
        RECT 51.515 -125.965 51.845 -125.635 ;
        RECT 51.515 -127.325 51.845 -126.995 ;
        RECT 51.515 -128.685 51.845 -128.355 ;
        RECT 51.515 -130.045 51.845 -129.715 ;
        RECT 51.515 -131.405 51.845 -131.075 ;
        RECT 51.515 -132.765 51.845 -132.435 ;
        RECT 51.515 -134.125 51.845 -133.795 ;
        RECT 51.515 -135.485 51.845 -135.155 ;
        RECT 51.515 -136.845 51.845 -136.515 ;
        RECT 51.515 -138.205 51.845 -137.875 ;
        RECT 51.515 -139.565 51.845 -139.235 ;
        RECT 51.515 -140.925 51.845 -140.595 ;
        RECT 51.515 -142.285 51.845 -141.955 ;
        RECT 51.515 -143.645 51.845 -143.315 ;
        RECT 51.515 -145.005 51.845 -144.675 ;
        RECT 51.515 -146.365 51.845 -146.035 ;
        RECT 51.515 -147.725 51.845 -147.395 ;
        RECT 51.515 -149.085 51.845 -148.755 ;
        RECT 51.515 -150.445 51.845 -150.115 ;
        RECT 51.515 -151.805 51.845 -151.475 ;
        RECT 51.515 -153.165 51.845 -152.835 ;
        RECT 51.515 -154.525 51.845 -154.195 ;
        RECT 51.515 -155.885 51.845 -155.555 ;
        RECT 51.515 -157.245 51.845 -156.915 ;
        RECT 51.515 -158.605 51.845 -158.275 ;
        RECT 51.515 -159.965 51.845 -159.635 ;
        RECT 51.515 -161.325 51.845 -160.995 ;
        RECT 51.515 -162.685 51.845 -162.355 ;
        RECT 51.515 -164.045 51.845 -163.715 ;
        RECT 51.515 -165.405 51.845 -165.075 ;
        RECT 51.515 -166.765 51.845 -166.435 ;
        RECT 51.515 -168.125 51.845 -167.795 ;
        RECT 51.515 -169.485 51.845 -169.155 ;
        RECT 51.515 -170.845 51.845 -170.515 ;
        RECT 51.515 -172.205 51.845 -171.875 ;
        RECT 51.515 -173.565 51.845 -173.235 ;
        RECT 51.515 -174.925 51.845 -174.595 ;
        RECT 51.515 -176.285 51.845 -175.955 ;
        RECT 51.515 -177.645 51.845 -177.315 ;
        RECT 51.515 -179.005 51.845 -178.675 ;
        RECT 51.515 -180.365 51.845 -180.035 ;
        RECT 51.515 -181.725 51.845 -181.395 ;
        RECT 51.515 -183.085 51.845 -182.755 ;
        RECT 51.515 -184.445 51.845 -184.115 ;
        RECT 51.515 -185.805 51.845 -185.475 ;
        RECT 51.515 -187.165 51.845 -186.835 ;
        RECT 51.515 -188.525 51.845 -188.195 ;
        RECT 51.515 -189.885 51.845 -189.555 ;
        RECT 51.515 -191.245 51.845 -190.915 ;
        RECT 51.515 -192.605 51.845 -192.275 ;
        RECT 51.515 -193.965 51.845 -193.635 ;
        RECT 51.515 -195.325 51.845 -194.995 ;
        RECT 51.515 -196.685 51.845 -196.355 ;
        RECT 51.515 -198.045 51.845 -197.715 ;
        RECT 51.515 -199.405 51.845 -199.075 ;
        RECT 51.515 -200.765 51.845 -200.435 ;
        RECT 51.515 -202.125 51.845 -201.795 ;
        RECT 51.515 -203.485 51.845 -203.155 ;
        RECT 51.515 -204.845 51.845 -204.515 ;
        RECT 51.515 -206.205 51.845 -205.875 ;
        RECT 51.515 -207.565 51.845 -207.235 ;
        RECT 51.515 -208.925 51.845 -208.595 ;
        RECT 51.515 -210.285 51.845 -209.955 ;
        RECT 51.515 -211.645 51.845 -211.315 ;
        RECT 51.515 -213.005 51.845 -212.675 ;
        RECT 51.515 -214.365 51.845 -214.035 ;
        RECT 51.515 -215.725 51.845 -215.395 ;
        RECT 51.515 -217.085 51.845 -216.755 ;
        RECT 51.515 -218.445 51.845 -218.115 ;
        RECT 51.515 -224.09 51.845 -222.96 ;
        RECT 51.52 -224.205 51.84 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.875 132.52 53.205 133.65 ;
        RECT 52.875 128.355 53.205 128.685 ;
        RECT 52.875 126.995 53.205 127.325 ;
        RECT 52.875 125.635 53.205 125.965 ;
        RECT 52.875 124.275 53.205 124.605 ;
        RECT 52.88 123.6 53.2 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.875 -0.845 53.205 -0.515 ;
        RECT 52.875 -2.205 53.205 -1.875 ;
        RECT 52.875 -3.565 53.205 -3.235 ;
        RECT 52.88 -3.565 53.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.235 132.52 54.565 133.65 ;
        RECT 54.235 128.355 54.565 128.685 ;
        RECT 54.235 126.995 54.565 127.325 ;
        RECT 54.235 125.635 54.565 125.965 ;
        RECT 54.235 124.275 54.565 124.605 ;
        RECT 54.24 123.6 54.56 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.235 -0.845 54.565 -0.515 ;
        RECT 54.235 -2.205 54.565 -1.875 ;
        RECT 54.235 -3.565 54.565 -3.235 ;
        RECT 54.24 -3.565 54.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.595 132.52 55.925 133.65 ;
        RECT 55.595 128.355 55.925 128.685 ;
        RECT 55.595 126.995 55.925 127.325 ;
        RECT 55.595 125.635 55.925 125.965 ;
        RECT 55.595 124.275 55.925 124.605 ;
        RECT 55.6 123.6 55.92 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.595 -0.845 55.925 -0.515 ;
        RECT 55.595 -2.205 55.925 -1.875 ;
        RECT 55.595 -3.565 55.925 -3.235 ;
        RECT 55.6 -3.565 55.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.955 132.52 57.285 133.65 ;
        RECT 56.955 128.355 57.285 128.685 ;
        RECT 56.955 126.995 57.285 127.325 ;
        RECT 56.955 125.635 57.285 125.965 ;
        RECT 56.955 124.275 57.285 124.605 ;
        RECT 56.96 123.6 57.28 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.955 -123.245 57.285 -122.915 ;
        RECT 56.955 -124.605 57.285 -124.275 ;
        RECT 56.955 -125.965 57.285 -125.635 ;
        RECT 56.955 -127.325 57.285 -126.995 ;
        RECT 56.955 -128.685 57.285 -128.355 ;
        RECT 56.955 -130.045 57.285 -129.715 ;
        RECT 56.955 -131.405 57.285 -131.075 ;
        RECT 56.955 -132.765 57.285 -132.435 ;
        RECT 56.955 -134.125 57.285 -133.795 ;
        RECT 56.955 -135.485 57.285 -135.155 ;
        RECT 56.955 -136.845 57.285 -136.515 ;
        RECT 56.955 -138.205 57.285 -137.875 ;
        RECT 56.955 -139.565 57.285 -139.235 ;
        RECT 56.955 -140.925 57.285 -140.595 ;
        RECT 56.955 -142.285 57.285 -141.955 ;
        RECT 56.955 -143.645 57.285 -143.315 ;
        RECT 56.955 -145.005 57.285 -144.675 ;
        RECT 56.955 -146.365 57.285 -146.035 ;
        RECT 56.955 -147.725 57.285 -147.395 ;
        RECT 56.955 -149.085 57.285 -148.755 ;
        RECT 56.955 -150.445 57.285 -150.115 ;
        RECT 56.955 -151.805 57.285 -151.475 ;
        RECT 56.955 -153.165 57.285 -152.835 ;
        RECT 56.955 -154.525 57.285 -154.195 ;
        RECT 56.955 -155.885 57.285 -155.555 ;
        RECT 56.955 -157.245 57.285 -156.915 ;
        RECT 56.955 -158.605 57.285 -158.275 ;
        RECT 56.955 -159.965 57.285 -159.635 ;
        RECT 56.955 -161.325 57.285 -160.995 ;
        RECT 56.955 -162.685 57.285 -162.355 ;
        RECT 56.955 -164.045 57.285 -163.715 ;
        RECT 56.955 -165.405 57.285 -165.075 ;
        RECT 56.955 -166.765 57.285 -166.435 ;
        RECT 56.955 -168.125 57.285 -167.795 ;
        RECT 56.955 -169.485 57.285 -169.155 ;
        RECT 56.955 -170.845 57.285 -170.515 ;
        RECT 56.955 -172.205 57.285 -171.875 ;
        RECT 56.955 -173.565 57.285 -173.235 ;
        RECT 56.955 -174.925 57.285 -174.595 ;
        RECT 56.955 -176.285 57.285 -175.955 ;
        RECT 56.955 -177.645 57.285 -177.315 ;
        RECT 56.955 -179.005 57.285 -178.675 ;
        RECT 56.955 -180.365 57.285 -180.035 ;
        RECT 56.955 -181.725 57.285 -181.395 ;
        RECT 56.955 -183.085 57.285 -182.755 ;
        RECT 56.955 -184.445 57.285 -184.115 ;
        RECT 56.955 -185.805 57.285 -185.475 ;
        RECT 56.955 -187.165 57.285 -186.835 ;
        RECT 56.955 -188.525 57.285 -188.195 ;
        RECT 56.955 -189.885 57.285 -189.555 ;
        RECT 56.955 -191.245 57.285 -190.915 ;
        RECT 56.955 -192.605 57.285 -192.275 ;
        RECT 56.955 -193.965 57.285 -193.635 ;
        RECT 56.955 -195.325 57.285 -194.995 ;
        RECT 56.955 -196.685 57.285 -196.355 ;
        RECT 56.955 -198.045 57.285 -197.715 ;
        RECT 56.955 -199.405 57.285 -199.075 ;
        RECT 56.955 -200.765 57.285 -200.435 ;
        RECT 56.955 -202.125 57.285 -201.795 ;
        RECT 56.955 -203.485 57.285 -203.155 ;
        RECT 56.955 -204.845 57.285 -204.515 ;
        RECT 56.955 -206.205 57.285 -205.875 ;
        RECT 56.955 -207.565 57.285 -207.235 ;
        RECT 56.955 -208.925 57.285 -208.595 ;
        RECT 56.955 -210.285 57.285 -209.955 ;
        RECT 56.955 -211.645 57.285 -211.315 ;
        RECT 56.955 -213.005 57.285 -212.675 ;
        RECT 56.955 -214.365 57.285 -214.035 ;
        RECT 56.955 -215.725 57.285 -215.395 ;
        RECT 56.955 -217.085 57.285 -216.755 ;
        RECT 56.955 -218.445 57.285 -218.115 ;
        RECT 56.955 -224.09 57.285 -222.96 ;
        RECT 56.96 -224.205 57.28 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.56 -121.535 57.89 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.315 132.52 58.645 133.65 ;
        RECT 58.315 128.355 58.645 128.685 ;
        RECT 58.315 126.995 58.645 127.325 ;
        RECT 58.315 125.635 58.645 125.965 ;
        RECT 58.315 124.275 58.645 124.605 ;
        RECT 58.32 123.6 58.64 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.675 132.52 60.005 133.65 ;
        RECT 59.675 128.355 60.005 128.685 ;
        RECT 59.675 126.995 60.005 127.325 ;
        RECT 59.675 125.635 60.005 125.965 ;
        RECT 59.675 124.275 60.005 124.605 ;
        RECT 59.68 123.6 60 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.675 -0.845 60.005 -0.515 ;
        RECT 59.675 -2.205 60.005 -1.875 ;
        RECT 59.675 -3.565 60.005 -3.235 ;
        RECT 59.68 -3.565 60 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.675 -119.165 60.005 -118.835 ;
        RECT 59.675 -120.525 60.005 -120.195 ;
        RECT 59.675 -121.885 60.005 -121.555 ;
        RECT 59.675 -123.245 60.005 -122.915 ;
        RECT 59.675 -124.605 60.005 -124.275 ;
        RECT 59.675 -125.965 60.005 -125.635 ;
        RECT 59.675 -127.325 60.005 -126.995 ;
        RECT 59.675 -128.685 60.005 -128.355 ;
        RECT 59.675 -130.045 60.005 -129.715 ;
        RECT 59.675 -131.405 60.005 -131.075 ;
        RECT 59.675 -132.765 60.005 -132.435 ;
        RECT 59.675 -134.125 60.005 -133.795 ;
        RECT 59.675 -135.485 60.005 -135.155 ;
        RECT 59.675 -136.845 60.005 -136.515 ;
        RECT 59.675 -138.205 60.005 -137.875 ;
        RECT 59.675 -139.565 60.005 -139.235 ;
        RECT 59.675 -140.925 60.005 -140.595 ;
        RECT 59.675 -142.285 60.005 -141.955 ;
        RECT 59.675 -143.645 60.005 -143.315 ;
        RECT 59.675 -145.005 60.005 -144.675 ;
        RECT 59.675 -146.365 60.005 -146.035 ;
        RECT 59.675 -147.725 60.005 -147.395 ;
        RECT 59.675 -149.085 60.005 -148.755 ;
        RECT 59.675 -150.445 60.005 -150.115 ;
        RECT 59.675 -151.805 60.005 -151.475 ;
        RECT 59.675 -153.165 60.005 -152.835 ;
        RECT 59.675 -154.525 60.005 -154.195 ;
        RECT 59.675 -155.885 60.005 -155.555 ;
        RECT 59.675 -157.245 60.005 -156.915 ;
        RECT 59.675 -158.605 60.005 -158.275 ;
        RECT 59.675 -159.965 60.005 -159.635 ;
        RECT 59.675 -161.325 60.005 -160.995 ;
        RECT 59.675 -162.685 60.005 -162.355 ;
        RECT 59.675 -164.045 60.005 -163.715 ;
        RECT 59.675 -165.405 60.005 -165.075 ;
        RECT 59.675 -166.765 60.005 -166.435 ;
        RECT 59.675 -168.125 60.005 -167.795 ;
        RECT 59.675 -169.485 60.005 -169.155 ;
        RECT 59.675 -170.845 60.005 -170.515 ;
        RECT 59.675 -172.205 60.005 -171.875 ;
        RECT 59.675 -173.565 60.005 -173.235 ;
        RECT 59.675 -174.925 60.005 -174.595 ;
        RECT 59.675 -176.285 60.005 -175.955 ;
        RECT 59.675 -177.645 60.005 -177.315 ;
        RECT 59.675 -179.005 60.005 -178.675 ;
        RECT 59.675 -180.365 60.005 -180.035 ;
        RECT 59.675 -181.725 60.005 -181.395 ;
        RECT 59.675 -183.085 60.005 -182.755 ;
        RECT 59.675 -184.445 60.005 -184.115 ;
        RECT 59.675 -185.805 60.005 -185.475 ;
        RECT 59.675 -187.165 60.005 -186.835 ;
        RECT 59.675 -188.525 60.005 -188.195 ;
        RECT 59.675 -189.885 60.005 -189.555 ;
        RECT 59.675 -191.245 60.005 -190.915 ;
        RECT 59.675 -192.605 60.005 -192.275 ;
        RECT 59.675 -193.965 60.005 -193.635 ;
        RECT 59.675 -195.325 60.005 -194.995 ;
        RECT 59.675 -196.685 60.005 -196.355 ;
        RECT 59.675 -198.045 60.005 -197.715 ;
        RECT 59.675 -199.405 60.005 -199.075 ;
        RECT 59.675 -200.765 60.005 -200.435 ;
        RECT 59.675 -202.125 60.005 -201.795 ;
        RECT 59.675 -203.485 60.005 -203.155 ;
        RECT 59.675 -204.845 60.005 -204.515 ;
        RECT 59.675 -206.205 60.005 -205.875 ;
        RECT 59.675 -207.565 60.005 -207.235 ;
        RECT 59.675 -208.925 60.005 -208.595 ;
        RECT 59.675 -210.285 60.005 -209.955 ;
        RECT 59.675 -211.645 60.005 -211.315 ;
        RECT 59.675 -213.005 60.005 -212.675 ;
        RECT 59.675 -214.365 60.005 -214.035 ;
        RECT 59.675 -215.725 60.005 -215.395 ;
        RECT 59.675 -217.085 60.005 -216.755 ;
        RECT 59.675 -218.445 60.005 -218.115 ;
        RECT 59.675 -224.09 60.005 -222.96 ;
        RECT 59.68 -224.205 60 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.035 132.52 61.365 133.65 ;
        RECT 61.035 128.355 61.365 128.685 ;
        RECT 61.035 126.995 61.365 127.325 ;
        RECT 61.035 125.635 61.365 125.965 ;
        RECT 61.035 124.275 61.365 124.605 ;
        RECT 61.04 123.6 61.36 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.035 -0.845 61.365 -0.515 ;
        RECT 61.035 -2.205 61.365 -1.875 ;
        RECT 61.035 -3.565 61.365 -3.235 ;
        RECT 61.04 -3.565 61.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.395 132.52 62.725 133.65 ;
        RECT 62.395 128.355 62.725 128.685 ;
        RECT 62.395 126.995 62.725 127.325 ;
        RECT 62.395 125.635 62.725 125.965 ;
        RECT 62.395 124.275 62.725 124.605 ;
        RECT 62.4 123.6 62.72 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.395 -0.845 62.725 -0.515 ;
        RECT 62.395 -2.205 62.725 -1.875 ;
        RECT 62.395 -3.565 62.725 -3.235 ;
        RECT 62.4 -3.565 62.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.395 -119.165 62.725 -118.835 ;
        RECT 62.395 -120.525 62.725 -120.195 ;
        RECT 62.395 -121.885 62.725 -121.555 ;
        RECT 62.395 -123.245 62.725 -122.915 ;
        RECT 62.395 -124.605 62.725 -124.275 ;
        RECT 62.395 -125.965 62.725 -125.635 ;
        RECT 62.395 -127.325 62.725 -126.995 ;
        RECT 62.395 -128.685 62.725 -128.355 ;
        RECT 62.395 -130.045 62.725 -129.715 ;
        RECT 62.395 -131.405 62.725 -131.075 ;
        RECT 62.395 -132.765 62.725 -132.435 ;
        RECT 62.395 -134.125 62.725 -133.795 ;
        RECT 62.395 -135.485 62.725 -135.155 ;
        RECT 62.395 -136.845 62.725 -136.515 ;
        RECT 62.395 -138.205 62.725 -137.875 ;
        RECT 62.395 -139.565 62.725 -139.235 ;
        RECT 62.395 -140.925 62.725 -140.595 ;
        RECT 62.395 -142.285 62.725 -141.955 ;
        RECT 62.395 -143.645 62.725 -143.315 ;
        RECT 62.395 -145.005 62.725 -144.675 ;
        RECT 62.395 -146.365 62.725 -146.035 ;
        RECT 62.395 -147.725 62.725 -147.395 ;
        RECT 62.395 -149.085 62.725 -148.755 ;
        RECT 62.395 -150.445 62.725 -150.115 ;
        RECT 62.395 -151.805 62.725 -151.475 ;
        RECT 62.395 -153.165 62.725 -152.835 ;
        RECT 62.395 -154.525 62.725 -154.195 ;
        RECT 62.395 -155.885 62.725 -155.555 ;
        RECT 62.395 -157.245 62.725 -156.915 ;
        RECT 62.395 -158.605 62.725 -158.275 ;
        RECT 62.395 -159.965 62.725 -159.635 ;
        RECT 62.395 -161.325 62.725 -160.995 ;
        RECT 62.395 -162.685 62.725 -162.355 ;
        RECT 62.395 -164.045 62.725 -163.715 ;
        RECT 62.395 -165.405 62.725 -165.075 ;
        RECT 62.395 -166.765 62.725 -166.435 ;
        RECT 62.395 -168.125 62.725 -167.795 ;
        RECT 62.395 -169.485 62.725 -169.155 ;
        RECT 62.395 -170.845 62.725 -170.515 ;
        RECT 62.395 -172.205 62.725 -171.875 ;
        RECT 62.395 -173.565 62.725 -173.235 ;
        RECT 62.395 -174.925 62.725 -174.595 ;
        RECT 62.395 -176.285 62.725 -175.955 ;
        RECT 62.395 -177.645 62.725 -177.315 ;
        RECT 62.395 -179.005 62.725 -178.675 ;
        RECT 62.395 -180.365 62.725 -180.035 ;
        RECT 62.395 -181.725 62.725 -181.395 ;
        RECT 62.395 -183.085 62.725 -182.755 ;
        RECT 62.395 -184.445 62.725 -184.115 ;
        RECT 62.395 -185.805 62.725 -185.475 ;
        RECT 62.395 -187.165 62.725 -186.835 ;
        RECT 62.395 -188.525 62.725 -188.195 ;
        RECT 62.395 -189.885 62.725 -189.555 ;
        RECT 62.395 -191.245 62.725 -190.915 ;
        RECT 62.395 -192.605 62.725 -192.275 ;
        RECT 62.395 -193.965 62.725 -193.635 ;
        RECT 62.395 -195.325 62.725 -194.995 ;
        RECT 62.395 -196.685 62.725 -196.355 ;
        RECT 62.395 -198.045 62.725 -197.715 ;
        RECT 62.395 -199.405 62.725 -199.075 ;
        RECT 62.395 -200.765 62.725 -200.435 ;
        RECT 62.395 -202.125 62.725 -201.795 ;
        RECT 62.395 -203.485 62.725 -203.155 ;
        RECT 62.395 -204.845 62.725 -204.515 ;
        RECT 62.395 -206.205 62.725 -205.875 ;
        RECT 62.395 -207.565 62.725 -207.235 ;
        RECT 62.395 -208.925 62.725 -208.595 ;
        RECT 62.395 -210.285 62.725 -209.955 ;
        RECT 62.395 -211.645 62.725 -211.315 ;
        RECT 62.395 -213.005 62.725 -212.675 ;
        RECT 62.395 -214.365 62.725 -214.035 ;
        RECT 62.395 -215.725 62.725 -215.395 ;
        RECT 62.395 -217.085 62.725 -216.755 ;
        RECT 62.395 -218.445 62.725 -218.115 ;
        RECT 62.395 -224.09 62.725 -222.96 ;
        RECT 62.4 -224.205 62.72 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.66 -121.535 63.99 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.755 132.52 64.085 133.65 ;
        RECT 63.755 128.355 64.085 128.685 ;
        RECT 63.755 126.995 64.085 127.325 ;
        RECT 63.755 125.635 64.085 125.965 ;
        RECT 63.755 124.275 64.085 124.605 ;
        RECT 63.76 123.6 64.08 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.755 -123.245 64.085 -122.915 ;
        RECT 63.755 -124.605 64.085 -124.275 ;
        RECT 63.755 -125.965 64.085 -125.635 ;
        RECT 63.755 -127.325 64.085 -126.995 ;
        RECT 63.755 -128.685 64.085 -128.355 ;
        RECT 63.755 -130.045 64.085 -129.715 ;
        RECT 63.755 -131.405 64.085 -131.075 ;
        RECT 63.755 -132.765 64.085 -132.435 ;
        RECT 63.755 -134.125 64.085 -133.795 ;
        RECT 63.755 -135.485 64.085 -135.155 ;
        RECT 63.755 -136.845 64.085 -136.515 ;
        RECT 63.755 -138.205 64.085 -137.875 ;
        RECT 63.755 -139.565 64.085 -139.235 ;
        RECT 63.755 -140.925 64.085 -140.595 ;
        RECT 63.755 -142.285 64.085 -141.955 ;
        RECT 63.755 -143.645 64.085 -143.315 ;
        RECT 63.755 -145.005 64.085 -144.675 ;
        RECT 63.755 -146.365 64.085 -146.035 ;
        RECT 63.755 -147.725 64.085 -147.395 ;
        RECT 63.755 -149.085 64.085 -148.755 ;
        RECT 63.755 -150.445 64.085 -150.115 ;
        RECT 63.755 -151.805 64.085 -151.475 ;
        RECT 63.755 -153.165 64.085 -152.835 ;
        RECT 63.755 -154.525 64.085 -154.195 ;
        RECT 63.755 -155.885 64.085 -155.555 ;
        RECT 63.755 -157.245 64.085 -156.915 ;
        RECT 63.755 -158.605 64.085 -158.275 ;
        RECT 63.755 -159.965 64.085 -159.635 ;
        RECT 63.755 -161.325 64.085 -160.995 ;
        RECT 63.755 -162.685 64.085 -162.355 ;
        RECT 63.755 -164.045 64.085 -163.715 ;
        RECT 63.755 -165.405 64.085 -165.075 ;
        RECT 63.755 -166.765 64.085 -166.435 ;
        RECT 63.755 -168.125 64.085 -167.795 ;
        RECT 63.755 -169.485 64.085 -169.155 ;
        RECT 63.755 -170.845 64.085 -170.515 ;
        RECT 63.755 -172.205 64.085 -171.875 ;
        RECT 63.755 -173.565 64.085 -173.235 ;
        RECT 63.755 -174.925 64.085 -174.595 ;
        RECT 63.755 -176.285 64.085 -175.955 ;
        RECT 63.755 -177.645 64.085 -177.315 ;
        RECT 63.755 -179.005 64.085 -178.675 ;
        RECT 63.755 -180.365 64.085 -180.035 ;
        RECT 63.755 -181.725 64.085 -181.395 ;
        RECT 63.755 -183.085 64.085 -182.755 ;
        RECT 63.755 -184.445 64.085 -184.115 ;
        RECT 63.755 -185.805 64.085 -185.475 ;
        RECT 63.755 -187.165 64.085 -186.835 ;
        RECT 63.755 -188.525 64.085 -188.195 ;
        RECT 63.755 -189.885 64.085 -189.555 ;
        RECT 63.755 -191.245 64.085 -190.915 ;
        RECT 63.755 -192.605 64.085 -192.275 ;
        RECT 63.755 -193.965 64.085 -193.635 ;
        RECT 63.755 -195.325 64.085 -194.995 ;
        RECT 63.755 -196.685 64.085 -196.355 ;
        RECT 63.755 -198.045 64.085 -197.715 ;
        RECT 63.755 -199.405 64.085 -199.075 ;
        RECT 63.755 -200.765 64.085 -200.435 ;
        RECT 63.755 -202.125 64.085 -201.795 ;
        RECT 63.755 -203.485 64.085 -203.155 ;
        RECT 63.755 -204.845 64.085 -204.515 ;
        RECT 63.755 -206.205 64.085 -205.875 ;
        RECT 63.755 -207.565 64.085 -207.235 ;
        RECT 63.755 -208.925 64.085 -208.595 ;
        RECT 63.755 -210.285 64.085 -209.955 ;
        RECT 63.755 -211.645 64.085 -211.315 ;
        RECT 63.755 -213.005 64.085 -212.675 ;
        RECT 63.755 -214.365 64.085 -214.035 ;
        RECT 63.755 -215.725 64.085 -215.395 ;
        RECT 63.755 -217.085 64.085 -216.755 ;
        RECT 63.755 -218.445 64.085 -218.115 ;
        RECT 63.755 -224.09 64.085 -222.96 ;
        RECT 63.76 -224.205 64.08 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.115 132.52 65.445 133.65 ;
        RECT 65.115 128.355 65.445 128.685 ;
        RECT 65.115 126.995 65.445 127.325 ;
        RECT 65.115 125.635 65.445 125.965 ;
        RECT 65.115 124.275 65.445 124.605 ;
        RECT 65.12 123.6 65.44 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.115 -0.845 65.445 -0.515 ;
        RECT 65.115 -2.205 65.445 -1.875 ;
        RECT 65.115 -3.565 65.445 -3.235 ;
        RECT 65.12 -3.565 65.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.475 132.52 66.805 133.65 ;
        RECT 66.475 128.355 66.805 128.685 ;
        RECT 66.475 126.995 66.805 127.325 ;
        RECT 66.475 125.635 66.805 125.965 ;
        RECT 66.475 124.275 66.805 124.605 ;
        RECT 66.48 123.6 66.8 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.475 -0.845 66.805 -0.515 ;
        RECT 66.475 -2.205 66.805 -1.875 ;
        RECT 66.475 -3.565 66.805 -3.235 ;
        RECT 66.48 -3.565 66.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.835 132.52 68.165 133.65 ;
        RECT 67.835 128.355 68.165 128.685 ;
        RECT 67.835 126.995 68.165 127.325 ;
        RECT 67.835 125.635 68.165 125.965 ;
        RECT 67.835 124.275 68.165 124.605 ;
        RECT 67.84 123.6 68.16 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.835 -0.845 68.165 -0.515 ;
        RECT 67.835 -2.205 68.165 -1.875 ;
        RECT 67.835 -3.565 68.165 -3.235 ;
        RECT 67.84 -3.565 68.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.835 -119.165 68.165 -118.835 ;
        RECT 67.835 -120.525 68.165 -120.195 ;
        RECT 67.835 -121.885 68.165 -121.555 ;
        RECT 67.835 -123.245 68.165 -122.915 ;
        RECT 67.835 -124.605 68.165 -124.275 ;
        RECT 67.835 -125.965 68.165 -125.635 ;
        RECT 67.835 -127.325 68.165 -126.995 ;
        RECT 67.835 -128.685 68.165 -128.355 ;
        RECT 67.835 -130.045 68.165 -129.715 ;
        RECT 67.835 -131.405 68.165 -131.075 ;
        RECT 67.835 -132.765 68.165 -132.435 ;
        RECT 67.835 -134.125 68.165 -133.795 ;
        RECT 67.835 -135.485 68.165 -135.155 ;
        RECT 67.835 -136.845 68.165 -136.515 ;
        RECT 67.835 -138.205 68.165 -137.875 ;
        RECT 67.835 -139.565 68.165 -139.235 ;
        RECT 67.835 -140.925 68.165 -140.595 ;
        RECT 67.835 -142.285 68.165 -141.955 ;
        RECT 67.835 -143.645 68.165 -143.315 ;
        RECT 67.835 -145.005 68.165 -144.675 ;
        RECT 67.835 -146.365 68.165 -146.035 ;
        RECT 67.835 -147.725 68.165 -147.395 ;
        RECT 67.835 -149.085 68.165 -148.755 ;
        RECT 67.835 -150.445 68.165 -150.115 ;
        RECT 67.835 -151.805 68.165 -151.475 ;
        RECT 67.835 -153.165 68.165 -152.835 ;
        RECT 67.835 -154.525 68.165 -154.195 ;
        RECT 67.835 -155.885 68.165 -155.555 ;
        RECT 67.835 -157.245 68.165 -156.915 ;
        RECT 67.835 -158.605 68.165 -158.275 ;
        RECT 67.835 -159.965 68.165 -159.635 ;
        RECT 67.835 -161.325 68.165 -160.995 ;
        RECT 67.835 -162.685 68.165 -162.355 ;
        RECT 67.835 -164.045 68.165 -163.715 ;
        RECT 67.835 -165.405 68.165 -165.075 ;
        RECT 67.835 -166.765 68.165 -166.435 ;
        RECT 67.835 -168.125 68.165 -167.795 ;
        RECT 67.835 -169.485 68.165 -169.155 ;
        RECT 67.835 -170.845 68.165 -170.515 ;
        RECT 67.835 -172.205 68.165 -171.875 ;
        RECT 67.835 -173.565 68.165 -173.235 ;
        RECT 67.835 -174.925 68.165 -174.595 ;
        RECT 67.835 -176.285 68.165 -175.955 ;
        RECT 67.835 -177.645 68.165 -177.315 ;
        RECT 67.835 -179.005 68.165 -178.675 ;
        RECT 67.835 -180.365 68.165 -180.035 ;
        RECT 67.835 -181.725 68.165 -181.395 ;
        RECT 67.835 -183.085 68.165 -182.755 ;
        RECT 67.835 -184.445 68.165 -184.115 ;
        RECT 67.835 -185.805 68.165 -185.475 ;
        RECT 67.835 -187.165 68.165 -186.835 ;
        RECT 67.835 -188.525 68.165 -188.195 ;
        RECT 67.835 -189.885 68.165 -189.555 ;
        RECT 67.835 -191.245 68.165 -190.915 ;
        RECT 67.835 -192.605 68.165 -192.275 ;
        RECT 67.835 -193.965 68.165 -193.635 ;
        RECT 67.835 -195.325 68.165 -194.995 ;
        RECT 67.835 -196.685 68.165 -196.355 ;
        RECT 67.835 -198.045 68.165 -197.715 ;
        RECT 67.835 -199.405 68.165 -199.075 ;
        RECT 67.835 -200.765 68.165 -200.435 ;
        RECT 67.835 -202.125 68.165 -201.795 ;
        RECT 67.835 -203.485 68.165 -203.155 ;
        RECT 67.835 -204.845 68.165 -204.515 ;
        RECT 67.835 -206.205 68.165 -205.875 ;
        RECT 67.835 -207.565 68.165 -207.235 ;
        RECT 67.835 -208.925 68.165 -208.595 ;
        RECT 67.835 -210.285 68.165 -209.955 ;
        RECT 67.835 -211.645 68.165 -211.315 ;
        RECT 67.835 -213.005 68.165 -212.675 ;
        RECT 67.835 -214.365 68.165 -214.035 ;
        RECT 67.835 -215.725 68.165 -215.395 ;
        RECT 67.835 -217.085 68.165 -216.755 ;
        RECT 67.835 -218.445 68.165 -218.115 ;
        RECT 67.835 -224.09 68.165 -222.96 ;
        RECT 67.84 -224.205 68.16 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.195 132.52 69.525 133.65 ;
        RECT 69.195 128.355 69.525 128.685 ;
        RECT 69.195 126.995 69.525 127.325 ;
        RECT 69.195 125.635 69.525 125.965 ;
        RECT 69.195 124.275 69.525 124.605 ;
        RECT 69.2 123.6 69.52 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.195 -123.245 69.525 -122.915 ;
        RECT 69.195 -124.605 69.525 -124.275 ;
        RECT 69.195 -125.965 69.525 -125.635 ;
        RECT 69.195 -127.325 69.525 -126.995 ;
        RECT 69.195 -128.685 69.525 -128.355 ;
        RECT 69.195 -130.045 69.525 -129.715 ;
        RECT 69.195 -131.405 69.525 -131.075 ;
        RECT 69.195 -132.765 69.525 -132.435 ;
        RECT 69.195 -134.125 69.525 -133.795 ;
        RECT 69.195 -135.485 69.525 -135.155 ;
        RECT 69.195 -136.845 69.525 -136.515 ;
        RECT 69.195 -138.205 69.525 -137.875 ;
        RECT 69.195 -139.565 69.525 -139.235 ;
        RECT 69.195 -140.925 69.525 -140.595 ;
        RECT 69.195 -142.285 69.525 -141.955 ;
        RECT 69.195 -143.645 69.525 -143.315 ;
        RECT 69.195 -145.005 69.525 -144.675 ;
        RECT 69.195 -146.365 69.525 -146.035 ;
        RECT 69.195 -147.725 69.525 -147.395 ;
        RECT 69.195 -149.085 69.525 -148.755 ;
        RECT 69.195 -150.445 69.525 -150.115 ;
        RECT 69.195 -151.805 69.525 -151.475 ;
        RECT 69.195 -153.165 69.525 -152.835 ;
        RECT 69.195 -154.525 69.525 -154.195 ;
        RECT 69.195 -155.885 69.525 -155.555 ;
        RECT 69.195 -157.245 69.525 -156.915 ;
        RECT 69.195 -158.605 69.525 -158.275 ;
        RECT 69.195 -159.965 69.525 -159.635 ;
        RECT 69.195 -161.325 69.525 -160.995 ;
        RECT 69.195 -162.685 69.525 -162.355 ;
        RECT 69.195 -164.045 69.525 -163.715 ;
        RECT 69.195 -165.405 69.525 -165.075 ;
        RECT 69.195 -166.765 69.525 -166.435 ;
        RECT 69.195 -168.125 69.525 -167.795 ;
        RECT 69.195 -169.485 69.525 -169.155 ;
        RECT 69.195 -170.845 69.525 -170.515 ;
        RECT 69.195 -172.205 69.525 -171.875 ;
        RECT 69.195 -173.565 69.525 -173.235 ;
        RECT 69.195 -174.925 69.525 -174.595 ;
        RECT 69.195 -176.285 69.525 -175.955 ;
        RECT 69.195 -177.645 69.525 -177.315 ;
        RECT 69.195 -179.005 69.525 -178.675 ;
        RECT 69.195 -180.365 69.525 -180.035 ;
        RECT 69.195 -181.725 69.525 -181.395 ;
        RECT 69.195 -183.085 69.525 -182.755 ;
        RECT 69.195 -184.445 69.525 -184.115 ;
        RECT 69.195 -185.805 69.525 -185.475 ;
        RECT 69.195 -187.165 69.525 -186.835 ;
        RECT 69.195 -188.525 69.525 -188.195 ;
        RECT 69.195 -189.885 69.525 -189.555 ;
        RECT 69.195 -191.245 69.525 -190.915 ;
        RECT 69.195 -192.605 69.525 -192.275 ;
        RECT 69.195 -193.965 69.525 -193.635 ;
        RECT 69.195 -195.325 69.525 -194.995 ;
        RECT 69.195 -196.685 69.525 -196.355 ;
        RECT 69.195 -198.045 69.525 -197.715 ;
        RECT 69.195 -199.405 69.525 -199.075 ;
        RECT 69.195 -200.765 69.525 -200.435 ;
        RECT 69.195 -202.125 69.525 -201.795 ;
        RECT 69.195 -203.485 69.525 -203.155 ;
        RECT 69.195 -204.845 69.525 -204.515 ;
        RECT 69.195 -206.205 69.525 -205.875 ;
        RECT 69.195 -207.565 69.525 -207.235 ;
        RECT 69.195 -208.925 69.525 -208.595 ;
        RECT 69.195 -210.285 69.525 -209.955 ;
        RECT 69.195 -211.645 69.525 -211.315 ;
        RECT 69.195 -213.005 69.525 -212.675 ;
        RECT 69.195 -214.365 69.525 -214.035 ;
        RECT 69.195 -215.725 69.525 -215.395 ;
        RECT 69.195 -217.085 69.525 -216.755 ;
        RECT 69.195 -218.445 69.525 -218.115 ;
        RECT 69.195 -224.09 69.525 -222.96 ;
        RECT 69.2 -224.205 69.52 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.76 -121.535 70.09 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.555 132.52 70.885 133.65 ;
        RECT 70.555 128.355 70.885 128.685 ;
        RECT 70.555 126.995 70.885 127.325 ;
        RECT 70.555 125.635 70.885 125.965 ;
        RECT 70.555 124.275 70.885 124.605 ;
        RECT 70.56 123.6 70.88 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 132.52 72.245 133.65 ;
        RECT 71.915 128.355 72.245 128.685 ;
        RECT 71.915 126.995 72.245 127.325 ;
        RECT 71.915 125.635 72.245 125.965 ;
        RECT 71.915 124.275 72.245 124.605 ;
        RECT 71.92 123.6 72.24 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 -0.845 72.245 -0.515 ;
        RECT 71.915 -2.205 72.245 -1.875 ;
        RECT 71.915 -3.565 72.245 -3.235 ;
        RECT 71.92 -3.565 72.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 -119.165 72.245 -118.835 ;
        RECT 71.915 -120.525 72.245 -120.195 ;
        RECT 71.915 -121.885 72.245 -121.555 ;
        RECT 71.915 -123.245 72.245 -122.915 ;
        RECT 71.915 -124.605 72.245 -124.275 ;
        RECT 71.915 -125.965 72.245 -125.635 ;
        RECT 71.915 -127.325 72.245 -126.995 ;
        RECT 71.915 -128.685 72.245 -128.355 ;
        RECT 71.915 -130.045 72.245 -129.715 ;
        RECT 71.915 -131.405 72.245 -131.075 ;
        RECT 71.915 -132.765 72.245 -132.435 ;
        RECT 71.915 -134.125 72.245 -133.795 ;
        RECT 71.915 -135.485 72.245 -135.155 ;
        RECT 71.915 -136.845 72.245 -136.515 ;
        RECT 71.915 -138.205 72.245 -137.875 ;
        RECT 71.915 -139.565 72.245 -139.235 ;
        RECT 71.915 -140.925 72.245 -140.595 ;
        RECT 71.915 -142.285 72.245 -141.955 ;
        RECT 71.915 -143.645 72.245 -143.315 ;
        RECT 71.915 -145.005 72.245 -144.675 ;
        RECT 71.915 -146.365 72.245 -146.035 ;
        RECT 71.915 -147.725 72.245 -147.395 ;
        RECT 71.915 -149.085 72.245 -148.755 ;
        RECT 71.915 -150.445 72.245 -150.115 ;
        RECT 71.915 -151.805 72.245 -151.475 ;
        RECT 71.915 -153.165 72.245 -152.835 ;
        RECT 71.915 -154.525 72.245 -154.195 ;
        RECT 71.915 -155.885 72.245 -155.555 ;
        RECT 71.915 -157.245 72.245 -156.915 ;
        RECT 71.915 -158.605 72.245 -158.275 ;
        RECT 71.915 -159.965 72.245 -159.635 ;
        RECT 71.915 -161.325 72.245 -160.995 ;
        RECT 71.915 -162.685 72.245 -162.355 ;
        RECT 71.915 -164.045 72.245 -163.715 ;
        RECT 71.915 -165.405 72.245 -165.075 ;
        RECT 71.915 -166.765 72.245 -166.435 ;
        RECT 71.915 -168.125 72.245 -167.795 ;
        RECT 71.915 -169.485 72.245 -169.155 ;
        RECT 71.915 -170.845 72.245 -170.515 ;
        RECT 71.915 -172.205 72.245 -171.875 ;
        RECT 71.915 -173.565 72.245 -173.235 ;
        RECT 71.915 -174.925 72.245 -174.595 ;
        RECT 71.915 -176.285 72.245 -175.955 ;
        RECT 71.915 -177.645 72.245 -177.315 ;
        RECT 71.915 -179.005 72.245 -178.675 ;
        RECT 71.915 -180.365 72.245 -180.035 ;
        RECT 71.915 -181.725 72.245 -181.395 ;
        RECT 71.915 -183.085 72.245 -182.755 ;
        RECT 71.915 -184.445 72.245 -184.115 ;
        RECT 71.915 -185.805 72.245 -185.475 ;
        RECT 71.915 -187.165 72.245 -186.835 ;
        RECT 71.915 -188.525 72.245 -188.195 ;
        RECT 71.915 -189.885 72.245 -189.555 ;
        RECT 71.915 -191.245 72.245 -190.915 ;
        RECT 71.915 -192.605 72.245 -192.275 ;
        RECT 71.915 -193.965 72.245 -193.635 ;
        RECT 71.915 -195.325 72.245 -194.995 ;
        RECT 71.915 -196.685 72.245 -196.355 ;
        RECT 71.915 -198.045 72.245 -197.715 ;
        RECT 71.915 -199.405 72.245 -199.075 ;
        RECT 71.915 -200.765 72.245 -200.435 ;
        RECT 71.915 -202.125 72.245 -201.795 ;
        RECT 71.915 -203.485 72.245 -203.155 ;
        RECT 71.915 -204.845 72.245 -204.515 ;
        RECT 71.915 -206.205 72.245 -205.875 ;
        RECT 71.915 -207.565 72.245 -207.235 ;
        RECT 71.915 -208.925 72.245 -208.595 ;
        RECT 71.915 -210.285 72.245 -209.955 ;
        RECT 71.915 -211.645 72.245 -211.315 ;
        RECT 71.915 -213.005 72.245 -212.675 ;
        RECT 71.915 -214.365 72.245 -214.035 ;
        RECT 71.915 -215.725 72.245 -215.395 ;
        RECT 71.915 -217.085 72.245 -216.755 ;
        RECT 71.915 -218.445 72.245 -218.115 ;
        RECT 71.915 -224.09 72.245 -222.96 ;
        RECT 71.92 -224.205 72.24 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.275 132.52 73.605 133.65 ;
        RECT 73.275 128.355 73.605 128.685 ;
        RECT 73.275 126.995 73.605 127.325 ;
        RECT 73.275 125.635 73.605 125.965 ;
        RECT 73.275 124.275 73.605 124.605 ;
        RECT 73.28 123.6 73.6 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.275 -0.845 73.605 -0.515 ;
        RECT 73.275 -2.205 73.605 -1.875 ;
        RECT 73.275 -3.565 73.605 -3.235 ;
        RECT 73.28 -3.565 73.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.635 132.52 74.965 133.65 ;
        RECT 74.635 128.355 74.965 128.685 ;
        RECT 74.635 126.995 74.965 127.325 ;
        RECT 74.635 125.635 74.965 125.965 ;
        RECT 74.635 124.275 74.965 124.605 ;
        RECT 74.64 123.6 74.96 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.635 -0.845 74.965 -0.515 ;
        RECT 74.635 -2.205 74.965 -1.875 ;
        RECT 74.635 -3.565 74.965 -3.235 ;
        RECT 74.64 -3.565 74.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.635 -138.205 74.965 -137.875 ;
        RECT 74.635 -139.565 74.965 -139.235 ;
        RECT 74.635 -140.925 74.965 -140.595 ;
        RECT 74.635 -142.285 74.965 -141.955 ;
        RECT 74.635 -143.645 74.965 -143.315 ;
        RECT 74.635 -145.005 74.965 -144.675 ;
        RECT 74.635 -146.365 74.965 -146.035 ;
        RECT 74.635 -147.725 74.965 -147.395 ;
        RECT 74.635 -149.085 74.965 -148.755 ;
        RECT 74.635 -150.445 74.965 -150.115 ;
        RECT 74.635 -151.805 74.965 -151.475 ;
        RECT 74.635 -153.165 74.965 -152.835 ;
        RECT 74.635 -154.525 74.965 -154.195 ;
        RECT 74.635 -155.885 74.965 -155.555 ;
        RECT 74.635 -157.245 74.965 -156.915 ;
        RECT 74.635 -158.605 74.965 -158.275 ;
        RECT 74.635 -159.965 74.965 -159.635 ;
        RECT 74.635 -161.325 74.965 -160.995 ;
        RECT 74.635 -162.685 74.965 -162.355 ;
        RECT 74.635 -164.045 74.965 -163.715 ;
        RECT 74.635 -165.405 74.965 -165.075 ;
        RECT 74.635 -166.765 74.965 -166.435 ;
        RECT 74.635 -168.125 74.965 -167.795 ;
        RECT 74.635 -169.485 74.965 -169.155 ;
        RECT 74.635 -170.845 74.965 -170.515 ;
        RECT 74.635 -172.205 74.965 -171.875 ;
        RECT 74.635 -173.565 74.965 -173.235 ;
        RECT 74.635 -174.925 74.965 -174.595 ;
        RECT 74.635 -176.285 74.965 -175.955 ;
        RECT 74.635 -177.645 74.965 -177.315 ;
        RECT 74.635 -179.005 74.965 -178.675 ;
        RECT 74.635 -180.365 74.965 -180.035 ;
        RECT 74.635 -181.725 74.965 -181.395 ;
        RECT 74.635 -183.085 74.965 -182.755 ;
        RECT 74.635 -184.445 74.965 -184.115 ;
        RECT 74.635 -185.805 74.965 -185.475 ;
        RECT 74.635 -187.165 74.965 -186.835 ;
        RECT 74.635 -188.525 74.965 -188.195 ;
        RECT 74.635 -189.885 74.965 -189.555 ;
        RECT 74.635 -191.245 74.965 -190.915 ;
        RECT 74.635 -192.605 74.965 -192.275 ;
        RECT 74.635 -193.965 74.965 -193.635 ;
        RECT 74.635 -195.325 74.965 -194.995 ;
        RECT 74.635 -196.685 74.965 -196.355 ;
        RECT 74.635 -198.045 74.965 -197.715 ;
        RECT 74.635 -199.405 74.965 -199.075 ;
        RECT 74.635 -200.765 74.965 -200.435 ;
        RECT 74.635 -202.125 74.965 -201.795 ;
        RECT 74.635 -203.485 74.965 -203.155 ;
        RECT 74.635 -204.845 74.965 -204.515 ;
        RECT 74.635 -206.205 74.965 -205.875 ;
        RECT 74.635 -207.565 74.965 -207.235 ;
        RECT 74.635 -208.925 74.965 -208.595 ;
        RECT 74.635 -210.285 74.965 -209.955 ;
        RECT 74.635 -211.645 74.965 -211.315 ;
        RECT 74.635 -213.005 74.965 -212.675 ;
        RECT 74.635 -214.365 74.965 -214.035 ;
        RECT 74.635 -215.725 74.965 -215.395 ;
        RECT 74.635 -217.085 74.965 -216.755 ;
        RECT 74.635 -218.445 74.965 -218.115 ;
        RECT 74.635 -224.09 74.965 -222.96 ;
        RECT 74.64 -224.205 74.96 -118.16 ;
        RECT 74.635 -119.165 74.965 -118.835 ;
        RECT 74.635 -120.525 74.965 -120.195 ;
        RECT 74.635 -121.885 74.965 -121.555 ;
        RECT 74.635 -123.245 74.965 -122.915 ;
        RECT 74.635 -124.605 74.965 -124.275 ;
        RECT 74.635 -125.965 74.965 -125.635 ;
        RECT 74.635 -127.325 74.965 -126.995 ;
        RECT 74.635 -128.685 74.965 -128.355 ;
        RECT 74.635 -130.045 74.965 -129.715 ;
        RECT 74.635 -131.405 74.965 -131.075 ;
        RECT 74.635 -132.765 74.965 -132.435 ;
        RECT 74.635 -134.125 74.965 -133.795 ;
        RECT 74.635 -135.485 74.965 -135.155 ;
        RECT 74.635 -136.845 74.965 -136.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.86 -121.535 15.19 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.155 132.52 16.485 133.65 ;
        RECT 16.155 128.355 16.485 128.685 ;
        RECT 16.155 126.995 16.485 127.325 ;
        RECT 16.155 125.635 16.485 125.965 ;
        RECT 16.155 124.275 16.485 124.605 ;
        RECT 16.16 123.6 16.48 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.515 132.52 17.845 133.65 ;
        RECT 17.515 128.355 17.845 128.685 ;
        RECT 17.515 126.995 17.845 127.325 ;
        RECT 17.515 125.635 17.845 125.965 ;
        RECT 17.515 124.275 17.845 124.605 ;
        RECT 17.52 123.6 17.84 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.515 -0.845 17.845 -0.515 ;
        RECT 17.515 -2.205 17.845 -1.875 ;
        RECT 17.515 -3.565 17.845 -3.235 ;
        RECT 17.52 -3.565 17.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.875 132.52 19.205 133.65 ;
        RECT 18.875 128.355 19.205 128.685 ;
        RECT 18.875 126.995 19.205 127.325 ;
        RECT 18.875 125.635 19.205 125.965 ;
        RECT 18.875 124.275 19.205 124.605 ;
        RECT 18.88 123.6 19.2 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.875 -0.845 19.205 -0.515 ;
        RECT 18.875 -2.205 19.205 -1.875 ;
        RECT 18.875 -3.565 19.205 -3.235 ;
        RECT 18.88 -3.565 19.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.875 -119.165 19.205 -118.835 ;
        RECT 18.875 -120.525 19.205 -120.195 ;
        RECT 18.875 -121.885 19.205 -121.555 ;
        RECT 18.875 -123.245 19.205 -122.915 ;
        RECT 18.875 -124.605 19.205 -124.275 ;
        RECT 18.875 -125.965 19.205 -125.635 ;
        RECT 18.875 -127.325 19.205 -126.995 ;
        RECT 18.875 -128.685 19.205 -128.355 ;
        RECT 18.875 -130.045 19.205 -129.715 ;
        RECT 18.875 -131.405 19.205 -131.075 ;
        RECT 18.875 -132.765 19.205 -132.435 ;
        RECT 18.875 -134.125 19.205 -133.795 ;
        RECT 18.875 -135.485 19.205 -135.155 ;
        RECT 18.875 -136.845 19.205 -136.515 ;
        RECT 18.875 -138.205 19.205 -137.875 ;
        RECT 18.875 -139.565 19.205 -139.235 ;
        RECT 18.875 -140.925 19.205 -140.595 ;
        RECT 18.875 -142.285 19.205 -141.955 ;
        RECT 18.875 -143.645 19.205 -143.315 ;
        RECT 18.875 -145.005 19.205 -144.675 ;
        RECT 18.875 -146.365 19.205 -146.035 ;
        RECT 18.875 -147.725 19.205 -147.395 ;
        RECT 18.875 -149.085 19.205 -148.755 ;
        RECT 18.875 -150.445 19.205 -150.115 ;
        RECT 18.875 -151.805 19.205 -151.475 ;
        RECT 18.875 -153.165 19.205 -152.835 ;
        RECT 18.875 -154.525 19.205 -154.195 ;
        RECT 18.875 -155.885 19.205 -155.555 ;
        RECT 18.875 -157.245 19.205 -156.915 ;
        RECT 18.875 -158.605 19.205 -158.275 ;
        RECT 18.875 -159.965 19.205 -159.635 ;
        RECT 18.875 -161.325 19.205 -160.995 ;
        RECT 18.875 -162.685 19.205 -162.355 ;
        RECT 18.875 -164.045 19.205 -163.715 ;
        RECT 18.875 -165.405 19.205 -165.075 ;
        RECT 18.875 -166.765 19.205 -166.435 ;
        RECT 18.875 -168.125 19.205 -167.795 ;
        RECT 18.875 -169.485 19.205 -169.155 ;
        RECT 18.875 -170.845 19.205 -170.515 ;
        RECT 18.875 -172.205 19.205 -171.875 ;
        RECT 18.875 -173.565 19.205 -173.235 ;
        RECT 18.875 -174.925 19.205 -174.595 ;
        RECT 18.875 -176.285 19.205 -175.955 ;
        RECT 18.875 -177.645 19.205 -177.315 ;
        RECT 18.875 -179.005 19.205 -178.675 ;
        RECT 18.875 -180.365 19.205 -180.035 ;
        RECT 18.875 -181.725 19.205 -181.395 ;
        RECT 18.875 -183.085 19.205 -182.755 ;
        RECT 18.875 -184.445 19.205 -184.115 ;
        RECT 18.875 -185.805 19.205 -185.475 ;
        RECT 18.875 -187.165 19.205 -186.835 ;
        RECT 18.875 -188.525 19.205 -188.195 ;
        RECT 18.875 -189.885 19.205 -189.555 ;
        RECT 18.875 -191.245 19.205 -190.915 ;
        RECT 18.875 -192.605 19.205 -192.275 ;
        RECT 18.875 -193.965 19.205 -193.635 ;
        RECT 18.875 -195.325 19.205 -194.995 ;
        RECT 18.875 -196.685 19.205 -196.355 ;
        RECT 18.875 -198.045 19.205 -197.715 ;
        RECT 18.875 -199.405 19.205 -199.075 ;
        RECT 18.875 -200.765 19.205 -200.435 ;
        RECT 18.875 -202.125 19.205 -201.795 ;
        RECT 18.875 -203.485 19.205 -203.155 ;
        RECT 18.875 -204.845 19.205 -204.515 ;
        RECT 18.875 -206.205 19.205 -205.875 ;
        RECT 18.875 -207.565 19.205 -207.235 ;
        RECT 18.875 -208.925 19.205 -208.595 ;
        RECT 18.875 -210.285 19.205 -209.955 ;
        RECT 18.875 -211.645 19.205 -211.315 ;
        RECT 18.875 -213.005 19.205 -212.675 ;
        RECT 18.875 -214.365 19.205 -214.035 ;
        RECT 18.875 -215.725 19.205 -215.395 ;
        RECT 18.875 -217.085 19.205 -216.755 ;
        RECT 18.875 -218.445 19.205 -218.115 ;
        RECT 18.875 -224.09 19.205 -222.96 ;
        RECT 18.88 -224.205 19.2 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.235 132.52 20.565 133.65 ;
        RECT 20.235 128.355 20.565 128.685 ;
        RECT 20.235 126.995 20.565 127.325 ;
        RECT 20.235 125.635 20.565 125.965 ;
        RECT 20.235 124.275 20.565 124.605 ;
        RECT 20.24 123.6 20.56 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.235 -0.845 20.565 -0.515 ;
        RECT 20.235 -2.205 20.565 -1.875 ;
        RECT 20.235 -3.565 20.565 -3.235 ;
        RECT 20.24 -3.565 20.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.235 -119.165 20.565 -118.835 ;
        RECT 20.235 -120.525 20.565 -120.195 ;
        RECT 20.235 -121.885 20.565 -121.555 ;
        RECT 20.235 -123.245 20.565 -122.915 ;
        RECT 20.235 -124.605 20.565 -124.275 ;
        RECT 20.235 -125.965 20.565 -125.635 ;
        RECT 20.235 -127.325 20.565 -126.995 ;
        RECT 20.235 -128.685 20.565 -128.355 ;
        RECT 20.235 -130.045 20.565 -129.715 ;
        RECT 20.235 -131.405 20.565 -131.075 ;
        RECT 20.235 -132.765 20.565 -132.435 ;
        RECT 20.235 -134.125 20.565 -133.795 ;
        RECT 20.235 -135.485 20.565 -135.155 ;
        RECT 20.235 -136.845 20.565 -136.515 ;
        RECT 20.235 -138.205 20.565 -137.875 ;
        RECT 20.235 -139.565 20.565 -139.235 ;
        RECT 20.235 -140.925 20.565 -140.595 ;
        RECT 20.235 -142.285 20.565 -141.955 ;
        RECT 20.235 -143.645 20.565 -143.315 ;
        RECT 20.235 -145.005 20.565 -144.675 ;
        RECT 20.235 -146.365 20.565 -146.035 ;
        RECT 20.235 -147.725 20.565 -147.395 ;
        RECT 20.235 -149.085 20.565 -148.755 ;
        RECT 20.235 -150.445 20.565 -150.115 ;
        RECT 20.235 -151.805 20.565 -151.475 ;
        RECT 20.235 -153.165 20.565 -152.835 ;
        RECT 20.235 -154.525 20.565 -154.195 ;
        RECT 20.235 -155.885 20.565 -155.555 ;
        RECT 20.235 -157.245 20.565 -156.915 ;
        RECT 20.235 -158.605 20.565 -158.275 ;
        RECT 20.235 -159.965 20.565 -159.635 ;
        RECT 20.235 -161.325 20.565 -160.995 ;
        RECT 20.235 -162.685 20.565 -162.355 ;
        RECT 20.235 -164.045 20.565 -163.715 ;
        RECT 20.235 -165.405 20.565 -165.075 ;
        RECT 20.235 -166.765 20.565 -166.435 ;
        RECT 20.235 -168.125 20.565 -167.795 ;
        RECT 20.235 -169.485 20.565 -169.155 ;
        RECT 20.235 -170.845 20.565 -170.515 ;
        RECT 20.235 -172.205 20.565 -171.875 ;
        RECT 20.235 -173.565 20.565 -173.235 ;
        RECT 20.235 -174.925 20.565 -174.595 ;
        RECT 20.235 -176.285 20.565 -175.955 ;
        RECT 20.235 -177.645 20.565 -177.315 ;
        RECT 20.235 -179.005 20.565 -178.675 ;
        RECT 20.235 -180.365 20.565 -180.035 ;
        RECT 20.235 -181.725 20.565 -181.395 ;
        RECT 20.235 -183.085 20.565 -182.755 ;
        RECT 20.235 -184.445 20.565 -184.115 ;
        RECT 20.235 -185.805 20.565 -185.475 ;
        RECT 20.235 -187.165 20.565 -186.835 ;
        RECT 20.235 -188.525 20.565 -188.195 ;
        RECT 20.235 -189.885 20.565 -189.555 ;
        RECT 20.235 -191.245 20.565 -190.915 ;
        RECT 20.235 -192.605 20.565 -192.275 ;
        RECT 20.235 -193.965 20.565 -193.635 ;
        RECT 20.235 -195.325 20.565 -194.995 ;
        RECT 20.235 -196.685 20.565 -196.355 ;
        RECT 20.235 -198.045 20.565 -197.715 ;
        RECT 20.235 -199.405 20.565 -199.075 ;
        RECT 20.235 -200.765 20.565 -200.435 ;
        RECT 20.235 -202.125 20.565 -201.795 ;
        RECT 20.235 -203.485 20.565 -203.155 ;
        RECT 20.235 -204.845 20.565 -204.515 ;
        RECT 20.235 -206.205 20.565 -205.875 ;
        RECT 20.235 -207.565 20.565 -207.235 ;
        RECT 20.235 -208.925 20.565 -208.595 ;
        RECT 20.235 -210.285 20.565 -209.955 ;
        RECT 20.235 -211.645 20.565 -211.315 ;
        RECT 20.235 -213.005 20.565 -212.675 ;
        RECT 20.235 -214.365 20.565 -214.035 ;
        RECT 20.235 -215.725 20.565 -215.395 ;
        RECT 20.235 -217.085 20.565 -216.755 ;
        RECT 20.235 -218.445 20.565 -218.115 ;
        RECT 20.235 -224.09 20.565 -222.96 ;
        RECT 20.24 -224.205 20.56 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.96 -121.535 21.29 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.595 132.52 21.925 133.65 ;
        RECT 21.595 128.355 21.925 128.685 ;
        RECT 21.595 126.995 21.925 127.325 ;
        RECT 21.595 125.635 21.925 125.965 ;
        RECT 21.595 124.275 21.925 124.605 ;
        RECT 21.6 123.6 21.92 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.595 -123.245 21.925 -122.915 ;
        RECT 21.595 -124.605 21.925 -124.275 ;
        RECT 21.595 -125.965 21.925 -125.635 ;
        RECT 21.595 -127.325 21.925 -126.995 ;
        RECT 21.595 -128.685 21.925 -128.355 ;
        RECT 21.595 -130.045 21.925 -129.715 ;
        RECT 21.595 -131.405 21.925 -131.075 ;
        RECT 21.595 -132.765 21.925 -132.435 ;
        RECT 21.595 -134.125 21.925 -133.795 ;
        RECT 21.595 -135.485 21.925 -135.155 ;
        RECT 21.595 -136.845 21.925 -136.515 ;
        RECT 21.595 -138.205 21.925 -137.875 ;
        RECT 21.595 -139.565 21.925 -139.235 ;
        RECT 21.595 -140.925 21.925 -140.595 ;
        RECT 21.595 -142.285 21.925 -141.955 ;
        RECT 21.595 -143.645 21.925 -143.315 ;
        RECT 21.595 -145.005 21.925 -144.675 ;
        RECT 21.595 -146.365 21.925 -146.035 ;
        RECT 21.595 -147.725 21.925 -147.395 ;
        RECT 21.595 -149.085 21.925 -148.755 ;
        RECT 21.595 -150.445 21.925 -150.115 ;
        RECT 21.595 -151.805 21.925 -151.475 ;
        RECT 21.595 -153.165 21.925 -152.835 ;
        RECT 21.595 -154.525 21.925 -154.195 ;
        RECT 21.595 -155.885 21.925 -155.555 ;
        RECT 21.595 -157.245 21.925 -156.915 ;
        RECT 21.595 -158.605 21.925 -158.275 ;
        RECT 21.595 -159.965 21.925 -159.635 ;
        RECT 21.595 -161.325 21.925 -160.995 ;
        RECT 21.595 -162.685 21.925 -162.355 ;
        RECT 21.595 -164.045 21.925 -163.715 ;
        RECT 21.595 -165.405 21.925 -165.075 ;
        RECT 21.595 -166.765 21.925 -166.435 ;
        RECT 21.595 -168.125 21.925 -167.795 ;
        RECT 21.595 -169.485 21.925 -169.155 ;
        RECT 21.595 -170.845 21.925 -170.515 ;
        RECT 21.595 -172.205 21.925 -171.875 ;
        RECT 21.595 -173.565 21.925 -173.235 ;
        RECT 21.595 -174.925 21.925 -174.595 ;
        RECT 21.595 -176.285 21.925 -175.955 ;
        RECT 21.595 -177.645 21.925 -177.315 ;
        RECT 21.595 -179.005 21.925 -178.675 ;
        RECT 21.595 -180.365 21.925 -180.035 ;
        RECT 21.595 -181.725 21.925 -181.395 ;
        RECT 21.595 -183.085 21.925 -182.755 ;
        RECT 21.595 -184.445 21.925 -184.115 ;
        RECT 21.595 -185.805 21.925 -185.475 ;
        RECT 21.595 -187.165 21.925 -186.835 ;
        RECT 21.595 -188.525 21.925 -188.195 ;
        RECT 21.595 -189.885 21.925 -189.555 ;
        RECT 21.595 -191.245 21.925 -190.915 ;
        RECT 21.595 -192.605 21.925 -192.275 ;
        RECT 21.595 -193.965 21.925 -193.635 ;
        RECT 21.595 -195.325 21.925 -194.995 ;
        RECT 21.595 -196.685 21.925 -196.355 ;
        RECT 21.595 -198.045 21.925 -197.715 ;
        RECT 21.595 -199.405 21.925 -199.075 ;
        RECT 21.595 -200.765 21.925 -200.435 ;
        RECT 21.595 -202.125 21.925 -201.795 ;
        RECT 21.595 -203.485 21.925 -203.155 ;
        RECT 21.595 -204.845 21.925 -204.515 ;
        RECT 21.595 -206.205 21.925 -205.875 ;
        RECT 21.595 -207.565 21.925 -207.235 ;
        RECT 21.595 -208.925 21.925 -208.595 ;
        RECT 21.595 -210.285 21.925 -209.955 ;
        RECT 21.595 -211.645 21.925 -211.315 ;
        RECT 21.595 -213.005 21.925 -212.675 ;
        RECT 21.595 -214.365 21.925 -214.035 ;
        RECT 21.595 -215.725 21.925 -215.395 ;
        RECT 21.595 -217.085 21.925 -216.755 ;
        RECT 21.595 -218.445 21.925 -218.115 ;
        RECT 21.595 -224.09 21.925 -222.96 ;
        RECT 21.6 -224.205 21.92 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.955 132.52 23.285 133.65 ;
        RECT 22.955 128.355 23.285 128.685 ;
        RECT 22.955 126.995 23.285 127.325 ;
        RECT 22.955 125.635 23.285 125.965 ;
        RECT 22.955 124.275 23.285 124.605 ;
        RECT 22.96 123.6 23.28 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.955 -0.845 23.285 -0.515 ;
        RECT 22.955 -2.205 23.285 -1.875 ;
        RECT 22.955 -3.565 23.285 -3.235 ;
        RECT 22.96 -3.565 23.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.315 132.52 24.645 133.65 ;
        RECT 24.315 128.355 24.645 128.685 ;
        RECT 24.315 126.995 24.645 127.325 ;
        RECT 24.315 125.635 24.645 125.965 ;
        RECT 24.315 124.275 24.645 124.605 ;
        RECT 24.32 123.6 24.64 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.315 -0.845 24.645 -0.515 ;
        RECT 24.315 -2.205 24.645 -1.875 ;
        RECT 24.315 -3.565 24.645 -3.235 ;
        RECT 24.32 -3.565 24.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.675 132.52 26.005 133.65 ;
        RECT 25.675 128.355 26.005 128.685 ;
        RECT 25.675 126.995 26.005 127.325 ;
        RECT 25.675 125.635 26.005 125.965 ;
        RECT 25.675 124.275 26.005 124.605 ;
        RECT 25.68 123.6 26 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.675 -0.845 26.005 -0.515 ;
        RECT 25.675 -2.205 26.005 -1.875 ;
        RECT 25.675 -3.565 26.005 -3.235 ;
        RECT 25.68 -3.565 26 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.675 -119.165 26.005 -118.835 ;
        RECT 25.675 -120.525 26.005 -120.195 ;
        RECT 25.675 -121.885 26.005 -121.555 ;
        RECT 25.675 -123.245 26.005 -122.915 ;
        RECT 25.675 -124.605 26.005 -124.275 ;
        RECT 25.675 -125.965 26.005 -125.635 ;
        RECT 25.675 -127.325 26.005 -126.995 ;
        RECT 25.675 -128.685 26.005 -128.355 ;
        RECT 25.675 -130.045 26.005 -129.715 ;
        RECT 25.675 -131.405 26.005 -131.075 ;
        RECT 25.675 -132.765 26.005 -132.435 ;
        RECT 25.675 -134.125 26.005 -133.795 ;
        RECT 25.675 -135.485 26.005 -135.155 ;
        RECT 25.675 -136.845 26.005 -136.515 ;
        RECT 25.675 -138.205 26.005 -137.875 ;
        RECT 25.675 -139.565 26.005 -139.235 ;
        RECT 25.675 -140.925 26.005 -140.595 ;
        RECT 25.675 -142.285 26.005 -141.955 ;
        RECT 25.675 -143.645 26.005 -143.315 ;
        RECT 25.675 -145.005 26.005 -144.675 ;
        RECT 25.675 -146.365 26.005 -146.035 ;
        RECT 25.675 -147.725 26.005 -147.395 ;
        RECT 25.675 -149.085 26.005 -148.755 ;
        RECT 25.675 -150.445 26.005 -150.115 ;
        RECT 25.675 -151.805 26.005 -151.475 ;
        RECT 25.675 -153.165 26.005 -152.835 ;
        RECT 25.675 -154.525 26.005 -154.195 ;
        RECT 25.675 -155.885 26.005 -155.555 ;
        RECT 25.675 -157.245 26.005 -156.915 ;
        RECT 25.675 -158.605 26.005 -158.275 ;
        RECT 25.675 -159.965 26.005 -159.635 ;
        RECT 25.675 -161.325 26.005 -160.995 ;
        RECT 25.675 -162.685 26.005 -162.355 ;
        RECT 25.675 -164.045 26.005 -163.715 ;
        RECT 25.675 -165.405 26.005 -165.075 ;
        RECT 25.675 -166.765 26.005 -166.435 ;
        RECT 25.675 -168.125 26.005 -167.795 ;
        RECT 25.675 -169.485 26.005 -169.155 ;
        RECT 25.675 -170.845 26.005 -170.515 ;
        RECT 25.675 -172.205 26.005 -171.875 ;
        RECT 25.675 -173.565 26.005 -173.235 ;
        RECT 25.675 -174.925 26.005 -174.595 ;
        RECT 25.675 -176.285 26.005 -175.955 ;
        RECT 25.675 -177.645 26.005 -177.315 ;
        RECT 25.675 -179.005 26.005 -178.675 ;
        RECT 25.675 -180.365 26.005 -180.035 ;
        RECT 25.675 -181.725 26.005 -181.395 ;
        RECT 25.675 -183.085 26.005 -182.755 ;
        RECT 25.675 -184.445 26.005 -184.115 ;
        RECT 25.675 -185.805 26.005 -185.475 ;
        RECT 25.675 -187.165 26.005 -186.835 ;
        RECT 25.675 -188.525 26.005 -188.195 ;
        RECT 25.675 -189.885 26.005 -189.555 ;
        RECT 25.675 -191.245 26.005 -190.915 ;
        RECT 25.675 -192.605 26.005 -192.275 ;
        RECT 25.675 -193.965 26.005 -193.635 ;
        RECT 25.675 -195.325 26.005 -194.995 ;
        RECT 25.675 -196.685 26.005 -196.355 ;
        RECT 25.675 -198.045 26.005 -197.715 ;
        RECT 25.675 -199.405 26.005 -199.075 ;
        RECT 25.675 -200.765 26.005 -200.435 ;
        RECT 25.675 -202.125 26.005 -201.795 ;
        RECT 25.675 -203.485 26.005 -203.155 ;
        RECT 25.675 -204.845 26.005 -204.515 ;
        RECT 25.675 -206.205 26.005 -205.875 ;
        RECT 25.675 -207.565 26.005 -207.235 ;
        RECT 25.675 -208.925 26.005 -208.595 ;
        RECT 25.675 -210.285 26.005 -209.955 ;
        RECT 25.675 -211.645 26.005 -211.315 ;
        RECT 25.675 -213.005 26.005 -212.675 ;
        RECT 25.675 -214.365 26.005 -214.035 ;
        RECT 25.675 -215.725 26.005 -215.395 ;
        RECT 25.675 -217.085 26.005 -216.755 ;
        RECT 25.675 -218.445 26.005 -218.115 ;
        RECT 25.675 -224.09 26.005 -222.96 ;
        RECT 25.68 -224.205 26 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.035 132.52 27.365 133.65 ;
        RECT 27.035 128.355 27.365 128.685 ;
        RECT 27.035 126.995 27.365 127.325 ;
        RECT 27.035 125.635 27.365 125.965 ;
        RECT 27.035 124.275 27.365 124.605 ;
        RECT 27.04 123.6 27.36 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.035 -123.245 27.365 -122.915 ;
        RECT 27.035 -124.605 27.365 -124.275 ;
        RECT 27.035 -125.965 27.365 -125.635 ;
        RECT 27.035 -127.325 27.365 -126.995 ;
        RECT 27.035 -128.685 27.365 -128.355 ;
        RECT 27.035 -130.045 27.365 -129.715 ;
        RECT 27.035 -131.405 27.365 -131.075 ;
        RECT 27.035 -132.765 27.365 -132.435 ;
        RECT 27.035 -134.125 27.365 -133.795 ;
        RECT 27.035 -135.485 27.365 -135.155 ;
        RECT 27.035 -136.845 27.365 -136.515 ;
        RECT 27.035 -138.205 27.365 -137.875 ;
        RECT 27.035 -139.565 27.365 -139.235 ;
        RECT 27.035 -140.925 27.365 -140.595 ;
        RECT 27.035 -142.285 27.365 -141.955 ;
        RECT 27.035 -143.645 27.365 -143.315 ;
        RECT 27.035 -145.005 27.365 -144.675 ;
        RECT 27.035 -146.365 27.365 -146.035 ;
        RECT 27.035 -147.725 27.365 -147.395 ;
        RECT 27.035 -149.085 27.365 -148.755 ;
        RECT 27.035 -150.445 27.365 -150.115 ;
        RECT 27.035 -151.805 27.365 -151.475 ;
        RECT 27.035 -153.165 27.365 -152.835 ;
        RECT 27.035 -154.525 27.365 -154.195 ;
        RECT 27.035 -155.885 27.365 -155.555 ;
        RECT 27.035 -157.245 27.365 -156.915 ;
        RECT 27.035 -158.605 27.365 -158.275 ;
        RECT 27.035 -159.965 27.365 -159.635 ;
        RECT 27.035 -161.325 27.365 -160.995 ;
        RECT 27.035 -162.685 27.365 -162.355 ;
        RECT 27.035 -164.045 27.365 -163.715 ;
        RECT 27.035 -165.405 27.365 -165.075 ;
        RECT 27.035 -166.765 27.365 -166.435 ;
        RECT 27.035 -168.125 27.365 -167.795 ;
        RECT 27.035 -169.485 27.365 -169.155 ;
        RECT 27.035 -170.845 27.365 -170.515 ;
        RECT 27.035 -172.205 27.365 -171.875 ;
        RECT 27.035 -173.565 27.365 -173.235 ;
        RECT 27.035 -174.925 27.365 -174.595 ;
        RECT 27.035 -176.285 27.365 -175.955 ;
        RECT 27.035 -177.645 27.365 -177.315 ;
        RECT 27.035 -179.005 27.365 -178.675 ;
        RECT 27.035 -180.365 27.365 -180.035 ;
        RECT 27.035 -181.725 27.365 -181.395 ;
        RECT 27.035 -183.085 27.365 -182.755 ;
        RECT 27.035 -184.445 27.365 -184.115 ;
        RECT 27.035 -185.805 27.365 -185.475 ;
        RECT 27.035 -187.165 27.365 -186.835 ;
        RECT 27.035 -188.525 27.365 -188.195 ;
        RECT 27.035 -189.885 27.365 -189.555 ;
        RECT 27.035 -191.245 27.365 -190.915 ;
        RECT 27.035 -192.605 27.365 -192.275 ;
        RECT 27.035 -193.965 27.365 -193.635 ;
        RECT 27.035 -195.325 27.365 -194.995 ;
        RECT 27.035 -196.685 27.365 -196.355 ;
        RECT 27.035 -198.045 27.365 -197.715 ;
        RECT 27.035 -199.405 27.365 -199.075 ;
        RECT 27.035 -200.765 27.365 -200.435 ;
        RECT 27.035 -202.125 27.365 -201.795 ;
        RECT 27.035 -203.485 27.365 -203.155 ;
        RECT 27.035 -204.845 27.365 -204.515 ;
        RECT 27.035 -206.205 27.365 -205.875 ;
        RECT 27.035 -207.565 27.365 -207.235 ;
        RECT 27.035 -208.925 27.365 -208.595 ;
        RECT 27.035 -210.285 27.365 -209.955 ;
        RECT 27.035 -211.645 27.365 -211.315 ;
        RECT 27.035 -213.005 27.365 -212.675 ;
        RECT 27.035 -214.365 27.365 -214.035 ;
        RECT 27.035 -215.725 27.365 -215.395 ;
        RECT 27.035 -217.085 27.365 -216.755 ;
        RECT 27.035 -218.445 27.365 -218.115 ;
        RECT 27.035 -224.09 27.365 -222.96 ;
        RECT 27.04 -224.205 27.36 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.06 -121.535 27.39 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.395 132.52 28.725 133.65 ;
        RECT 28.395 128.355 28.725 128.685 ;
        RECT 28.395 126.995 28.725 127.325 ;
        RECT 28.395 125.635 28.725 125.965 ;
        RECT 28.395 124.275 28.725 124.605 ;
        RECT 28.4 123.6 28.72 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.395 -0.845 28.725 -0.515 ;
        RECT 28.395 -2.205 28.725 -1.875 ;
        RECT 28.395 -3.565 28.725 -3.235 ;
        RECT 28.4 -3.565 28.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.755 132.52 30.085 133.65 ;
        RECT 29.755 128.355 30.085 128.685 ;
        RECT 29.755 126.995 30.085 127.325 ;
        RECT 29.755 125.635 30.085 125.965 ;
        RECT 29.755 124.275 30.085 124.605 ;
        RECT 29.76 123.6 30.08 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.755 -0.845 30.085 -0.515 ;
        RECT 29.755 -2.205 30.085 -1.875 ;
        RECT 29.755 -3.565 30.085 -3.235 ;
        RECT 29.76 -3.565 30.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.115 132.52 31.445 133.65 ;
        RECT 31.115 128.355 31.445 128.685 ;
        RECT 31.115 126.995 31.445 127.325 ;
        RECT 31.115 125.635 31.445 125.965 ;
        RECT 31.115 124.275 31.445 124.605 ;
        RECT 31.12 123.6 31.44 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.115 -0.845 31.445 -0.515 ;
        RECT 31.115 -2.205 31.445 -1.875 ;
        RECT 31.115 -3.565 31.445 -3.235 ;
        RECT 31.12 -3.565 31.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.115 -119.165 31.445 -118.835 ;
        RECT 31.115 -120.525 31.445 -120.195 ;
        RECT 31.115 -121.885 31.445 -121.555 ;
        RECT 31.115 -123.245 31.445 -122.915 ;
        RECT 31.115 -124.605 31.445 -124.275 ;
        RECT 31.115 -125.965 31.445 -125.635 ;
        RECT 31.115 -127.325 31.445 -126.995 ;
        RECT 31.115 -128.685 31.445 -128.355 ;
        RECT 31.115 -130.045 31.445 -129.715 ;
        RECT 31.115 -131.405 31.445 -131.075 ;
        RECT 31.115 -132.765 31.445 -132.435 ;
        RECT 31.115 -134.125 31.445 -133.795 ;
        RECT 31.115 -135.485 31.445 -135.155 ;
        RECT 31.115 -136.845 31.445 -136.515 ;
        RECT 31.115 -138.205 31.445 -137.875 ;
        RECT 31.115 -139.565 31.445 -139.235 ;
        RECT 31.115 -140.925 31.445 -140.595 ;
        RECT 31.115 -142.285 31.445 -141.955 ;
        RECT 31.115 -143.645 31.445 -143.315 ;
        RECT 31.115 -145.005 31.445 -144.675 ;
        RECT 31.115 -146.365 31.445 -146.035 ;
        RECT 31.115 -147.725 31.445 -147.395 ;
        RECT 31.115 -149.085 31.445 -148.755 ;
        RECT 31.115 -150.445 31.445 -150.115 ;
        RECT 31.115 -151.805 31.445 -151.475 ;
        RECT 31.115 -153.165 31.445 -152.835 ;
        RECT 31.115 -154.525 31.445 -154.195 ;
        RECT 31.115 -155.885 31.445 -155.555 ;
        RECT 31.115 -157.245 31.445 -156.915 ;
        RECT 31.115 -158.605 31.445 -158.275 ;
        RECT 31.115 -159.965 31.445 -159.635 ;
        RECT 31.115 -161.325 31.445 -160.995 ;
        RECT 31.115 -162.685 31.445 -162.355 ;
        RECT 31.115 -164.045 31.445 -163.715 ;
        RECT 31.115 -165.405 31.445 -165.075 ;
        RECT 31.115 -166.765 31.445 -166.435 ;
        RECT 31.115 -168.125 31.445 -167.795 ;
        RECT 31.115 -169.485 31.445 -169.155 ;
        RECT 31.115 -170.845 31.445 -170.515 ;
        RECT 31.115 -172.205 31.445 -171.875 ;
        RECT 31.115 -173.565 31.445 -173.235 ;
        RECT 31.115 -174.925 31.445 -174.595 ;
        RECT 31.115 -176.285 31.445 -175.955 ;
        RECT 31.115 -177.645 31.445 -177.315 ;
        RECT 31.115 -179.005 31.445 -178.675 ;
        RECT 31.115 -180.365 31.445 -180.035 ;
        RECT 31.115 -181.725 31.445 -181.395 ;
        RECT 31.115 -183.085 31.445 -182.755 ;
        RECT 31.115 -184.445 31.445 -184.115 ;
        RECT 31.115 -185.805 31.445 -185.475 ;
        RECT 31.115 -187.165 31.445 -186.835 ;
        RECT 31.115 -188.525 31.445 -188.195 ;
        RECT 31.115 -189.885 31.445 -189.555 ;
        RECT 31.115 -191.245 31.445 -190.915 ;
        RECT 31.115 -192.605 31.445 -192.275 ;
        RECT 31.115 -193.965 31.445 -193.635 ;
        RECT 31.115 -195.325 31.445 -194.995 ;
        RECT 31.115 -196.685 31.445 -196.355 ;
        RECT 31.115 -198.045 31.445 -197.715 ;
        RECT 31.115 -199.405 31.445 -199.075 ;
        RECT 31.115 -200.765 31.445 -200.435 ;
        RECT 31.115 -202.125 31.445 -201.795 ;
        RECT 31.115 -203.485 31.445 -203.155 ;
        RECT 31.115 -204.845 31.445 -204.515 ;
        RECT 31.115 -206.205 31.445 -205.875 ;
        RECT 31.115 -207.565 31.445 -207.235 ;
        RECT 31.115 -208.925 31.445 -208.595 ;
        RECT 31.115 -210.285 31.445 -209.955 ;
        RECT 31.115 -211.645 31.445 -211.315 ;
        RECT 31.115 -213.005 31.445 -212.675 ;
        RECT 31.115 -214.365 31.445 -214.035 ;
        RECT 31.115 -215.725 31.445 -215.395 ;
        RECT 31.115 -217.085 31.445 -216.755 ;
        RECT 31.115 -218.445 31.445 -218.115 ;
        RECT 31.115 -224.09 31.445 -222.96 ;
        RECT 31.12 -224.205 31.44 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.475 132.52 32.805 133.65 ;
        RECT 32.475 128.355 32.805 128.685 ;
        RECT 32.475 126.995 32.805 127.325 ;
        RECT 32.475 125.635 32.805 125.965 ;
        RECT 32.475 124.275 32.805 124.605 ;
        RECT 32.48 123.6 32.8 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.475 -0.845 32.805 -0.515 ;
        RECT 32.475 -2.205 32.805 -1.875 ;
        RECT 32.475 -3.565 32.805 -3.235 ;
        RECT 32.48 -3.565 32.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.475 -119.165 32.805 -118.835 ;
        RECT 32.475 -120.525 32.805 -120.195 ;
        RECT 32.475 -121.885 32.805 -121.555 ;
        RECT 32.475 -123.245 32.805 -122.915 ;
        RECT 32.475 -124.605 32.805 -124.275 ;
        RECT 32.475 -125.965 32.805 -125.635 ;
        RECT 32.475 -127.325 32.805 -126.995 ;
        RECT 32.475 -128.685 32.805 -128.355 ;
        RECT 32.475 -130.045 32.805 -129.715 ;
        RECT 32.475 -131.405 32.805 -131.075 ;
        RECT 32.475 -132.765 32.805 -132.435 ;
        RECT 32.475 -134.125 32.805 -133.795 ;
        RECT 32.475 -135.485 32.805 -135.155 ;
        RECT 32.475 -136.845 32.805 -136.515 ;
        RECT 32.475 -138.205 32.805 -137.875 ;
        RECT 32.475 -139.565 32.805 -139.235 ;
        RECT 32.475 -140.925 32.805 -140.595 ;
        RECT 32.475 -142.285 32.805 -141.955 ;
        RECT 32.475 -143.645 32.805 -143.315 ;
        RECT 32.475 -145.005 32.805 -144.675 ;
        RECT 32.475 -146.365 32.805 -146.035 ;
        RECT 32.475 -147.725 32.805 -147.395 ;
        RECT 32.475 -149.085 32.805 -148.755 ;
        RECT 32.475 -150.445 32.805 -150.115 ;
        RECT 32.475 -151.805 32.805 -151.475 ;
        RECT 32.475 -153.165 32.805 -152.835 ;
        RECT 32.475 -154.525 32.805 -154.195 ;
        RECT 32.475 -155.885 32.805 -155.555 ;
        RECT 32.475 -157.245 32.805 -156.915 ;
        RECT 32.475 -158.605 32.805 -158.275 ;
        RECT 32.475 -159.965 32.805 -159.635 ;
        RECT 32.475 -161.325 32.805 -160.995 ;
        RECT 32.475 -162.685 32.805 -162.355 ;
        RECT 32.475 -164.045 32.805 -163.715 ;
        RECT 32.475 -165.405 32.805 -165.075 ;
        RECT 32.475 -166.765 32.805 -166.435 ;
        RECT 32.475 -168.125 32.805 -167.795 ;
        RECT 32.475 -169.485 32.805 -169.155 ;
        RECT 32.475 -170.845 32.805 -170.515 ;
        RECT 32.475 -172.205 32.805 -171.875 ;
        RECT 32.475 -173.565 32.805 -173.235 ;
        RECT 32.475 -174.925 32.805 -174.595 ;
        RECT 32.475 -176.285 32.805 -175.955 ;
        RECT 32.475 -177.645 32.805 -177.315 ;
        RECT 32.475 -179.005 32.805 -178.675 ;
        RECT 32.475 -180.365 32.805 -180.035 ;
        RECT 32.475 -181.725 32.805 -181.395 ;
        RECT 32.475 -183.085 32.805 -182.755 ;
        RECT 32.475 -184.445 32.805 -184.115 ;
        RECT 32.475 -185.805 32.805 -185.475 ;
        RECT 32.475 -187.165 32.805 -186.835 ;
        RECT 32.475 -188.525 32.805 -188.195 ;
        RECT 32.475 -189.885 32.805 -189.555 ;
        RECT 32.475 -191.245 32.805 -190.915 ;
        RECT 32.475 -192.605 32.805 -192.275 ;
        RECT 32.475 -193.965 32.805 -193.635 ;
        RECT 32.475 -195.325 32.805 -194.995 ;
        RECT 32.475 -196.685 32.805 -196.355 ;
        RECT 32.475 -198.045 32.805 -197.715 ;
        RECT 32.475 -199.405 32.805 -199.075 ;
        RECT 32.475 -200.765 32.805 -200.435 ;
        RECT 32.475 -202.125 32.805 -201.795 ;
        RECT 32.475 -203.485 32.805 -203.155 ;
        RECT 32.475 -204.845 32.805 -204.515 ;
        RECT 32.475 -206.205 32.805 -205.875 ;
        RECT 32.475 -207.565 32.805 -207.235 ;
        RECT 32.475 -208.925 32.805 -208.595 ;
        RECT 32.475 -210.285 32.805 -209.955 ;
        RECT 32.475 -211.645 32.805 -211.315 ;
        RECT 32.475 -213.005 32.805 -212.675 ;
        RECT 32.475 -214.365 32.805 -214.035 ;
        RECT 32.475 -215.725 32.805 -215.395 ;
        RECT 32.475 -217.085 32.805 -216.755 ;
        RECT 32.475 -218.445 32.805 -218.115 ;
        RECT 32.475 -224.09 32.805 -222.96 ;
        RECT 32.48 -224.205 32.8 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.16 -121.535 33.49 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.835 132.52 34.165 133.65 ;
        RECT 33.835 128.355 34.165 128.685 ;
        RECT 33.835 126.995 34.165 127.325 ;
        RECT 33.835 125.635 34.165 125.965 ;
        RECT 33.835 124.275 34.165 124.605 ;
        RECT 33.84 123.6 34.16 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.195 132.52 35.525 133.65 ;
        RECT 35.195 128.355 35.525 128.685 ;
        RECT 35.195 126.995 35.525 127.325 ;
        RECT 35.195 125.635 35.525 125.965 ;
        RECT 35.195 124.275 35.525 124.605 ;
        RECT 35.2 123.6 35.52 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.195 -0.845 35.525 -0.515 ;
        RECT 35.195 -2.205 35.525 -1.875 ;
        RECT 35.195 -3.565 35.525 -3.235 ;
        RECT 35.2 -3.565 35.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.555 132.52 36.885 133.65 ;
        RECT 36.555 128.355 36.885 128.685 ;
        RECT 36.555 126.995 36.885 127.325 ;
        RECT 36.555 125.635 36.885 125.965 ;
        RECT 36.555 124.275 36.885 124.605 ;
        RECT 36.56 123.6 36.88 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.555 -0.845 36.885 -0.515 ;
        RECT 36.555 -2.205 36.885 -1.875 ;
        RECT 36.555 -3.565 36.885 -3.235 ;
        RECT 36.56 -3.565 36.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.915 132.52 38.245 133.65 ;
        RECT 37.915 128.355 38.245 128.685 ;
        RECT 37.915 126.995 38.245 127.325 ;
        RECT 37.915 125.635 38.245 125.965 ;
        RECT 37.915 124.275 38.245 124.605 ;
        RECT 37.92 123.6 38.24 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.915 -0.845 38.245 -0.515 ;
        RECT 37.915 -2.205 38.245 -1.875 ;
        RECT 37.915 -3.565 38.245 -3.235 ;
        RECT 37.92 -3.565 38.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.915 -119.165 38.245 -118.835 ;
        RECT 37.915 -120.525 38.245 -120.195 ;
        RECT 37.915 -121.885 38.245 -121.555 ;
        RECT 37.915 -123.245 38.245 -122.915 ;
        RECT 37.915 -124.605 38.245 -124.275 ;
        RECT 37.915 -125.965 38.245 -125.635 ;
        RECT 37.915 -127.325 38.245 -126.995 ;
        RECT 37.915 -128.685 38.245 -128.355 ;
        RECT 37.915 -130.045 38.245 -129.715 ;
        RECT 37.915 -131.405 38.245 -131.075 ;
        RECT 37.915 -132.765 38.245 -132.435 ;
        RECT 37.915 -134.125 38.245 -133.795 ;
        RECT 37.915 -135.485 38.245 -135.155 ;
        RECT 37.915 -136.845 38.245 -136.515 ;
        RECT 37.915 -138.205 38.245 -137.875 ;
        RECT 37.915 -139.565 38.245 -139.235 ;
        RECT 37.915 -140.925 38.245 -140.595 ;
        RECT 37.915 -142.285 38.245 -141.955 ;
        RECT 37.915 -143.645 38.245 -143.315 ;
        RECT 37.915 -145.005 38.245 -144.675 ;
        RECT 37.915 -146.365 38.245 -146.035 ;
        RECT 37.915 -147.725 38.245 -147.395 ;
        RECT 37.915 -149.085 38.245 -148.755 ;
        RECT 37.915 -150.445 38.245 -150.115 ;
        RECT 37.915 -151.805 38.245 -151.475 ;
        RECT 37.915 -153.165 38.245 -152.835 ;
        RECT 37.915 -154.525 38.245 -154.195 ;
        RECT 37.915 -155.885 38.245 -155.555 ;
        RECT 37.915 -157.245 38.245 -156.915 ;
        RECT 37.915 -158.605 38.245 -158.275 ;
        RECT 37.915 -159.965 38.245 -159.635 ;
        RECT 37.915 -161.325 38.245 -160.995 ;
        RECT 37.915 -162.685 38.245 -162.355 ;
        RECT 37.915 -164.045 38.245 -163.715 ;
        RECT 37.915 -165.405 38.245 -165.075 ;
        RECT 37.915 -166.765 38.245 -166.435 ;
        RECT 37.915 -168.125 38.245 -167.795 ;
        RECT 37.915 -169.485 38.245 -169.155 ;
        RECT 37.915 -170.845 38.245 -170.515 ;
        RECT 37.915 -172.205 38.245 -171.875 ;
        RECT 37.915 -173.565 38.245 -173.235 ;
        RECT 37.915 -174.925 38.245 -174.595 ;
        RECT 37.915 -176.285 38.245 -175.955 ;
        RECT 37.915 -177.645 38.245 -177.315 ;
        RECT 37.915 -179.005 38.245 -178.675 ;
        RECT 37.915 -180.365 38.245 -180.035 ;
        RECT 37.915 -181.725 38.245 -181.395 ;
        RECT 37.915 -183.085 38.245 -182.755 ;
        RECT 37.915 -184.445 38.245 -184.115 ;
        RECT 37.915 -185.805 38.245 -185.475 ;
        RECT 37.915 -187.165 38.245 -186.835 ;
        RECT 37.915 -188.525 38.245 -188.195 ;
        RECT 37.915 -189.885 38.245 -189.555 ;
        RECT 37.915 -191.245 38.245 -190.915 ;
        RECT 37.915 -192.605 38.245 -192.275 ;
        RECT 37.915 -193.965 38.245 -193.635 ;
        RECT 37.915 -195.325 38.245 -194.995 ;
        RECT 37.915 -196.685 38.245 -196.355 ;
        RECT 37.915 -198.045 38.245 -197.715 ;
        RECT 37.915 -199.405 38.245 -199.075 ;
        RECT 37.915 -200.765 38.245 -200.435 ;
        RECT 37.915 -202.125 38.245 -201.795 ;
        RECT 37.915 -203.485 38.245 -203.155 ;
        RECT 37.915 -204.845 38.245 -204.515 ;
        RECT 37.915 -206.205 38.245 -205.875 ;
        RECT 37.915 -207.565 38.245 -207.235 ;
        RECT 37.915 -208.925 38.245 -208.595 ;
        RECT 37.915 -210.285 38.245 -209.955 ;
        RECT 37.915 -211.645 38.245 -211.315 ;
        RECT 37.915 -213.005 38.245 -212.675 ;
        RECT 37.915 -214.365 38.245 -214.035 ;
        RECT 37.915 -215.725 38.245 -215.395 ;
        RECT 37.915 -217.085 38.245 -216.755 ;
        RECT 37.915 -218.445 38.245 -218.115 ;
        RECT 37.915 -224.09 38.245 -222.96 ;
        RECT 37.92 -224.205 38.24 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.26 -121.535 39.59 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.275 132.52 39.605 133.65 ;
        RECT 39.275 128.355 39.605 128.685 ;
        RECT 39.275 126.995 39.605 127.325 ;
        RECT 39.275 125.635 39.605 125.965 ;
        RECT 39.275 124.275 39.605 124.605 ;
        RECT 39.28 123.6 39.6 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.275 -123.245 39.605 -122.915 ;
        RECT 39.275 -124.605 39.605 -124.275 ;
        RECT 39.275 -125.965 39.605 -125.635 ;
        RECT 39.275 -127.325 39.605 -126.995 ;
        RECT 39.275 -128.685 39.605 -128.355 ;
        RECT 39.275 -130.045 39.605 -129.715 ;
        RECT 39.275 -131.405 39.605 -131.075 ;
        RECT 39.275 -132.765 39.605 -132.435 ;
        RECT 39.275 -134.125 39.605 -133.795 ;
        RECT 39.275 -135.485 39.605 -135.155 ;
        RECT 39.275 -136.845 39.605 -136.515 ;
        RECT 39.275 -138.205 39.605 -137.875 ;
        RECT 39.275 -139.565 39.605 -139.235 ;
        RECT 39.275 -140.925 39.605 -140.595 ;
        RECT 39.275 -142.285 39.605 -141.955 ;
        RECT 39.275 -143.645 39.605 -143.315 ;
        RECT 39.275 -145.005 39.605 -144.675 ;
        RECT 39.275 -146.365 39.605 -146.035 ;
        RECT 39.275 -147.725 39.605 -147.395 ;
        RECT 39.275 -149.085 39.605 -148.755 ;
        RECT 39.275 -150.445 39.605 -150.115 ;
        RECT 39.275 -151.805 39.605 -151.475 ;
        RECT 39.275 -153.165 39.605 -152.835 ;
        RECT 39.275 -154.525 39.605 -154.195 ;
        RECT 39.275 -155.885 39.605 -155.555 ;
        RECT 39.275 -157.245 39.605 -156.915 ;
        RECT 39.275 -158.605 39.605 -158.275 ;
        RECT 39.275 -159.965 39.605 -159.635 ;
        RECT 39.275 -161.325 39.605 -160.995 ;
        RECT 39.275 -162.685 39.605 -162.355 ;
        RECT 39.275 -164.045 39.605 -163.715 ;
        RECT 39.275 -165.405 39.605 -165.075 ;
        RECT 39.275 -166.765 39.605 -166.435 ;
        RECT 39.275 -168.125 39.605 -167.795 ;
        RECT 39.275 -169.485 39.605 -169.155 ;
        RECT 39.275 -170.845 39.605 -170.515 ;
        RECT 39.275 -172.205 39.605 -171.875 ;
        RECT 39.275 -173.565 39.605 -173.235 ;
        RECT 39.275 -174.925 39.605 -174.595 ;
        RECT 39.275 -176.285 39.605 -175.955 ;
        RECT 39.275 -177.645 39.605 -177.315 ;
        RECT 39.275 -179.005 39.605 -178.675 ;
        RECT 39.275 -180.365 39.605 -180.035 ;
        RECT 39.275 -181.725 39.605 -181.395 ;
        RECT 39.275 -183.085 39.605 -182.755 ;
        RECT 39.275 -184.445 39.605 -184.115 ;
        RECT 39.275 -185.805 39.605 -185.475 ;
        RECT 39.275 -187.165 39.605 -186.835 ;
        RECT 39.275 -188.525 39.605 -188.195 ;
        RECT 39.275 -189.885 39.605 -189.555 ;
        RECT 39.275 -191.245 39.605 -190.915 ;
        RECT 39.275 -192.605 39.605 -192.275 ;
        RECT 39.275 -193.965 39.605 -193.635 ;
        RECT 39.275 -195.325 39.605 -194.995 ;
        RECT 39.275 -196.685 39.605 -196.355 ;
        RECT 39.275 -198.045 39.605 -197.715 ;
        RECT 39.275 -199.405 39.605 -199.075 ;
        RECT 39.275 -200.765 39.605 -200.435 ;
        RECT 39.275 -202.125 39.605 -201.795 ;
        RECT 39.275 -203.485 39.605 -203.155 ;
        RECT 39.275 -204.845 39.605 -204.515 ;
        RECT 39.275 -206.205 39.605 -205.875 ;
        RECT 39.275 -207.565 39.605 -207.235 ;
        RECT 39.275 -208.925 39.605 -208.595 ;
        RECT 39.275 -210.285 39.605 -209.955 ;
        RECT 39.275 -211.645 39.605 -211.315 ;
        RECT 39.275 -213.005 39.605 -212.675 ;
        RECT 39.275 -214.365 39.605 -214.035 ;
        RECT 39.275 -215.725 39.605 -215.395 ;
        RECT 39.275 -217.085 39.605 -216.755 ;
        RECT 39.275 -218.445 39.605 -218.115 ;
        RECT 39.275 -224.09 39.605 -222.96 ;
        RECT 39.28 -224.205 39.6 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.635 132.52 40.965 133.65 ;
        RECT 40.635 128.355 40.965 128.685 ;
        RECT 40.635 126.995 40.965 127.325 ;
        RECT 40.635 125.635 40.965 125.965 ;
        RECT 40.635 124.275 40.965 124.605 ;
        RECT 40.64 123.6 40.96 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.635 -0.845 40.965 -0.515 ;
        RECT 40.635 -2.205 40.965 -1.875 ;
        RECT 40.635 -3.565 40.965 -3.235 ;
        RECT 40.64 -3.565 40.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.995 132.52 42.325 133.65 ;
        RECT 41.995 128.355 42.325 128.685 ;
        RECT 41.995 126.995 42.325 127.325 ;
        RECT 41.995 125.635 42.325 125.965 ;
        RECT 41.995 124.275 42.325 124.605 ;
        RECT 42 123.6 42.32 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.995 -0.845 42.325 -0.515 ;
        RECT 41.995 -2.205 42.325 -1.875 ;
        RECT 41.995 -3.565 42.325 -3.235 ;
        RECT 42 -3.565 42.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.355 132.52 43.685 133.65 ;
        RECT 43.355 128.355 43.685 128.685 ;
        RECT 43.355 126.995 43.685 127.325 ;
        RECT 43.355 125.635 43.685 125.965 ;
        RECT 43.355 124.275 43.685 124.605 ;
        RECT 43.36 123.6 43.68 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.355 -0.845 43.685 -0.515 ;
        RECT 43.355 -2.205 43.685 -1.875 ;
        RECT 43.355 -3.565 43.685 -3.235 ;
        RECT 43.36 -3.565 43.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.355 -119.165 43.685 -118.835 ;
        RECT 43.355 -120.525 43.685 -120.195 ;
        RECT 43.355 -121.885 43.685 -121.555 ;
        RECT 43.355 -123.245 43.685 -122.915 ;
        RECT 43.355 -124.605 43.685 -124.275 ;
        RECT 43.355 -125.965 43.685 -125.635 ;
        RECT 43.355 -127.325 43.685 -126.995 ;
        RECT 43.355 -128.685 43.685 -128.355 ;
        RECT 43.355 -130.045 43.685 -129.715 ;
        RECT 43.355 -131.405 43.685 -131.075 ;
        RECT 43.355 -132.765 43.685 -132.435 ;
        RECT 43.355 -134.125 43.685 -133.795 ;
        RECT 43.355 -135.485 43.685 -135.155 ;
        RECT 43.355 -136.845 43.685 -136.515 ;
        RECT 43.355 -138.205 43.685 -137.875 ;
        RECT 43.355 -139.565 43.685 -139.235 ;
        RECT 43.355 -140.925 43.685 -140.595 ;
        RECT 43.355 -142.285 43.685 -141.955 ;
        RECT 43.355 -143.645 43.685 -143.315 ;
        RECT 43.355 -145.005 43.685 -144.675 ;
        RECT 43.355 -146.365 43.685 -146.035 ;
        RECT 43.355 -147.725 43.685 -147.395 ;
        RECT 43.355 -149.085 43.685 -148.755 ;
        RECT 43.355 -150.445 43.685 -150.115 ;
        RECT 43.355 -151.805 43.685 -151.475 ;
        RECT 43.355 -153.165 43.685 -152.835 ;
        RECT 43.355 -154.525 43.685 -154.195 ;
        RECT 43.355 -155.885 43.685 -155.555 ;
        RECT 43.355 -157.245 43.685 -156.915 ;
        RECT 43.355 -158.605 43.685 -158.275 ;
        RECT 43.355 -159.965 43.685 -159.635 ;
        RECT 43.355 -161.325 43.685 -160.995 ;
        RECT 43.355 -162.685 43.685 -162.355 ;
        RECT 43.355 -164.045 43.685 -163.715 ;
        RECT 43.355 -165.405 43.685 -165.075 ;
        RECT 43.355 -166.765 43.685 -166.435 ;
        RECT 43.355 -168.125 43.685 -167.795 ;
        RECT 43.355 -169.485 43.685 -169.155 ;
        RECT 43.355 -170.845 43.685 -170.515 ;
        RECT 43.355 -172.205 43.685 -171.875 ;
        RECT 43.355 -173.565 43.685 -173.235 ;
        RECT 43.355 -174.925 43.685 -174.595 ;
        RECT 43.355 -176.285 43.685 -175.955 ;
        RECT 43.355 -177.645 43.685 -177.315 ;
        RECT 43.355 -179.005 43.685 -178.675 ;
        RECT 43.355 -180.365 43.685 -180.035 ;
        RECT 43.355 -181.725 43.685 -181.395 ;
        RECT 43.355 -183.085 43.685 -182.755 ;
        RECT 43.355 -184.445 43.685 -184.115 ;
        RECT 43.355 -185.805 43.685 -185.475 ;
        RECT 43.355 -187.165 43.685 -186.835 ;
        RECT 43.355 -188.525 43.685 -188.195 ;
        RECT 43.355 -189.885 43.685 -189.555 ;
        RECT 43.355 -191.245 43.685 -190.915 ;
        RECT 43.355 -192.605 43.685 -192.275 ;
        RECT 43.355 -193.965 43.685 -193.635 ;
        RECT 43.355 -195.325 43.685 -194.995 ;
        RECT 43.355 -196.685 43.685 -196.355 ;
        RECT 43.355 -198.045 43.685 -197.715 ;
        RECT 43.355 -199.405 43.685 -199.075 ;
        RECT 43.355 -200.765 43.685 -200.435 ;
        RECT 43.355 -202.125 43.685 -201.795 ;
        RECT 43.355 -203.485 43.685 -203.155 ;
        RECT 43.355 -204.845 43.685 -204.515 ;
        RECT 43.355 -206.205 43.685 -205.875 ;
        RECT 43.355 -207.565 43.685 -207.235 ;
        RECT 43.355 -208.925 43.685 -208.595 ;
        RECT 43.355 -210.285 43.685 -209.955 ;
        RECT 43.355 -211.645 43.685 -211.315 ;
        RECT 43.355 -213.005 43.685 -212.675 ;
        RECT 43.355 -214.365 43.685 -214.035 ;
        RECT 43.355 -215.725 43.685 -215.395 ;
        RECT 43.355 -217.085 43.685 -216.755 ;
        RECT 43.355 -218.445 43.685 -218.115 ;
        RECT 43.355 -224.09 43.685 -222.96 ;
        RECT 43.36 -224.205 43.68 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.715 132.52 45.045 133.65 ;
        RECT 44.715 128.355 45.045 128.685 ;
        RECT 44.715 126.995 45.045 127.325 ;
        RECT 44.715 125.635 45.045 125.965 ;
        RECT 44.715 124.275 45.045 124.605 ;
        RECT 44.72 123.6 45.04 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.715 -217.085 45.045 -216.755 ;
        RECT 44.715 -218.445 45.045 -218.115 ;
        RECT 44.715 -224.09 45.045 -222.96 ;
        RECT 44.72 -224.205 45.04 -122.24 ;
        RECT 44.715 -123.245 45.045 -122.915 ;
        RECT 44.715 -124.605 45.045 -124.275 ;
        RECT 44.715 -125.965 45.045 -125.635 ;
        RECT 44.715 -127.325 45.045 -126.995 ;
        RECT 44.715 -128.685 45.045 -128.355 ;
        RECT 44.715 -130.045 45.045 -129.715 ;
        RECT 44.715 -131.405 45.045 -131.075 ;
        RECT 44.715 -132.765 45.045 -132.435 ;
        RECT 44.715 -134.125 45.045 -133.795 ;
        RECT 44.715 -135.485 45.045 -135.155 ;
        RECT 44.715 -136.845 45.045 -136.515 ;
        RECT 44.715 -138.205 45.045 -137.875 ;
        RECT 44.715 -139.565 45.045 -139.235 ;
        RECT 44.715 -140.925 45.045 -140.595 ;
        RECT 44.715 -142.285 45.045 -141.955 ;
        RECT 44.715 -143.645 45.045 -143.315 ;
        RECT 44.715 -145.005 45.045 -144.675 ;
        RECT 44.715 -146.365 45.045 -146.035 ;
        RECT 44.715 -147.725 45.045 -147.395 ;
        RECT 44.715 -149.085 45.045 -148.755 ;
        RECT 44.715 -150.445 45.045 -150.115 ;
        RECT 44.715 -151.805 45.045 -151.475 ;
        RECT 44.715 -153.165 45.045 -152.835 ;
        RECT 44.715 -154.525 45.045 -154.195 ;
        RECT 44.715 -155.885 45.045 -155.555 ;
        RECT 44.715 -157.245 45.045 -156.915 ;
        RECT 44.715 -158.605 45.045 -158.275 ;
        RECT 44.715 -159.965 45.045 -159.635 ;
        RECT 44.715 -161.325 45.045 -160.995 ;
        RECT 44.715 -162.685 45.045 -162.355 ;
        RECT 44.715 -164.045 45.045 -163.715 ;
        RECT 44.715 -165.405 45.045 -165.075 ;
        RECT 44.715 -166.765 45.045 -166.435 ;
        RECT 44.715 -168.125 45.045 -167.795 ;
        RECT 44.715 -169.485 45.045 -169.155 ;
        RECT 44.715 -170.845 45.045 -170.515 ;
        RECT 44.715 -172.205 45.045 -171.875 ;
        RECT 44.715 -173.565 45.045 -173.235 ;
        RECT 44.715 -174.925 45.045 -174.595 ;
        RECT 44.715 -176.285 45.045 -175.955 ;
        RECT 44.715 -177.645 45.045 -177.315 ;
        RECT 44.715 -179.005 45.045 -178.675 ;
        RECT 44.715 -180.365 45.045 -180.035 ;
        RECT 44.715 -181.725 45.045 -181.395 ;
        RECT 44.715 -183.085 45.045 -182.755 ;
        RECT 44.715 -184.445 45.045 -184.115 ;
        RECT 44.715 -185.805 45.045 -185.475 ;
        RECT 44.715 -187.165 45.045 -186.835 ;
        RECT 44.715 -188.525 45.045 -188.195 ;
        RECT 44.715 -189.885 45.045 -189.555 ;
        RECT 44.715 -191.245 45.045 -190.915 ;
        RECT 44.715 -192.605 45.045 -192.275 ;
        RECT 44.715 -193.965 45.045 -193.635 ;
        RECT 44.715 -195.325 45.045 -194.995 ;
        RECT 44.715 -196.685 45.045 -196.355 ;
        RECT 44.715 -198.045 45.045 -197.715 ;
        RECT 44.715 -199.405 45.045 -199.075 ;
        RECT 44.715 -200.765 45.045 -200.435 ;
        RECT 44.715 -202.125 45.045 -201.795 ;
        RECT 44.715 -203.485 45.045 -203.155 ;
        RECT 44.715 -204.845 45.045 -204.515 ;
        RECT 44.715 -206.205 45.045 -205.875 ;
        RECT 44.715 -207.565 45.045 -207.235 ;
        RECT 44.715 -208.925 45.045 -208.595 ;
        RECT 44.715 -210.285 45.045 -209.955 ;
        RECT 44.715 -211.645 45.045 -211.315 ;
        RECT 44.715 -213.005 45.045 -212.675 ;
        RECT 44.715 -214.365 45.045 -214.035 ;
        RECT 44.715 -215.725 45.045 -215.395 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.525 132.52 -1.195 133.65 ;
        RECT -1.525 128.355 -1.195 128.685 ;
        RECT -1.525 126.995 -1.195 127.325 ;
        RECT -1.525 125.635 -1.195 125.965 ;
        RECT -1.525 124.275 -1.195 124.605 ;
        RECT -1.525 121.41 -1.195 121.74 ;
        RECT -1.525 119.235 -1.195 119.565 ;
        RECT -1.525 117.655 -1.195 117.985 ;
        RECT -1.525 116.805 -1.195 117.135 ;
        RECT -1.525 114.495 -1.195 114.825 ;
        RECT -1.525 113.645 -1.195 113.975 ;
        RECT -1.525 111.335 -1.195 111.665 ;
        RECT -1.525 110.485 -1.195 110.815 ;
        RECT -1.525 108.175 -1.195 108.505 ;
        RECT -1.525 107.325 -1.195 107.655 ;
        RECT -1.525 105.015 -1.195 105.345 ;
        RECT -1.525 103.435 -1.195 103.765 ;
        RECT -1.525 102.585 -1.195 102.915 ;
        RECT -1.525 100.275 -1.195 100.605 ;
        RECT -1.525 99.425 -1.195 99.755 ;
        RECT -1.525 97.115 -1.195 97.445 ;
        RECT -1.525 96.265 -1.195 96.595 ;
        RECT -1.525 93.955 -1.195 94.285 ;
        RECT -1.525 93.105 -1.195 93.435 ;
        RECT -1.525 90.795 -1.195 91.125 ;
        RECT -1.525 89.215 -1.195 89.545 ;
        RECT -1.525 88.365 -1.195 88.695 ;
        RECT -1.525 86.055 -1.195 86.385 ;
        RECT -1.525 85.205 -1.195 85.535 ;
        RECT -1.525 82.895 -1.195 83.225 ;
        RECT -1.525 82.045 -1.195 82.375 ;
        RECT -1.525 79.735 -1.195 80.065 ;
        RECT -1.525 78.885 -1.195 79.215 ;
        RECT -1.525 76.575 -1.195 76.905 ;
        RECT -1.525 74.995 -1.195 75.325 ;
        RECT -1.525 74.145 -1.195 74.475 ;
        RECT -1.525 71.835 -1.195 72.165 ;
        RECT -1.525 70.985 -1.195 71.315 ;
        RECT -1.525 68.675 -1.195 69.005 ;
        RECT -1.525 67.825 -1.195 68.155 ;
        RECT -1.525 65.515 -1.195 65.845 ;
        RECT -1.525 64.665 -1.195 64.995 ;
        RECT -1.525 62.355 -1.195 62.685 ;
        RECT -1.525 60.775 -1.195 61.105 ;
        RECT -1.525 59.925 -1.195 60.255 ;
        RECT -1.525 57.615 -1.195 57.945 ;
        RECT -1.525 56.765 -1.195 57.095 ;
        RECT -1.525 54.455 -1.195 54.785 ;
        RECT -1.525 53.605 -1.195 53.935 ;
        RECT -1.525 51.295 -1.195 51.625 ;
        RECT -1.525 50.445 -1.195 50.775 ;
        RECT -1.525 48.135 -1.195 48.465 ;
        RECT -1.525 46.555 -1.195 46.885 ;
        RECT -1.525 45.705 -1.195 46.035 ;
        RECT -1.525 43.395 -1.195 43.725 ;
        RECT -1.525 42.545 -1.195 42.875 ;
        RECT -1.525 40.235 -1.195 40.565 ;
        RECT -1.525 39.385 -1.195 39.715 ;
        RECT -1.525 37.075 -1.195 37.405 ;
        RECT -1.525 36.225 -1.195 36.555 ;
        RECT -1.525 33.915 -1.195 34.245 ;
        RECT -1.525 32.335 -1.195 32.665 ;
        RECT -1.525 31.485 -1.195 31.815 ;
        RECT -1.525 29.175 -1.195 29.505 ;
        RECT -1.525 28.325 -1.195 28.655 ;
        RECT -1.525 26.015 -1.195 26.345 ;
        RECT -1.525 25.165 -1.195 25.495 ;
        RECT -1.525 22.855 -1.195 23.185 ;
        RECT -1.525 22.005 -1.195 22.335 ;
        RECT -1.525 19.695 -1.195 20.025 ;
        RECT -1.525 18.115 -1.195 18.445 ;
        RECT -1.525 17.265 -1.195 17.595 ;
        RECT -1.525 14.955 -1.195 15.285 ;
        RECT -1.525 14.105 -1.195 14.435 ;
        RECT -1.525 11.795 -1.195 12.125 ;
        RECT -1.525 10.945 -1.195 11.275 ;
        RECT -1.525 8.635 -1.195 8.965 ;
        RECT -1.525 7.785 -1.195 8.115 ;
        RECT -1.525 5.475 -1.195 5.805 ;
        RECT -1.525 3.895 -1.195 4.225 ;
        RECT -1.525 3.045 -1.195 3.375 ;
        RECT -1.525 0.87 -1.195 1.2 ;
        RECT -1.525 -0.845 -1.195 -0.515 ;
        RECT -1.525 -2.205 -1.195 -1.875 ;
        RECT -1.525 -3.565 -1.195 -3.235 ;
        RECT -1.525 -4.925 -1.195 -4.595 ;
        RECT -1.525 -6.285 -1.195 -5.955 ;
        RECT -1.525 -7.645 -1.195 -7.315 ;
        RECT -1.525 -9.005 -1.195 -8.675 ;
        RECT -1.525 -10.365 -1.195 -10.035 ;
        RECT -1.525 -11.725 -1.195 -11.395 ;
        RECT -1.525 -13.085 -1.195 -12.755 ;
        RECT -1.525 -14.445 -1.195 -14.115 ;
        RECT -1.525 -15.805 -1.195 -15.475 ;
        RECT -1.525 -17.165 -1.195 -16.835 ;
        RECT -1.525 -18.525 -1.195 -18.195 ;
        RECT -1.525 -21.245 -1.195 -20.915 ;
        RECT -1.525 -22.605 -1.195 -22.275 ;
        RECT -1.525 -23.965 -1.195 -23.635 ;
        RECT -1.525 -25.325 -1.195 -24.995 ;
        RECT -1.525 -26.685 -1.195 -26.355 ;
        RECT -1.525 -28.045 -1.195 -27.715 ;
        RECT -1.525 -29.405 -1.195 -29.075 ;
        RECT -1.525 -30.765 -1.195 -30.435 ;
        RECT -1.525 -32.125 -1.195 -31.795 ;
        RECT -1.525 -33.485 -1.195 -33.155 ;
        RECT -1.525 -34.845 -1.195 -34.515 ;
        RECT -1.525 -36.205 -1.195 -35.875 ;
        RECT -1.525 -37.565 -1.195 -37.235 ;
        RECT -1.525 -38.925 -1.195 -38.595 ;
        RECT -1.525 -40.285 -1.195 -39.955 ;
        RECT -1.525 -41.645 -1.195 -41.315 ;
        RECT -1.525 -43.005 -1.195 -42.675 ;
        RECT -1.525 -44.365 -1.195 -44.035 ;
        RECT -1.525 -45.725 -1.195 -45.395 ;
        RECT -1.525 -47.085 -1.195 -46.755 ;
        RECT -1.525 -48.445 -1.195 -48.115 ;
        RECT -1.525 -49.805 -1.195 -49.475 ;
        RECT -1.525 -51.165 -1.195 -50.835 ;
        RECT -1.525 -52.525 -1.195 -52.195 ;
        RECT -1.525 -53.885 -1.195 -53.555 ;
        RECT -1.525 -55.245 -1.195 -54.915 ;
        RECT -1.525 -56.605 -1.195 -56.275 ;
        RECT -1.525 -57.965 -1.195 -57.635 ;
        RECT -1.525 -59.325 -1.195 -58.995 ;
        RECT -1.525 -62.045 -1.195 -61.715 ;
        RECT -1.525 -66.125 -1.195 -65.795 ;
        RECT -1.525 -68.845 -1.195 -68.515 ;
        RECT -1.525 -70.205 -1.195 -69.875 ;
        RECT -1.525 -71.565 -1.195 -71.235 ;
        RECT -1.525 -72.925 -1.195 -72.595 ;
        RECT -1.525 -74.285 -1.195 -73.955 ;
        RECT -1.525 -75.645 -1.195 -75.315 ;
        RECT -1.525 -77.005 -1.195 -76.675 ;
        RECT -1.525 -78.365 -1.195 -78.035 ;
        RECT -1.525 -79.725 -1.195 -79.395 ;
        RECT -1.525 -81.085 -1.195 -80.755 ;
        RECT -1.525 -82.445 -1.195 -82.115 ;
        RECT -1.525 -83.805 -1.195 -83.475 ;
        RECT -1.525 -85.165 -1.195 -84.835 ;
        RECT -1.525 -86.525 -1.195 -86.195 ;
        RECT -1.525 -87.885 -1.195 -87.555 ;
        RECT -1.525 -89.245 -1.195 -88.915 ;
        RECT -1.525 -90.605 -1.195 -90.275 ;
        RECT -1.525 -91.965 -1.195 -91.635 ;
        RECT -1.525 -93.325 -1.195 -92.995 ;
        RECT -1.525 -94.685 -1.195 -94.355 ;
        RECT -1.525 -96.045 -1.195 -95.715 ;
        RECT -1.525 -97.405 -1.195 -97.075 ;
        RECT -1.525 -98.765 -1.195 -98.435 ;
        RECT -1.525 -100.125 -1.195 -99.795 ;
        RECT -1.525 -101.485 -1.195 -101.155 ;
        RECT -1.525 -102.845 -1.195 -102.515 ;
        RECT -1.525 -104.205 -1.195 -103.875 ;
        RECT -1.525 -105.565 -1.195 -105.235 ;
        RECT -1.525 -106.925 -1.195 -106.595 ;
        RECT -1.525 -108.285 -1.195 -107.955 ;
        RECT -1.525 -109.645 -1.195 -109.315 ;
        RECT -1.525 -111.005 -1.195 -110.675 ;
        RECT -1.525 -115.085 -1.195 -114.755 ;
        RECT -1.525 -116.445 -1.195 -116.115 ;
        RECT -1.525 -117.805 -1.195 -117.475 ;
        RECT -1.525 -119.165 -1.195 -118.835 ;
        RECT -1.525 -120.525 -1.195 -120.195 ;
        RECT -1.525 -121.885 -1.195 -121.555 ;
        RECT -1.525 -123.245 -1.195 -122.915 ;
        RECT -1.525 -124.605 -1.195 -124.275 ;
        RECT -1.525 -125.965 -1.195 -125.635 ;
        RECT -1.525 -127.325 -1.195 -126.995 ;
        RECT -1.525 -128.685 -1.195 -128.355 ;
        RECT -1.525 -130.045 -1.195 -129.715 ;
        RECT -1.525 -131.405 -1.195 -131.075 ;
        RECT -1.525 -132.765 -1.195 -132.435 ;
        RECT -1.525 -134.125 -1.195 -133.795 ;
        RECT -1.525 -135.485 -1.195 -135.155 ;
        RECT -1.525 -136.845 -1.195 -136.515 ;
        RECT -1.525 -138.205 -1.195 -137.875 ;
        RECT -1.525 -139.565 -1.195 -139.235 ;
        RECT -1.525 -140.925 -1.195 -140.595 ;
        RECT -1.525 -142.285 -1.195 -141.955 ;
        RECT -1.525 -143.645 -1.195 -143.315 ;
        RECT -1.525 -145.005 -1.195 -144.675 ;
        RECT -1.525 -146.365 -1.195 -146.035 ;
        RECT -1.525 -147.725 -1.195 -147.395 ;
        RECT -1.525 -149.085 -1.195 -148.755 ;
        RECT -1.525 -150.445 -1.195 -150.115 ;
        RECT -1.525 -151.805 -1.195 -151.475 ;
        RECT -1.525 -153.165 -1.195 -152.835 ;
        RECT -1.525 -154.525 -1.195 -154.195 ;
        RECT -1.525 -155.885 -1.195 -155.555 ;
        RECT -1.525 -157.245 -1.195 -156.915 ;
        RECT -1.525 -158.605 -1.195 -158.275 ;
        RECT -1.525 -159.965 -1.195 -159.635 ;
        RECT -1.525 -161.325 -1.195 -160.995 ;
        RECT -1.525 -162.685 -1.195 -162.355 ;
        RECT -1.525 -164.045 -1.195 -163.715 ;
        RECT -1.525 -165.405 -1.195 -165.075 ;
        RECT -1.525 -166.765 -1.195 -166.435 ;
        RECT -1.525 -168.125 -1.195 -167.795 ;
        RECT -1.525 -169.485 -1.195 -169.155 ;
        RECT -1.525 -170.845 -1.195 -170.515 ;
        RECT -1.525 -172.205 -1.195 -171.875 ;
        RECT -1.525 -173.565 -1.195 -173.235 ;
        RECT -1.525 -174.925 -1.195 -174.595 ;
        RECT -1.525 -176.285 -1.195 -175.955 ;
        RECT -1.525 -177.645 -1.195 -177.315 ;
        RECT -1.525 -179.005 -1.195 -178.675 ;
        RECT -1.525 -180.365 -1.195 -180.035 ;
        RECT -1.525 -181.725 -1.195 -181.395 ;
        RECT -1.525 -183.085 -1.195 -182.755 ;
        RECT -1.525 -184.445 -1.195 -184.115 ;
        RECT -1.525 -185.805 -1.195 -185.475 ;
        RECT -1.525 -187.165 -1.195 -186.835 ;
        RECT -1.525 -188.525 -1.195 -188.195 ;
        RECT -1.525 -189.885 -1.195 -189.555 ;
        RECT -1.525 -191.245 -1.195 -190.915 ;
        RECT -1.525 -192.605 -1.195 -192.275 ;
        RECT -1.525 -193.965 -1.195 -193.635 ;
        RECT -1.525 -195.325 -1.195 -194.995 ;
        RECT -1.525 -196.685 -1.195 -196.355 ;
        RECT -1.525 -198.045 -1.195 -197.715 ;
        RECT -1.525 -199.405 -1.195 -199.075 ;
        RECT -1.525 -200.765 -1.195 -200.435 ;
        RECT -1.525 -202.125 -1.195 -201.795 ;
        RECT -1.525 -203.485 -1.195 -203.155 ;
        RECT -1.525 -204.845 -1.195 -204.515 ;
        RECT -1.525 -206.205 -1.195 -205.875 ;
        RECT -1.525 -207.565 -1.195 -207.235 ;
        RECT -1.525 -208.925 -1.195 -208.595 ;
        RECT -1.525 -210.285 -1.195 -209.955 ;
        RECT -1.525 -211.645 -1.195 -211.315 ;
        RECT -1.525 -213.005 -1.195 -212.675 ;
        RECT -1.525 -214.365 -1.195 -214.035 ;
        RECT -1.525 -215.725 -1.195 -215.395 ;
        RECT -1.525 -217.085 -1.195 -216.755 ;
        RECT -1.525 -218.445 -1.195 -218.115 ;
        RECT -1.525 -224.09 -1.195 -222.96 ;
        RECT -1.52 -224.205 -1.2 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.165 132.52 0.165 133.65 ;
        RECT -0.165 128.355 0.165 128.685 ;
        RECT -0.165 126.995 0.165 127.325 ;
        RECT -0.165 125.635 0.165 125.965 ;
        RECT -0.165 124.275 0.165 124.605 ;
        RECT -0.16 123.6 0.16 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.165 -0.845 0.165 -0.515 ;
        RECT -0.165 -2.205 0.165 -1.875 ;
        RECT -0.165 -3.565 0.165 -3.235 ;
        RECT -0.16 -3.565 0.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.165 -119.165 0.165 -118.835 ;
        RECT -0.165 -120.525 0.165 -120.195 ;
        RECT -0.165 -121.885 0.165 -121.555 ;
        RECT -0.165 -123.245 0.165 -122.915 ;
        RECT -0.165 -124.605 0.165 -124.275 ;
        RECT -0.165 -125.965 0.165 -125.635 ;
        RECT -0.165 -127.325 0.165 -126.995 ;
        RECT -0.165 -128.685 0.165 -128.355 ;
        RECT -0.165 -130.045 0.165 -129.715 ;
        RECT -0.165 -131.405 0.165 -131.075 ;
        RECT -0.165 -132.765 0.165 -132.435 ;
        RECT -0.165 -134.125 0.165 -133.795 ;
        RECT -0.165 -135.485 0.165 -135.155 ;
        RECT -0.165 -136.845 0.165 -136.515 ;
        RECT -0.165 -138.205 0.165 -137.875 ;
        RECT -0.165 -139.565 0.165 -139.235 ;
        RECT -0.165 -140.925 0.165 -140.595 ;
        RECT -0.165 -142.285 0.165 -141.955 ;
        RECT -0.165 -143.645 0.165 -143.315 ;
        RECT -0.165 -145.005 0.165 -144.675 ;
        RECT -0.165 -146.365 0.165 -146.035 ;
        RECT -0.165 -147.725 0.165 -147.395 ;
        RECT -0.165 -149.085 0.165 -148.755 ;
        RECT -0.165 -150.445 0.165 -150.115 ;
        RECT -0.165 -151.805 0.165 -151.475 ;
        RECT -0.165 -153.165 0.165 -152.835 ;
        RECT -0.165 -154.525 0.165 -154.195 ;
        RECT -0.165 -155.885 0.165 -155.555 ;
        RECT -0.165 -157.245 0.165 -156.915 ;
        RECT -0.165 -158.605 0.165 -158.275 ;
        RECT -0.165 -159.965 0.165 -159.635 ;
        RECT -0.165 -161.325 0.165 -160.995 ;
        RECT -0.165 -162.685 0.165 -162.355 ;
        RECT -0.165 -164.045 0.165 -163.715 ;
        RECT -0.165 -165.405 0.165 -165.075 ;
        RECT -0.165 -166.765 0.165 -166.435 ;
        RECT -0.165 -168.125 0.165 -167.795 ;
        RECT -0.165 -169.485 0.165 -169.155 ;
        RECT -0.165 -170.845 0.165 -170.515 ;
        RECT -0.165 -172.205 0.165 -171.875 ;
        RECT -0.165 -173.565 0.165 -173.235 ;
        RECT -0.165 -174.925 0.165 -174.595 ;
        RECT -0.165 -176.285 0.165 -175.955 ;
        RECT -0.165 -177.645 0.165 -177.315 ;
        RECT -0.165 -179.005 0.165 -178.675 ;
        RECT -0.165 -180.365 0.165 -180.035 ;
        RECT -0.165 -181.725 0.165 -181.395 ;
        RECT -0.165 -183.085 0.165 -182.755 ;
        RECT -0.165 -184.445 0.165 -184.115 ;
        RECT -0.165 -185.805 0.165 -185.475 ;
        RECT -0.165 -187.165 0.165 -186.835 ;
        RECT -0.165 -188.525 0.165 -188.195 ;
        RECT -0.165 -189.885 0.165 -189.555 ;
        RECT -0.165 -191.245 0.165 -190.915 ;
        RECT -0.165 -192.605 0.165 -192.275 ;
        RECT -0.165 -193.965 0.165 -193.635 ;
        RECT -0.165 -195.325 0.165 -194.995 ;
        RECT -0.165 -196.685 0.165 -196.355 ;
        RECT -0.165 -198.045 0.165 -197.715 ;
        RECT -0.165 -199.405 0.165 -199.075 ;
        RECT -0.165 -200.765 0.165 -200.435 ;
        RECT -0.165 -202.125 0.165 -201.795 ;
        RECT -0.165 -203.485 0.165 -203.155 ;
        RECT -0.165 -204.845 0.165 -204.515 ;
        RECT -0.165 -206.205 0.165 -205.875 ;
        RECT -0.165 -207.565 0.165 -207.235 ;
        RECT -0.165 -208.925 0.165 -208.595 ;
        RECT -0.165 -210.285 0.165 -209.955 ;
        RECT -0.165 -211.645 0.165 -211.315 ;
        RECT -0.165 -213.005 0.165 -212.675 ;
        RECT -0.165 -214.365 0.165 -214.035 ;
        RECT -0.165 -215.725 0.165 -215.395 ;
        RECT -0.165 -217.085 0.165 -216.755 ;
        RECT -0.165 -218.445 0.165 -218.115 ;
        RECT -0.165 -224.09 0.165 -222.96 ;
        RECT -0.16 -224.205 0.16 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.195 132.52 1.525 133.65 ;
        RECT 1.195 128.355 1.525 128.685 ;
        RECT 1.195 126.995 1.525 127.325 ;
        RECT 1.195 125.635 1.525 125.965 ;
        RECT 1.195 124.275 1.525 124.605 ;
        RECT 1.2 123.6 1.52 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.195 -0.845 1.525 -0.515 ;
        RECT 1.195 -2.205 1.525 -1.875 ;
        RECT 1.195 -3.565 1.525 -3.235 ;
        RECT 1.2 -3.565 1.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.195 -119.165 1.525 -118.835 ;
        RECT 1.195 -120.525 1.525 -120.195 ;
        RECT 1.195 -121.885 1.525 -121.555 ;
        RECT 1.195 -123.245 1.525 -122.915 ;
        RECT 1.195 -124.605 1.525 -124.275 ;
        RECT 1.195 -125.965 1.525 -125.635 ;
        RECT 1.195 -127.325 1.525 -126.995 ;
        RECT 1.195 -128.685 1.525 -128.355 ;
        RECT 1.195 -130.045 1.525 -129.715 ;
        RECT 1.195 -131.405 1.525 -131.075 ;
        RECT 1.195 -132.765 1.525 -132.435 ;
        RECT 1.195 -134.125 1.525 -133.795 ;
        RECT 1.195 -135.485 1.525 -135.155 ;
        RECT 1.195 -136.845 1.525 -136.515 ;
        RECT 1.195 -138.205 1.525 -137.875 ;
        RECT 1.195 -139.565 1.525 -139.235 ;
        RECT 1.195 -140.925 1.525 -140.595 ;
        RECT 1.195 -142.285 1.525 -141.955 ;
        RECT 1.195 -143.645 1.525 -143.315 ;
        RECT 1.195 -145.005 1.525 -144.675 ;
        RECT 1.195 -146.365 1.525 -146.035 ;
        RECT 1.195 -147.725 1.525 -147.395 ;
        RECT 1.195 -149.085 1.525 -148.755 ;
        RECT 1.195 -150.445 1.525 -150.115 ;
        RECT 1.195 -151.805 1.525 -151.475 ;
        RECT 1.195 -153.165 1.525 -152.835 ;
        RECT 1.195 -154.525 1.525 -154.195 ;
        RECT 1.195 -155.885 1.525 -155.555 ;
        RECT 1.195 -157.245 1.525 -156.915 ;
        RECT 1.195 -158.605 1.525 -158.275 ;
        RECT 1.195 -159.965 1.525 -159.635 ;
        RECT 1.195 -161.325 1.525 -160.995 ;
        RECT 1.195 -162.685 1.525 -162.355 ;
        RECT 1.195 -164.045 1.525 -163.715 ;
        RECT 1.195 -165.405 1.525 -165.075 ;
        RECT 1.195 -166.765 1.525 -166.435 ;
        RECT 1.195 -168.125 1.525 -167.795 ;
        RECT 1.195 -169.485 1.525 -169.155 ;
        RECT 1.195 -170.845 1.525 -170.515 ;
        RECT 1.195 -172.205 1.525 -171.875 ;
        RECT 1.195 -173.565 1.525 -173.235 ;
        RECT 1.195 -174.925 1.525 -174.595 ;
        RECT 1.195 -176.285 1.525 -175.955 ;
        RECT 1.195 -177.645 1.525 -177.315 ;
        RECT 1.195 -179.005 1.525 -178.675 ;
        RECT 1.195 -180.365 1.525 -180.035 ;
        RECT 1.195 -181.725 1.525 -181.395 ;
        RECT 1.195 -183.085 1.525 -182.755 ;
        RECT 1.195 -184.445 1.525 -184.115 ;
        RECT 1.195 -185.805 1.525 -185.475 ;
        RECT 1.195 -187.165 1.525 -186.835 ;
        RECT 1.195 -188.525 1.525 -188.195 ;
        RECT 1.195 -189.885 1.525 -189.555 ;
        RECT 1.195 -191.245 1.525 -190.915 ;
        RECT 1.195 -192.605 1.525 -192.275 ;
        RECT 1.195 -193.965 1.525 -193.635 ;
        RECT 1.195 -195.325 1.525 -194.995 ;
        RECT 1.195 -196.685 1.525 -196.355 ;
        RECT 1.195 -198.045 1.525 -197.715 ;
        RECT 1.195 -199.405 1.525 -199.075 ;
        RECT 1.195 -200.765 1.525 -200.435 ;
        RECT 1.195 -202.125 1.525 -201.795 ;
        RECT 1.195 -203.485 1.525 -203.155 ;
        RECT 1.195 -204.845 1.525 -204.515 ;
        RECT 1.195 -206.205 1.525 -205.875 ;
        RECT 1.195 -207.565 1.525 -207.235 ;
        RECT 1.195 -208.925 1.525 -208.595 ;
        RECT 1.195 -210.285 1.525 -209.955 ;
        RECT 1.195 -211.645 1.525 -211.315 ;
        RECT 1.195 -213.005 1.525 -212.675 ;
        RECT 1.195 -214.365 1.525 -214.035 ;
        RECT 1.195 -215.725 1.525 -215.395 ;
        RECT 1.195 -217.085 1.525 -216.755 ;
        RECT 1.195 -218.445 1.525 -218.115 ;
        RECT 1.195 -224.09 1.525 -222.96 ;
        RECT 1.2 -224.205 1.52 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 132.52 2.885 133.65 ;
        RECT 2.555 128.355 2.885 128.685 ;
        RECT 2.555 126.995 2.885 127.325 ;
        RECT 2.555 125.635 2.885 125.965 ;
        RECT 2.555 124.275 2.885 124.605 ;
        RECT 2.56 123.6 2.88 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 -123.245 2.885 -122.915 ;
        RECT 2.555 -124.605 2.885 -124.275 ;
        RECT 2.555 -125.965 2.885 -125.635 ;
        RECT 2.555 -127.325 2.885 -126.995 ;
        RECT 2.555 -128.685 2.885 -128.355 ;
        RECT 2.555 -130.045 2.885 -129.715 ;
        RECT 2.555 -131.405 2.885 -131.075 ;
        RECT 2.555 -132.765 2.885 -132.435 ;
        RECT 2.555 -134.125 2.885 -133.795 ;
        RECT 2.555 -135.485 2.885 -135.155 ;
        RECT 2.555 -136.845 2.885 -136.515 ;
        RECT 2.555 -138.205 2.885 -137.875 ;
        RECT 2.555 -139.565 2.885 -139.235 ;
        RECT 2.555 -140.925 2.885 -140.595 ;
        RECT 2.555 -142.285 2.885 -141.955 ;
        RECT 2.555 -143.645 2.885 -143.315 ;
        RECT 2.555 -145.005 2.885 -144.675 ;
        RECT 2.555 -146.365 2.885 -146.035 ;
        RECT 2.555 -147.725 2.885 -147.395 ;
        RECT 2.555 -149.085 2.885 -148.755 ;
        RECT 2.555 -150.445 2.885 -150.115 ;
        RECT 2.555 -151.805 2.885 -151.475 ;
        RECT 2.555 -153.165 2.885 -152.835 ;
        RECT 2.555 -154.525 2.885 -154.195 ;
        RECT 2.555 -155.885 2.885 -155.555 ;
        RECT 2.555 -157.245 2.885 -156.915 ;
        RECT 2.555 -158.605 2.885 -158.275 ;
        RECT 2.555 -159.965 2.885 -159.635 ;
        RECT 2.555 -161.325 2.885 -160.995 ;
        RECT 2.555 -162.685 2.885 -162.355 ;
        RECT 2.555 -164.045 2.885 -163.715 ;
        RECT 2.555 -165.405 2.885 -165.075 ;
        RECT 2.555 -166.765 2.885 -166.435 ;
        RECT 2.555 -168.125 2.885 -167.795 ;
        RECT 2.555 -169.485 2.885 -169.155 ;
        RECT 2.555 -170.845 2.885 -170.515 ;
        RECT 2.555 -172.205 2.885 -171.875 ;
        RECT 2.555 -173.565 2.885 -173.235 ;
        RECT 2.555 -174.925 2.885 -174.595 ;
        RECT 2.555 -176.285 2.885 -175.955 ;
        RECT 2.555 -177.645 2.885 -177.315 ;
        RECT 2.555 -179.005 2.885 -178.675 ;
        RECT 2.555 -180.365 2.885 -180.035 ;
        RECT 2.555 -181.725 2.885 -181.395 ;
        RECT 2.555 -183.085 2.885 -182.755 ;
        RECT 2.555 -184.445 2.885 -184.115 ;
        RECT 2.555 -185.805 2.885 -185.475 ;
        RECT 2.555 -187.165 2.885 -186.835 ;
        RECT 2.555 -188.525 2.885 -188.195 ;
        RECT 2.555 -189.885 2.885 -189.555 ;
        RECT 2.555 -191.245 2.885 -190.915 ;
        RECT 2.555 -192.605 2.885 -192.275 ;
        RECT 2.555 -193.965 2.885 -193.635 ;
        RECT 2.555 -195.325 2.885 -194.995 ;
        RECT 2.555 -196.685 2.885 -196.355 ;
        RECT 2.555 -198.045 2.885 -197.715 ;
        RECT 2.555 -199.405 2.885 -199.075 ;
        RECT 2.555 -200.765 2.885 -200.435 ;
        RECT 2.555 -202.125 2.885 -201.795 ;
        RECT 2.555 -203.485 2.885 -203.155 ;
        RECT 2.555 -204.845 2.885 -204.515 ;
        RECT 2.555 -206.205 2.885 -205.875 ;
        RECT 2.555 -207.565 2.885 -207.235 ;
        RECT 2.555 -208.925 2.885 -208.595 ;
        RECT 2.555 -210.285 2.885 -209.955 ;
        RECT 2.555 -211.645 2.885 -211.315 ;
        RECT 2.555 -213.005 2.885 -212.675 ;
        RECT 2.555 -214.365 2.885 -214.035 ;
        RECT 2.555 -215.725 2.885 -215.395 ;
        RECT 2.555 -217.085 2.885 -216.755 ;
        RECT 2.555 -218.445 2.885 -218.115 ;
        RECT 2.555 -224.09 2.885 -222.96 ;
        RECT 2.56 -224.205 2.88 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.66 -121.535 2.99 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.915 132.52 4.245 133.65 ;
        RECT 3.915 128.355 4.245 128.685 ;
        RECT 3.915 126.995 4.245 127.325 ;
        RECT 3.915 125.635 4.245 125.965 ;
        RECT 3.915 124.275 4.245 124.605 ;
        RECT 3.92 123.6 4.24 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.275 132.52 5.605 133.65 ;
        RECT 5.275 128.355 5.605 128.685 ;
        RECT 5.275 126.995 5.605 127.325 ;
        RECT 5.275 125.635 5.605 125.965 ;
        RECT 5.275 124.275 5.605 124.605 ;
        RECT 5.28 123.6 5.6 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.275 -0.845 5.605 -0.515 ;
        RECT 5.275 -2.205 5.605 -1.875 ;
        RECT 5.275 -3.565 5.605 -3.235 ;
        RECT 5.28 -3.565 5.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 132.52 6.965 133.65 ;
        RECT 6.635 128.355 6.965 128.685 ;
        RECT 6.635 126.995 6.965 127.325 ;
        RECT 6.635 125.635 6.965 125.965 ;
        RECT 6.635 124.275 6.965 124.605 ;
        RECT 6.64 123.6 6.96 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 -0.845 6.965 -0.515 ;
        RECT 6.635 -2.205 6.965 -1.875 ;
        RECT 6.635 -3.565 6.965 -3.235 ;
        RECT 6.64 -3.565 6.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.995 132.52 8.325 133.65 ;
        RECT 7.995 128.355 8.325 128.685 ;
        RECT 7.995 126.995 8.325 127.325 ;
        RECT 7.995 125.635 8.325 125.965 ;
        RECT 7.995 124.275 8.325 124.605 ;
        RECT 8 123.6 8.32 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.995 -0.845 8.325 -0.515 ;
        RECT 7.995 -2.205 8.325 -1.875 ;
        RECT 7.995 -3.565 8.325 -3.235 ;
        RECT 8 -3.565 8.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.995 -119.165 8.325 -118.835 ;
        RECT 7.995 -120.525 8.325 -120.195 ;
        RECT 7.995 -121.885 8.325 -121.555 ;
        RECT 7.995 -123.245 8.325 -122.915 ;
        RECT 7.995 -124.605 8.325 -124.275 ;
        RECT 7.995 -125.965 8.325 -125.635 ;
        RECT 7.995 -127.325 8.325 -126.995 ;
        RECT 7.995 -128.685 8.325 -128.355 ;
        RECT 7.995 -130.045 8.325 -129.715 ;
        RECT 7.995 -131.405 8.325 -131.075 ;
        RECT 7.995 -132.765 8.325 -132.435 ;
        RECT 7.995 -134.125 8.325 -133.795 ;
        RECT 7.995 -135.485 8.325 -135.155 ;
        RECT 7.995 -136.845 8.325 -136.515 ;
        RECT 7.995 -138.205 8.325 -137.875 ;
        RECT 7.995 -139.565 8.325 -139.235 ;
        RECT 7.995 -140.925 8.325 -140.595 ;
        RECT 7.995 -142.285 8.325 -141.955 ;
        RECT 7.995 -143.645 8.325 -143.315 ;
        RECT 7.995 -145.005 8.325 -144.675 ;
        RECT 7.995 -146.365 8.325 -146.035 ;
        RECT 7.995 -147.725 8.325 -147.395 ;
        RECT 7.995 -149.085 8.325 -148.755 ;
        RECT 7.995 -150.445 8.325 -150.115 ;
        RECT 7.995 -151.805 8.325 -151.475 ;
        RECT 7.995 -153.165 8.325 -152.835 ;
        RECT 7.995 -154.525 8.325 -154.195 ;
        RECT 7.995 -155.885 8.325 -155.555 ;
        RECT 7.995 -157.245 8.325 -156.915 ;
        RECT 7.995 -158.605 8.325 -158.275 ;
        RECT 7.995 -159.965 8.325 -159.635 ;
        RECT 7.995 -161.325 8.325 -160.995 ;
        RECT 7.995 -162.685 8.325 -162.355 ;
        RECT 7.995 -164.045 8.325 -163.715 ;
        RECT 7.995 -165.405 8.325 -165.075 ;
        RECT 7.995 -166.765 8.325 -166.435 ;
        RECT 7.995 -168.125 8.325 -167.795 ;
        RECT 7.995 -169.485 8.325 -169.155 ;
        RECT 7.995 -170.845 8.325 -170.515 ;
        RECT 7.995 -172.205 8.325 -171.875 ;
        RECT 7.995 -173.565 8.325 -173.235 ;
        RECT 7.995 -174.925 8.325 -174.595 ;
        RECT 7.995 -176.285 8.325 -175.955 ;
        RECT 7.995 -177.645 8.325 -177.315 ;
        RECT 7.995 -179.005 8.325 -178.675 ;
        RECT 7.995 -180.365 8.325 -180.035 ;
        RECT 7.995 -181.725 8.325 -181.395 ;
        RECT 7.995 -183.085 8.325 -182.755 ;
        RECT 7.995 -184.445 8.325 -184.115 ;
        RECT 7.995 -185.805 8.325 -185.475 ;
        RECT 7.995 -187.165 8.325 -186.835 ;
        RECT 7.995 -188.525 8.325 -188.195 ;
        RECT 7.995 -189.885 8.325 -189.555 ;
        RECT 7.995 -191.245 8.325 -190.915 ;
        RECT 7.995 -192.605 8.325 -192.275 ;
        RECT 7.995 -193.965 8.325 -193.635 ;
        RECT 7.995 -195.325 8.325 -194.995 ;
        RECT 7.995 -196.685 8.325 -196.355 ;
        RECT 7.995 -198.045 8.325 -197.715 ;
        RECT 7.995 -199.405 8.325 -199.075 ;
        RECT 7.995 -200.765 8.325 -200.435 ;
        RECT 7.995 -202.125 8.325 -201.795 ;
        RECT 7.995 -203.485 8.325 -203.155 ;
        RECT 7.995 -204.845 8.325 -204.515 ;
        RECT 7.995 -206.205 8.325 -205.875 ;
        RECT 7.995 -207.565 8.325 -207.235 ;
        RECT 7.995 -208.925 8.325 -208.595 ;
        RECT 7.995 -210.285 8.325 -209.955 ;
        RECT 7.995 -211.645 8.325 -211.315 ;
        RECT 7.995 -213.005 8.325 -212.675 ;
        RECT 7.995 -214.365 8.325 -214.035 ;
        RECT 7.995 -215.725 8.325 -215.395 ;
        RECT 7.995 -217.085 8.325 -216.755 ;
        RECT 7.995 -218.445 8.325 -218.115 ;
        RECT 7.995 -224.09 8.325 -222.96 ;
        RECT 8 -224.205 8.32 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.76 -121.535 9.09 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 132.52 9.685 133.65 ;
        RECT 9.355 128.355 9.685 128.685 ;
        RECT 9.355 126.995 9.685 127.325 ;
        RECT 9.355 125.635 9.685 125.965 ;
        RECT 9.355 124.275 9.685 124.605 ;
        RECT 9.36 123.6 9.68 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 -123.245 9.685 -122.915 ;
        RECT 9.355 -124.605 9.685 -124.275 ;
        RECT 9.355 -125.965 9.685 -125.635 ;
        RECT 9.355 -127.325 9.685 -126.995 ;
        RECT 9.355 -128.685 9.685 -128.355 ;
        RECT 9.355 -130.045 9.685 -129.715 ;
        RECT 9.355 -131.405 9.685 -131.075 ;
        RECT 9.355 -132.765 9.685 -132.435 ;
        RECT 9.355 -134.125 9.685 -133.795 ;
        RECT 9.355 -135.485 9.685 -135.155 ;
        RECT 9.355 -136.845 9.685 -136.515 ;
        RECT 9.355 -138.205 9.685 -137.875 ;
        RECT 9.355 -139.565 9.685 -139.235 ;
        RECT 9.355 -140.925 9.685 -140.595 ;
        RECT 9.355 -142.285 9.685 -141.955 ;
        RECT 9.355 -143.645 9.685 -143.315 ;
        RECT 9.355 -145.005 9.685 -144.675 ;
        RECT 9.355 -146.365 9.685 -146.035 ;
        RECT 9.355 -147.725 9.685 -147.395 ;
        RECT 9.355 -149.085 9.685 -148.755 ;
        RECT 9.355 -150.445 9.685 -150.115 ;
        RECT 9.355 -151.805 9.685 -151.475 ;
        RECT 9.355 -153.165 9.685 -152.835 ;
        RECT 9.355 -154.525 9.685 -154.195 ;
        RECT 9.355 -155.885 9.685 -155.555 ;
        RECT 9.355 -157.245 9.685 -156.915 ;
        RECT 9.355 -158.605 9.685 -158.275 ;
        RECT 9.355 -159.965 9.685 -159.635 ;
        RECT 9.355 -161.325 9.685 -160.995 ;
        RECT 9.355 -162.685 9.685 -162.355 ;
        RECT 9.355 -164.045 9.685 -163.715 ;
        RECT 9.355 -165.405 9.685 -165.075 ;
        RECT 9.355 -166.765 9.685 -166.435 ;
        RECT 9.355 -168.125 9.685 -167.795 ;
        RECT 9.355 -169.485 9.685 -169.155 ;
        RECT 9.355 -170.845 9.685 -170.515 ;
        RECT 9.355 -172.205 9.685 -171.875 ;
        RECT 9.355 -173.565 9.685 -173.235 ;
        RECT 9.355 -174.925 9.685 -174.595 ;
        RECT 9.355 -176.285 9.685 -175.955 ;
        RECT 9.355 -177.645 9.685 -177.315 ;
        RECT 9.355 -179.005 9.685 -178.675 ;
        RECT 9.355 -180.365 9.685 -180.035 ;
        RECT 9.355 -181.725 9.685 -181.395 ;
        RECT 9.355 -183.085 9.685 -182.755 ;
        RECT 9.355 -184.445 9.685 -184.115 ;
        RECT 9.355 -185.805 9.685 -185.475 ;
        RECT 9.355 -187.165 9.685 -186.835 ;
        RECT 9.355 -188.525 9.685 -188.195 ;
        RECT 9.355 -189.885 9.685 -189.555 ;
        RECT 9.355 -191.245 9.685 -190.915 ;
        RECT 9.355 -192.605 9.685 -192.275 ;
        RECT 9.355 -193.965 9.685 -193.635 ;
        RECT 9.355 -195.325 9.685 -194.995 ;
        RECT 9.355 -196.685 9.685 -196.355 ;
        RECT 9.355 -198.045 9.685 -197.715 ;
        RECT 9.355 -199.405 9.685 -199.075 ;
        RECT 9.355 -200.765 9.685 -200.435 ;
        RECT 9.355 -202.125 9.685 -201.795 ;
        RECT 9.355 -203.485 9.685 -203.155 ;
        RECT 9.355 -204.845 9.685 -204.515 ;
        RECT 9.355 -206.205 9.685 -205.875 ;
        RECT 9.355 -207.565 9.685 -207.235 ;
        RECT 9.355 -208.925 9.685 -208.595 ;
        RECT 9.355 -210.285 9.685 -209.955 ;
        RECT 9.355 -211.645 9.685 -211.315 ;
        RECT 9.355 -213.005 9.685 -212.675 ;
        RECT 9.355 -214.365 9.685 -214.035 ;
        RECT 9.355 -215.725 9.685 -215.395 ;
        RECT 9.355 -217.085 9.685 -216.755 ;
        RECT 9.355 -218.445 9.685 -218.115 ;
        RECT 9.355 -224.09 9.685 -222.96 ;
        RECT 9.36 -224.205 9.68 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.715 132.52 11.045 133.65 ;
        RECT 10.715 128.355 11.045 128.685 ;
        RECT 10.715 126.995 11.045 127.325 ;
        RECT 10.715 125.635 11.045 125.965 ;
        RECT 10.715 124.275 11.045 124.605 ;
        RECT 10.72 123.6 11.04 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.715 -0.845 11.045 -0.515 ;
        RECT 10.715 -2.205 11.045 -1.875 ;
        RECT 10.715 -3.565 11.045 -3.235 ;
        RECT 10.72 -3.565 11.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.075 132.52 12.405 133.65 ;
        RECT 12.075 128.355 12.405 128.685 ;
        RECT 12.075 126.995 12.405 127.325 ;
        RECT 12.075 125.635 12.405 125.965 ;
        RECT 12.075 124.275 12.405 124.605 ;
        RECT 12.08 123.6 12.4 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.075 -0.845 12.405 -0.515 ;
        RECT 12.075 -2.205 12.405 -1.875 ;
        RECT 12.075 -3.565 12.405 -3.235 ;
        RECT 12.08 -3.565 12.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.435 132.52 13.765 133.65 ;
        RECT 13.435 128.355 13.765 128.685 ;
        RECT 13.435 126.995 13.765 127.325 ;
        RECT 13.435 125.635 13.765 125.965 ;
        RECT 13.435 124.275 13.765 124.605 ;
        RECT 13.44 123.6 13.76 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.435 -0.845 13.765 -0.515 ;
        RECT 13.435 -2.205 13.765 -1.875 ;
        RECT 13.435 -3.565 13.765 -3.235 ;
        RECT 13.44 -3.565 13.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.435 -119.165 13.765 -118.835 ;
        RECT 13.435 -120.525 13.765 -120.195 ;
        RECT 13.435 -121.885 13.765 -121.555 ;
        RECT 13.435 -123.245 13.765 -122.915 ;
        RECT 13.435 -124.605 13.765 -124.275 ;
        RECT 13.435 -125.965 13.765 -125.635 ;
        RECT 13.435 -127.325 13.765 -126.995 ;
        RECT 13.435 -128.685 13.765 -128.355 ;
        RECT 13.435 -130.045 13.765 -129.715 ;
        RECT 13.435 -131.405 13.765 -131.075 ;
        RECT 13.435 -132.765 13.765 -132.435 ;
        RECT 13.435 -134.125 13.765 -133.795 ;
        RECT 13.435 -135.485 13.765 -135.155 ;
        RECT 13.435 -136.845 13.765 -136.515 ;
        RECT 13.435 -138.205 13.765 -137.875 ;
        RECT 13.435 -139.565 13.765 -139.235 ;
        RECT 13.435 -140.925 13.765 -140.595 ;
        RECT 13.435 -142.285 13.765 -141.955 ;
        RECT 13.435 -143.645 13.765 -143.315 ;
        RECT 13.435 -145.005 13.765 -144.675 ;
        RECT 13.435 -146.365 13.765 -146.035 ;
        RECT 13.435 -147.725 13.765 -147.395 ;
        RECT 13.435 -149.085 13.765 -148.755 ;
        RECT 13.435 -150.445 13.765 -150.115 ;
        RECT 13.435 -151.805 13.765 -151.475 ;
        RECT 13.435 -153.165 13.765 -152.835 ;
        RECT 13.435 -154.525 13.765 -154.195 ;
        RECT 13.435 -155.885 13.765 -155.555 ;
        RECT 13.435 -157.245 13.765 -156.915 ;
        RECT 13.435 -158.605 13.765 -158.275 ;
        RECT 13.435 -159.965 13.765 -159.635 ;
        RECT 13.435 -161.325 13.765 -160.995 ;
        RECT 13.435 -162.685 13.765 -162.355 ;
        RECT 13.435 -164.045 13.765 -163.715 ;
        RECT 13.435 -165.405 13.765 -165.075 ;
        RECT 13.435 -166.765 13.765 -166.435 ;
        RECT 13.435 -168.125 13.765 -167.795 ;
        RECT 13.435 -169.485 13.765 -169.155 ;
        RECT 13.435 -170.845 13.765 -170.515 ;
        RECT 13.435 -172.205 13.765 -171.875 ;
        RECT 13.435 -173.565 13.765 -173.235 ;
        RECT 13.435 -174.925 13.765 -174.595 ;
        RECT 13.435 -176.285 13.765 -175.955 ;
        RECT 13.435 -177.645 13.765 -177.315 ;
        RECT 13.435 -179.005 13.765 -178.675 ;
        RECT 13.435 -180.365 13.765 -180.035 ;
        RECT 13.435 -181.725 13.765 -181.395 ;
        RECT 13.435 -183.085 13.765 -182.755 ;
        RECT 13.435 -184.445 13.765 -184.115 ;
        RECT 13.435 -185.805 13.765 -185.475 ;
        RECT 13.435 -187.165 13.765 -186.835 ;
        RECT 13.435 -188.525 13.765 -188.195 ;
        RECT 13.435 -189.885 13.765 -189.555 ;
        RECT 13.435 -191.245 13.765 -190.915 ;
        RECT 13.435 -192.605 13.765 -192.275 ;
        RECT 13.435 -193.965 13.765 -193.635 ;
        RECT 13.435 -195.325 13.765 -194.995 ;
        RECT 13.435 -196.685 13.765 -196.355 ;
        RECT 13.435 -198.045 13.765 -197.715 ;
        RECT 13.435 -199.405 13.765 -199.075 ;
        RECT 13.435 -200.765 13.765 -200.435 ;
        RECT 13.435 -202.125 13.765 -201.795 ;
        RECT 13.435 -203.485 13.765 -203.155 ;
        RECT 13.435 -204.845 13.765 -204.515 ;
        RECT 13.435 -206.205 13.765 -205.875 ;
        RECT 13.435 -207.565 13.765 -207.235 ;
        RECT 13.435 -208.925 13.765 -208.595 ;
        RECT 13.435 -210.285 13.765 -209.955 ;
        RECT 13.435 -211.645 13.765 -211.315 ;
        RECT 13.435 -213.005 13.765 -212.675 ;
        RECT 13.435 -214.365 13.765 -214.035 ;
        RECT 13.435 -215.725 13.765 -215.395 ;
        RECT 13.435 -217.085 13.765 -216.755 ;
        RECT 13.435 -218.445 13.765 -218.115 ;
        RECT 13.435 -224.09 13.765 -222.96 ;
        RECT 13.44 -224.205 13.76 -118.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 132.52 15.125 133.65 ;
        RECT 14.795 128.355 15.125 128.685 ;
        RECT 14.795 126.995 15.125 127.325 ;
        RECT 14.795 125.635 15.125 125.965 ;
        RECT 14.795 124.275 15.125 124.605 ;
        RECT 14.8 123.6 15.12 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 -183.085 15.125 -182.755 ;
        RECT 14.795 -184.445 15.125 -184.115 ;
        RECT 14.795 -185.805 15.125 -185.475 ;
        RECT 14.795 -187.165 15.125 -186.835 ;
        RECT 14.795 -188.525 15.125 -188.195 ;
        RECT 14.795 -189.885 15.125 -189.555 ;
        RECT 14.795 -191.245 15.125 -190.915 ;
        RECT 14.795 -192.605 15.125 -192.275 ;
        RECT 14.795 -193.965 15.125 -193.635 ;
        RECT 14.795 -195.325 15.125 -194.995 ;
        RECT 14.795 -196.685 15.125 -196.355 ;
        RECT 14.795 -198.045 15.125 -197.715 ;
        RECT 14.795 -199.405 15.125 -199.075 ;
        RECT 14.795 -200.765 15.125 -200.435 ;
        RECT 14.795 -202.125 15.125 -201.795 ;
        RECT 14.795 -203.485 15.125 -203.155 ;
        RECT 14.795 -204.845 15.125 -204.515 ;
        RECT 14.795 -206.205 15.125 -205.875 ;
        RECT 14.795 -207.565 15.125 -207.235 ;
        RECT 14.795 -208.925 15.125 -208.595 ;
        RECT 14.795 -210.285 15.125 -209.955 ;
        RECT 14.795 -211.645 15.125 -211.315 ;
        RECT 14.795 -213.005 15.125 -212.675 ;
        RECT 14.795 -214.365 15.125 -214.035 ;
        RECT 14.795 -215.725 15.125 -215.395 ;
        RECT 14.795 -217.085 15.125 -216.755 ;
        RECT 14.795 -218.445 15.125 -218.115 ;
        RECT 14.795 -224.09 15.125 -222.96 ;
        RECT 14.8 -224.205 15.12 -122.24 ;
        RECT 14.795 -123.245 15.125 -122.915 ;
        RECT 14.795 -124.605 15.125 -124.275 ;
        RECT 14.795 -125.965 15.125 -125.635 ;
        RECT 14.795 -127.325 15.125 -126.995 ;
        RECT 14.795 -128.685 15.125 -128.355 ;
        RECT 14.795 -130.045 15.125 -129.715 ;
        RECT 14.795 -131.405 15.125 -131.075 ;
        RECT 14.795 -132.765 15.125 -132.435 ;
        RECT 14.795 -134.125 15.125 -133.795 ;
        RECT 14.795 -135.485 15.125 -135.155 ;
        RECT 14.795 -136.845 15.125 -136.515 ;
        RECT 14.795 -138.205 15.125 -137.875 ;
        RECT 14.795 -139.565 15.125 -139.235 ;
        RECT 14.795 -140.925 15.125 -140.595 ;
        RECT 14.795 -142.285 15.125 -141.955 ;
        RECT 14.795 -143.645 15.125 -143.315 ;
        RECT 14.795 -145.005 15.125 -144.675 ;
        RECT 14.795 -146.365 15.125 -146.035 ;
        RECT 14.795 -147.725 15.125 -147.395 ;
        RECT 14.795 -149.085 15.125 -148.755 ;
        RECT 14.795 -150.445 15.125 -150.115 ;
        RECT 14.795 -151.805 15.125 -151.475 ;
        RECT 14.795 -153.165 15.125 -152.835 ;
        RECT 14.795 -154.525 15.125 -154.195 ;
        RECT 14.795 -155.885 15.125 -155.555 ;
        RECT 14.795 -157.245 15.125 -156.915 ;
        RECT 14.795 -158.605 15.125 -158.275 ;
        RECT 14.795 -159.965 15.125 -159.635 ;
        RECT 14.795 -161.325 15.125 -160.995 ;
        RECT 14.795 -162.685 15.125 -162.355 ;
        RECT 14.795 -164.045 15.125 -163.715 ;
        RECT 14.795 -165.405 15.125 -165.075 ;
        RECT 14.795 -166.765 15.125 -166.435 ;
        RECT 14.795 -168.125 15.125 -167.795 ;
        RECT 14.795 -169.485 15.125 -169.155 ;
        RECT 14.795 -170.845 15.125 -170.515 ;
        RECT 14.795 -172.205 15.125 -171.875 ;
        RECT 14.795 -173.565 15.125 -173.235 ;
        RECT 14.795 -174.925 15.125 -174.595 ;
        RECT 14.795 -176.285 15.125 -175.955 ;
        RECT 14.795 -177.645 15.125 -177.315 ;
        RECT 14.795 -179.005 15.125 -178.675 ;
        RECT 14.795 -180.365 15.125 -180.035 ;
        RECT 14.795 -181.725 15.125 -181.395 ;
    END
    PORT
      LAYER met3 ;
        RECT -8.325 132.52 -7.995 133.65 ;
        RECT -8.325 128.355 -7.995 128.685 ;
        RECT -8.325 126.995 -7.995 127.325 ;
        RECT -8.325 125.635 -7.995 125.965 ;
        RECT -8.325 124.275 -7.995 124.605 ;
        RECT -8.325 122.915 -7.995 123.245 ;
        RECT -8.325 121.555 -7.995 121.885 ;
        RECT -8.325 120.195 -7.995 120.525 ;
        RECT -8.325 118.835 -7.995 119.165 ;
        RECT -8.325 117.475 -7.995 117.805 ;
        RECT -8.325 110.675 -7.995 111.005 ;
        RECT -8.325 107.955 -7.995 108.285 ;
        RECT -8.325 103.875 -7.995 104.205 ;
        RECT -8.325 99.795 -7.995 100.125 ;
        RECT -8.325 97.075 -7.995 97.405 ;
        RECT -8.325 90.275 -7.995 90.605 ;
        RECT -8.325 88.915 -7.995 89.245 ;
        RECT -8.325 82.115 -7.995 82.445 ;
        RECT -8.325 79.395 -7.995 79.725 ;
        RECT -8.325 75.315 -7.995 75.645 ;
        RECT -8.325 71.235 -7.995 71.565 ;
        RECT -8.325 68.515 -7.995 68.845 ;
        RECT -8.325 61.715 -7.995 62.045 ;
        RECT -8.325 60.355 -7.995 60.685 ;
        RECT -8.325 50.835 -7.995 51.165 ;
        RECT -8.325 46.755 -7.995 47.085 ;
        RECT -8.325 42.675 -7.995 43.005 ;
        RECT -8.325 39.955 -7.995 40.285 ;
        RECT -8.325 33.155 -7.995 33.485 ;
        RECT -8.325 31.795 -7.995 32.125 ;
        RECT -8.325 29.075 -7.995 29.405 ;
        RECT -8.325 22.275 -7.995 22.605 ;
        RECT -8.325 19.555 -7.995 19.885 ;
        RECT -8.325 18.195 -7.995 18.525 ;
        RECT -8.325 11.395 -7.995 11.725 ;
        RECT -8.325 4.595 -7.995 4.925 ;
        RECT -8.325 3.235 -7.995 3.565 ;
        RECT -8.325 1.875 -7.995 2.205 ;
        RECT -8.325 0.515 -7.995 0.845 ;
        RECT -8.325 -0.845 -7.995 -0.515 ;
        RECT -8.325 -2.205 -7.995 -1.875 ;
        RECT -8.325 -3.565 -7.995 -3.235 ;
        RECT -8.325 -4.925 -7.995 -4.595 ;
        RECT -8.325 -6.285 -7.995 -5.955 ;
        RECT -8.325 -7.645 -7.995 -7.315 ;
        RECT -8.325 -9.005 -7.995 -8.675 ;
        RECT -8.325 -10.365 -7.995 -10.035 ;
        RECT -8.325 -11.725 -7.995 -11.395 ;
        RECT -8.325 -13.085 -7.995 -12.755 ;
        RECT -8.325 -14.445 -7.995 -14.115 ;
        RECT -8.325 -15.805 -7.995 -15.475 ;
        RECT -8.325 -17.165 -7.995 -16.835 ;
        RECT -8.325 -18.525 -7.995 -18.195 ;
        RECT -8.325 -21.245 -7.995 -20.915 ;
        RECT -8.325 -22.605 -7.995 -22.275 ;
        RECT -8.325 -23.965 -7.995 -23.635 ;
        RECT -8.325 -25.325 -7.995 -24.995 ;
        RECT -8.325 -26.685 -7.995 -26.355 ;
        RECT -8.325 -28.045 -7.995 -27.715 ;
        RECT -8.325 -29.405 -7.995 -29.075 ;
        RECT -8.325 -30.765 -7.995 -30.435 ;
        RECT -8.325 -32.125 -7.995 -31.795 ;
        RECT -8.325 -33.485 -7.995 -33.155 ;
        RECT -8.325 -34.845 -7.995 -34.515 ;
        RECT -8.325 -36.205 -7.995 -35.875 ;
        RECT -8.325 -37.565 -7.995 -37.235 ;
        RECT -8.325 -38.925 -7.995 -38.595 ;
        RECT -8.325 -40.285 -7.995 -39.955 ;
        RECT -8.325 -41.645 -7.995 -41.315 ;
        RECT -8.325 -43.005 -7.995 -42.675 ;
        RECT -8.325 -44.365 -7.995 -44.035 ;
        RECT -8.325 -45.725 -7.995 -45.395 ;
        RECT -8.325 -47.085 -7.995 -46.755 ;
        RECT -8.325 -48.445 -7.995 -48.115 ;
        RECT -8.325 -49.805 -7.995 -49.475 ;
        RECT -8.325 -51.165 -7.995 -50.835 ;
        RECT -8.325 -52.525 -7.995 -52.195 ;
        RECT -8.325 -53.885 -7.995 -53.555 ;
        RECT -8.325 -55.245 -7.995 -54.915 ;
        RECT -8.325 -56.605 -7.995 -56.275 ;
        RECT -8.325 -57.965 -7.995 -57.635 ;
        RECT -8.325 -59.325 -7.995 -58.995 ;
        RECT -8.325 -62.045 -7.995 -61.715 ;
        RECT -8.325 -66.125 -7.995 -65.795 ;
        RECT -8.325 -68.845 -7.995 -68.515 ;
        RECT -8.325 -70.205 -7.995 -69.875 ;
        RECT -8.325 -71.565 -7.995 -71.235 ;
        RECT -8.325 -72.925 -7.995 -72.595 ;
        RECT -8.325 -74.285 -7.995 -73.955 ;
        RECT -8.325 -75.645 -7.995 -75.315 ;
        RECT -8.325 -77.005 -7.995 -76.675 ;
        RECT -8.325 -78.365 -7.995 -78.035 ;
        RECT -8.325 -79.725 -7.995 -79.395 ;
        RECT -8.325 -81.085 -7.995 -80.755 ;
        RECT -8.325 -82.445 -7.995 -82.115 ;
        RECT -8.325 -83.805 -7.995 -83.475 ;
        RECT -8.325 -85.165 -7.995 -84.835 ;
        RECT -8.325 -86.525 -7.995 -86.195 ;
        RECT -8.325 -87.885 -7.995 -87.555 ;
        RECT -8.325 -89.245 -7.995 -88.915 ;
        RECT -8.325 -90.605 -7.995 -90.275 ;
        RECT -8.325 -91.965 -7.995 -91.635 ;
        RECT -8.325 -93.325 -7.995 -92.995 ;
        RECT -8.325 -94.685 -7.995 -94.355 ;
        RECT -8.325 -96.045 -7.995 -95.715 ;
        RECT -8.325 -97.405 -7.995 -97.075 ;
        RECT -8.325 -98.765 -7.995 -98.435 ;
        RECT -8.325 -100.125 -7.995 -99.795 ;
        RECT -8.325 -101.485 -7.995 -101.155 ;
        RECT -8.325 -102.845 -7.995 -102.515 ;
        RECT -8.325 -104.205 -7.995 -103.875 ;
        RECT -8.325 -105.565 -7.995 -105.235 ;
        RECT -8.325 -106.925 -7.995 -106.595 ;
        RECT -8.325 -108.285 -7.995 -107.955 ;
        RECT -8.325 -109.645 -7.995 -109.315 ;
        RECT -8.325 -111.005 -7.995 -110.675 ;
        RECT -8.325 -115.085 -7.995 -114.755 ;
        RECT -8.325 -116.445 -7.995 -116.115 ;
        RECT -8.325 -117.805 -7.995 -117.475 ;
        RECT -8.325 -119.165 -7.995 -118.835 ;
        RECT -8.325 -120.525 -7.995 -120.195 ;
        RECT -8.325 -121.885 -7.995 -121.555 ;
        RECT -8.325 -123.245 -7.995 -122.915 ;
        RECT -8.325 -124.605 -7.995 -124.275 ;
        RECT -8.325 -125.965 -7.995 -125.635 ;
        RECT -8.325 -127.325 -7.995 -126.995 ;
        RECT -8.325 -128.685 -7.995 -128.355 ;
        RECT -8.325 -130.045 -7.995 -129.715 ;
        RECT -8.325 -131.405 -7.995 -131.075 ;
        RECT -8.325 -132.765 -7.995 -132.435 ;
        RECT -8.325 -134.125 -7.995 -133.795 ;
        RECT -8.325 -135.485 -7.995 -135.155 ;
        RECT -8.325 -136.845 -7.995 -136.515 ;
        RECT -8.325 -138.205 -7.995 -137.875 ;
        RECT -8.325 -139.565 -7.995 -139.235 ;
        RECT -8.325 -140.925 -7.995 -140.595 ;
        RECT -8.325 -142.285 -7.995 -141.955 ;
        RECT -8.325 -143.645 -7.995 -143.315 ;
        RECT -8.325 -145.005 -7.995 -144.675 ;
        RECT -8.325 -146.365 -7.995 -146.035 ;
        RECT -8.325 -147.725 -7.995 -147.395 ;
        RECT -8.325 -149.085 -7.995 -148.755 ;
        RECT -8.325 -150.445 -7.995 -150.115 ;
        RECT -8.325 -151.805 -7.995 -151.475 ;
        RECT -8.325 -153.165 -7.995 -152.835 ;
        RECT -8.325 -154.525 -7.995 -154.195 ;
        RECT -8.325 -155.885 -7.995 -155.555 ;
        RECT -8.325 -157.245 -7.995 -156.915 ;
        RECT -8.325 -158.605 -7.995 -158.275 ;
        RECT -8.325 -159.965 -7.995 -159.635 ;
        RECT -8.325 -161.325 -7.995 -160.995 ;
        RECT -8.325 -162.685 -7.995 -162.355 ;
        RECT -8.325 -164.045 -7.995 -163.715 ;
        RECT -8.325 -165.405 -7.995 -165.075 ;
        RECT -8.325 -166.765 -7.995 -166.435 ;
        RECT -8.325 -168.125 -7.995 -167.795 ;
        RECT -8.325 -169.485 -7.995 -169.155 ;
        RECT -8.325 -170.845 -7.995 -170.515 ;
        RECT -8.325 -172.205 -7.995 -171.875 ;
        RECT -8.325 -173.565 -7.995 -173.235 ;
        RECT -8.325 -174.925 -7.995 -174.595 ;
        RECT -8.325 -176.285 -7.995 -175.955 ;
        RECT -8.325 -177.645 -7.995 -177.315 ;
        RECT -8.325 -179.005 -7.995 -178.675 ;
        RECT -8.325 -180.365 -7.995 -180.035 ;
        RECT -8.325 -181.725 -7.995 -181.395 ;
        RECT -8.325 -183.085 -7.995 -182.755 ;
        RECT -8.325 -184.445 -7.995 -184.115 ;
        RECT -8.325 -185.805 -7.995 -185.475 ;
        RECT -8.325 -187.165 -7.995 -186.835 ;
        RECT -8.325 -188.525 -7.995 -188.195 ;
        RECT -8.325 -189.885 -7.995 -189.555 ;
        RECT -8.325 -191.245 -7.995 -190.915 ;
        RECT -8.325 -192.605 -7.995 -192.275 ;
        RECT -8.325 -193.965 -7.995 -193.635 ;
        RECT -8.325 -195.325 -7.995 -194.995 ;
        RECT -8.325 -196.685 -7.995 -196.355 ;
        RECT -8.325 -198.045 -7.995 -197.715 ;
        RECT -8.325 -199.405 -7.995 -199.075 ;
        RECT -8.325 -200.765 -7.995 -200.435 ;
        RECT -8.325 -202.125 -7.995 -201.795 ;
        RECT -8.325 -203.485 -7.995 -203.155 ;
        RECT -8.325 -204.845 -7.995 -204.515 ;
        RECT -8.325 -206.205 -7.995 -205.875 ;
        RECT -8.325 -207.565 -7.995 -207.235 ;
        RECT -8.325 -208.925 -7.995 -208.595 ;
        RECT -8.325 -210.285 -7.995 -209.955 ;
        RECT -8.325 -211.645 -7.995 -211.315 ;
        RECT -8.325 -213.005 -7.995 -212.675 ;
        RECT -8.325 -214.365 -7.995 -214.035 ;
        RECT -8.325 -215.725 -7.995 -215.395 ;
        RECT -8.325 -217.085 -7.995 -216.755 ;
        RECT -8.325 -218.445 -7.995 -218.115 ;
        RECT -8.325 -224.09 -7.995 -222.96 ;
        RECT -8.32 -224.205 -8 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -6.965 132.52 -6.635 133.65 ;
        RECT -6.965 128.355 -6.635 128.685 ;
        RECT -6.965 126.995 -6.635 127.325 ;
        RECT -6.965 125.635 -6.635 125.965 ;
        RECT -6.965 124.275 -6.635 124.605 ;
        RECT -6.965 122.915 -6.635 123.245 ;
        RECT -6.965 121.555 -6.635 121.885 ;
        RECT -6.965 120.195 -6.635 120.525 ;
        RECT -6.965 118.835 -6.635 119.165 ;
        RECT -6.965 117.475 -6.635 117.805 ;
        RECT -6.965 110.675 -6.635 111.005 ;
        RECT -6.965 107.955 -6.635 108.285 ;
        RECT -6.965 103.875 -6.635 104.205 ;
        RECT -6.965 99.795 -6.635 100.125 ;
        RECT -6.965 97.075 -6.635 97.405 ;
        RECT -6.965 90.275 -6.635 90.605 ;
        RECT -6.965 88.915 -6.635 89.245 ;
        RECT -6.965 82.115 -6.635 82.445 ;
        RECT -6.965 79.395 -6.635 79.725 ;
        RECT -6.965 75.315 -6.635 75.645 ;
        RECT -6.965 71.235 -6.635 71.565 ;
        RECT -6.965 68.515 -6.635 68.845 ;
        RECT -6.965 61.715 -6.635 62.045 ;
        RECT -6.965 60.355 -6.635 60.685 ;
        RECT -6.965 50.835 -6.635 51.165 ;
        RECT -6.965 46.755 -6.635 47.085 ;
        RECT -6.965 42.675 -6.635 43.005 ;
        RECT -6.965 39.955 -6.635 40.285 ;
        RECT -6.965 33.155 -6.635 33.485 ;
        RECT -6.965 31.795 -6.635 32.125 ;
        RECT -6.965 29.075 -6.635 29.405 ;
        RECT -6.965 22.275 -6.635 22.605 ;
        RECT -6.965 19.555 -6.635 19.885 ;
        RECT -6.965 18.195 -6.635 18.525 ;
        RECT -6.965 11.395 -6.635 11.725 ;
        RECT -6.965 4.595 -6.635 4.925 ;
        RECT -6.965 3.235 -6.635 3.565 ;
        RECT -6.965 1.875 -6.635 2.205 ;
        RECT -6.965 0.515 -6.635 0.845 ;
        RECT -6.965 -0.845 -6.635 -0.515 ;
        RECT -6.965 -2.205 -6.635 -1.875 ;
        RECT -6.965 -3.565 -6.635 -3.235 ;
        RECT -6.965 -4.925 -6.635 -4.595 ;
        RECT -6.965 -6.285 -6.635 -5.955 ;
        RECT -6.965 -7.645 -6.635 -7.315 ;
        RECT -6.965 -9.005 -6.635 -8.675 ;
        RECT -6.965 -10.365 -6.635 -10.035 ;
        RECT -6.965 -11.725 -6.635 -11.395 ;
        RECT -6.965 -13.085 -6.635 -12.755 ;
        RECT -6.965 -14.445 -6.635 -14.115 ;
        RECT -6.965 -15.805 -6.635 -15.475 ;
        RECT -6.965 -17.165 -6.635 -16.835 ;
        RECT -6.965 -18.525 -6.635 -18.195 ;
        RECT -6.965 -21.245 -6.635 -20.915 ;
        RECT -6.965 -22.605 -6.635 -22.275 ;
        RECT -6.965 -23.965 -6.635 -23.635 ;
        RECT -6.965 -25.325 -6.635 -24.995 ;
        RECT -6.965 -26.685 -6.635 -26.355 ;
        RECT -6.965 -28.045 -6.635 -27.715 ;
        RECT -6.965 -29.405 -6.635 -29.075 ;
        RECT -6.965 -30.765 -6.635 -30.435 ;
        RECT -6.965 -32.125 -6.635 -31.795 ;
        RECT -6.965 -33.485 -6.635 -33.155 ;
        RECT -6.965 -34.845 -6.635 -34.515 ;
        RECT -6.965 -36.205 -6.635 -35.875 ;
        RECT -6.965 -37.565 -6.635 -37.235 ;
        RECT -6.965 -38.925 -6.635 -38.595 ;
        RECT -6.965 -40.285 -6.635 -39.955 ;
        RECT -6.965 -41.645 -6.635 -41.315 ;
        RECT -6.965 -43.005 -6.635 -42.675 ;
        RECT -6.965 -44.365 -6.635 -44.035 ;
        RECT -6.965 -45.725 -6.635 -45.395 ;
        RECT -6.965 -47.085 -6.635 -46.755 ;
        RECT -6.965 -48.445 -6.635 -48.115 ;
        RECT -6.965 -49.805 -6.635 -49.475 ;
        RECT -6.965 -51.165 -6.635 -50.835 ;
        RECT -6.965 -52.525 -6.635 -52.195 ;
        RECT -6.965 -53.885 -6.635 -53.555 ;
        RECT -6.965 -55.245 -6.635 -54.915 ;
        RECT -6.965 -56.605 -6.635 -56.275 ;
        RECT -6.965 -57.965 -6.635 -57.635 ;
        RECT -6.965 -59.325 -6.635 -58.995 ;
        RECT -6.965 -62.045 -6.635 -61.715 ;
        RECT -6.965 -66.125 -6.635 -65.795 ;
        RECT -6.965 -68.845 -6.635 -68.515 ;
        RECT -6.965 -70.205 -6.635 -69.875 ;
        RECT -6.965 -71.565 -6.635 -71.235 ;
        RECT -6.965 -72.925 -6.635 -72.595 ;
        RECT -6.965 -74.285 -6.635 -73.955 ;
        RECT -6.965 -75.645 -6.635 -75.315 ;
        RECT -6.965 -77.005 -6.635 -76.675 ;
        RECT -6.965 -78.365 -6.635 -78.035 ;
        RECT -6.965 -79.725 -6.635 -79.395 ;
        RECT -6.965 -81.085 -6.635 -80.755 ;
        RECT -6.965 -82.445 -6.635 -82.115 ;
        RECT -6.965 -83.805 -6.635 -83.475 ;
        RECT -6.965 -85.165 -6.635 -84.835 ;
        RECT -6.965 -86.525 -6.635 -86.195 ;
        RECT -6.965 -87.885 -6.635 -87.555 ;
        RECT -6.965 -89.245 -6.635 -88.915 ;
        RECT -6.965 -90.605 -6.635 -90.275 ;
        RECT -6.965 -91.965 -6.635 -91.635 ;
        RECT -6.965 -93.325 -6.635 -92.995 ;
        RECT -6.965 -94.685 -6.635 -94.355 ;
        RECT -6.965 -96.045 -6.635 -95.715 ;
        RECT -6.965 -97.405 -6.635 -97.075 ;
        RECT -6.965 -98.765 -6.635 -98.435 ;
        RECT -6.965 -100.125 -6.635 -99.795 ;
        RECT -6.965 -101.485 -6.635 -101.155 ;
        RECT -6.965 -102.845 -6.635 -102.515 ;
        RECT -6.965 -104.205 -6.635 -103.875 ;
        RECT -6.965 -105.565 -6.635 -105.235 ;
        RECT -6.965 -106.925 -6.635 -106.595 ;
        RECT -6.965 -108.285 -6.635 -107.955 ;
        RECT -6.965 -109.645 -6.635 -109.315 ;
        RECT -6.965 -111.005 -6.635 -110.675 ;
        RECT -6.965 -115.085 -6.635 -114.755 ;
        RECT -6.965 -116.445 -6.635 -116.115 ;
        RECT -6.965 -117.805 -6.635 -117.475 ;
        RECT -6.965 -119.165 -6.635 -118.835 ;
        RECT -6.965 -120.525 -6.635 -120.195 ;
        RECT -6.965 -121.885 -6.635 -121.555 ;
        RECT -6.965 -123.245 -6.635 -122.915 ;
        RECT -6.965 -124.605 -6.635 -124.275 ;
        RECT -6.965 -125.965 -6.635 -125.635 ;
        RECT -6.965 -127.325 -6.635 -126.995 ;
        RECT -6.965 -128.685 -6.635 -128.355 ;
        RECT -6.965 -130.045 -6.635 -129.715 ;
        RECT -6.965 -131.405 -6.635 -131.075 ;
        RECT -6.965 -132.765 -6.635 -132.435 ;
        RECT -6.965 -134.125 -6.635 -133.795 ;
        RECT -6.965 -135.485 -6.635 -135.155 ;
        RECT -6.965 -136.845 -6.635 -136.515 ;
        RECT -6.965 -138.205 -6.635 -137.875 ;
        RECT -6.965 -139.565 -6.635 -139.235 ;
        RECT -6.965 -140.925 -6.635 -140.595 ;
        RECT -6.965 -142.285 -6.635 -141.955 ;
        RECT -6.965 -143.645 -6.635 -143.315 ;
        RECT -6.965 -145.005 -6.635 -144.675 ;
        RECT -6.965 -146.365 -6.635 -146.035 ;
        RECT -6.965 -147.725 -6.635 -147.395 ;
        RECT -6.965 -149.085 -6.635 -148.755 ;
        RECT -6.965 -150.445 -6.635 -150.115 ;
        RECT -6.965 -151.805 -6.635 -151.475 ;
        RECT -6.965 -153.165 -6.635 -152.835 ;
        RECT -6.965 -154.525 -6.635 -154.195 ;
        RECT -6.965 -155.885 -6.635 -155.555 ;
        RECT -6.965 -157.245 -6.635 -156.915 ;
        RECT -6.965 -158.605 -6.635 -158.275 ;
        RECT -6.965 -159.965 -6.635 -159.635 ;
        RECT -6.965 -161.325 -6.635 -160.995 ;
        RECT -6.965 -162.685 -6.635 -162.355 ;
        RECT -6.965 -164.045 -6.635 -163.715 ;
        RECT -6.965 -165.405 -6.635 -165.075 ;
        RECT -6.965 -166.765 -6.635 -166.435 ;
        RECT -6.965 -168.125 -6.635 -167.795 ;
        RECT -6.965 -169.485 -6.635 -169.155 ;
        RECT -6.965 -170.845 -6.635 -170.515 ;
        RECT -6.965 -172.205 -6.635 -171.875 ;
        RECT -6.965 -173.565 -6.635 -173.235 ;
        RECT -6.965 -174.925 -6.635 -174.595 ;
        RECT -6.965 -176.285 -6.635 -175.955 ;
        RECT -6.965 -177.645 -6.635 -177.315 ;
        RECT -6.965 -179.005 -6.635 -178.675 ;
        RECT -6.965 -180.365 -6.635 -180.035 ;
        RECT -6.965 -181.725 -6.635 -181.395 ;
        RECT -6.965 -183.085 -6.635 -182.755 ;
        RECT -6.965 -184.445 -6.635 -184.115 ;
        RECT -6.965 -185.805 -6.635 -185.475 ;
        RECT -6.965 -187.165 -6.635 -186.835 ;
        RECT -6.965 -188.525 -6.635 -188.195 ;
        RECT -6.965 -189.885 -6.635 -189.555 ;
        RECT -6.965 -191.245 -6.635 -190.915 ;
        RECT -6.965 -192.605 -6.635 -192.275 ;
        RECT -6.965 -193.965 -6.635 -193.635 ;
        RECT -6.965 -195.325 -6.635 -194.995 ;
        RECT -6.965 -196.685 -6.635 -196.355 ;
        RECT -6.965 -198.045 -6.635 -197.715 ;
        RECT -6.965 -199.405 -6.635 -199.075 ;
        RECT -6.965 -200.765 -6.635 -200.435 ;
        RECT -6.965 -202.125 -6.635 -201.795 ;
        RECT -6.965 -203.485 -6.635 -203.155 ;
        RECT -6.965 -204.845 -6.635 -204.515 ;
        RECT -6.965 -206.205 -6.635 -205.875 ;
        RECT -6.965 -207.565 -6.635 -207.235 ;
        RECT -6.965 -208.925 -6.635 -208.595 ;
        RECT -6.965 -210.285 -6.635 -209.955 ;
        RECT -6.965 -211.645 -6.635 -211.315 ;
        RECT -6.965 -213.005 -6.635 -212.675 ;
        RECT -6.965 -214.365 -6.635 -214.035 ;
        RECT -6.965 -215.725 -6.635 -215.395 ;
        RECT -6.965 -217.085 -6.635 -216.755 ;
        RECT -6.965 -218.445 -6.635 -218.115 ;
        RECT -6.965 -224.09 -6.635 -222.96 ;
        RECT -6.96 -224.205 -6.64 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.605 132.52 -5.275 133.65 ;
        RECT -5.605 128.355 -5.275 128.685 ;
        RECT -5.605 126.995 -5.275 127.325 ;
        RECT -5.605 125.635 -5.275 125.965 ;
        RECT -5.605 124.275 -5.275 124.605 ;
        RECT -5.605 121.41 -5.275 121.74 ;
        RECT -5.605 119.235 -5.275 119.565 ;
        RECT -5.605 117.655 -5.275 117.985 ;
        RECT -5.605 116.805 -5.275 117.135 ;
        RECT -5.605 114.495 -5.275 114.825 ;
        RECT -5.605 113.645 -5.275 113.975 ;
        RECT -5.605 111.335 -5.275 111.665 ;
        RECT -5.605 110.485 -5.275 110.815 ;
        RECT -5.605 108.175 -5.275 108.505 ;
        RECT -5.605 107.325 -5.275 107.655 ;
        RECT -5.605 105.015 -5.275 105.345 ;
        RECT -5.605 103.435 -5.275 103.765 ;
        RECT -5.605 102.585 -5.275 102.915 ;
        RECT -5.605 100.275 -5.275 100.605 ;
        RECT -5.605 99.425 -5.275 99.755 ;
        RECT -5.605 97.115 -5.275 97.445 ;
        RECT -5.605 96.265 -5.275 96.595 ;
        RECT -5.605 93.955 -5.275 94.285 ;
        RECT -5.605 93.105 -5.275 93.435 ;
        RECT -5.605 90.795 -5.275 91.125 ;
        RECT -5.605 89.215 -5.275 89.545 ;
        RECT -5.605 88.365 -5.275 88.695 ;
        RECT -5.605 86.055 -5.275 86.385 ;
        RECT -5.605 85.205 -5.275 85.535 ;
        RECT -5.605 82.895 -5.275 83.225 ;
        RECT -5.605 82.045 -5.275 82.375 ;
        RECT -5.605 79.735 -5.275 80.065 ;
        RECT -5.605 78.885 -5.275 79.215 ;
        RECT -5.605 76.575 -5.275 76.905 ;
        RECT -5.605 74.995 -5.275 75.325 ;
        RECT -5.605 74.145 -5.275 74.475 ;
        RECT -5.605 71.835 -5.275 72.165 ;
        RECT -5.605 70.985 -5.275 71.315 ;
        RECT -5.605 68.675 -5.275 69.005 ;
        RECT -5.605 67.825 -5.275 68.155 ;
        RECT -5.605 65.515 -5.275 65.845 ;
        RECT -5.605 64.665 -5.275 64.995 ;
        RECT -5.605 62.355 -5.275 62.685 ;
        RECT -5.605 60.775 -5.275 61.105 ;
        RECT -5.605 59.925 -5.275 60.255 ;
        RECT -5.605 57.615 -5.275 57.945 ;
        RECT -5.605 56.765 -5.275 57.095 ;
        RECT -5.605 54.455 -5.275 54.785 ;
        RECT -5.605 53.605 -5.275 53.935 ;
        RECT -5.605 51.295 -5.275 51.625 ;
        RECT -5.605 50.445 -5.275 50.775 ;
        RECT -5.605 48.135 -5.275 48.465 ;
        RECT -5.605 46.555 -5.275 46.885 ;
        RECT -5.605 45.705 -5.275 46.035 ;
        RECT -5.605 43.395 -5.275 43.725 ;
        RECT -5.605 42.545 -5.275 42.875 ;
        RECT -5.605 40.235 -5.275 40.565 ;
        RECT -5.605 39.385 -5.275 39.715 ;
        RECT -5.605 37.075 -5.275 37.405 ;
        RECT -5.605 36.225 -5.275 36.555 ;
        RECT -5.605 33.915 -5.275 34.245 ;
        RECT -5.605 32.335 -5.275 32.665 ;
        RECT -5.605 31.485 -5.275 31.815 ;
        RECT -5.605 29.175 -5.275 29.505 ;
        RECT -5.605 28.325 -5.275 28.655 ;
        RECT -5.605 26.015 -5.275 26.345 ;
        RECT -5.605 25.165 -5.275 25.495 ;
        RECT -5.605 22.855 -5.275 23.185 ;
        RECT -5.605 22.005 -5.275 22.335 ;
        RECT -5.605 19.695 -5.275 20.025 ;
        RECT -5.605 18.115 -5.275 18.445 ;
        RECT -5.605 17.265 -5.275 17.595 ;
        RECT -5.605 14.955 -5.275 15.285 ;
        RECT -5.605 14.105 -5.275 14.435 ;
        RECT -5.605 11.795 -5.275 12.125 ;
        RECT -5.605 10.945 -5.275 11.275 ;
        RECT -5.605 8.635 -5.275 8.965 ;
        RECT -5.605 7.785 -5.275 8.115 ;
        RECT -5.605 5.475 -5.275 5.805 ;
        RECT -5.605 3.895 -5.275 4.225 ;
        RECT -5.605 3.045 -5.275 3.375 ;
        RECT -5.605 0.87 -5.275 1.2 ;
        RECT -5.605 -0.845 -5.275 -0.515 ;
        RECT -5.605 -2.205 -5.275 -1.875 ;
        RECT -5.605 -3.565 -5.275 -3.235 ;
        RECT -5.605 -4.925 -5.275 -4.595 ;
        RECT -5.605 -6.285 -5.275 -5.955 ;
        RECT -5.605 -7.645 -5.275 -7.315 ;
        RECT -5.605 -9.005 -5.275 -8.675 ;
        RECT -5.605 -10.365 -5.275 -10.035 ;
        RECT -5.605 -11.725 -5.275 -11.395 ;
        RECT -5.605 -13.085 -5.275 -12.755 ;
        RECT -5.605 -14.445 -5.275 -14.115 ;
        RECT -5.605 -15.805 -5.275 -15.475 ;
        RECT -5.605 -17.165 -5.275 -16.835 ;
        RECT -5.605 -18.525 -5.275 -18.195 ;
        RECT -5.605 -21.245 -5.275 -20.915 ;
        RECT -5.605 -22.605 -5.275 -22.275 ;
        RECT -5.605 -23.965 -5.275 -23.635 ;
        RECT -5.605 -25.325 -5.275 -24.995 ;
        RECT -5.605 -26.685 -5.275 -26.355 ;
        RECT -5.605 -28.045 -5.275 -27.715 ;
        RECT -5.605 -29.405 -5.275 -29.075 ;
        RECT -5.605 -30.765 -5.275 -30.435 ;
        RECT -5.605 -32.125 -5.275 -31.795 ;
        RECT -5.605 -33.485 -5.275 -33.155 ;
        RECT -5.605 -34.845 -5.275 -34.515 ;
        RECT -5.605 -36.205 -5.275 -35.875 ;
        RECT -5.605 -37.565 -5.275 -37.235 ;
        RECT -5.605 -38.925 -5.275 -38.595 ;
        RECT -5.605 -40.285 -5.275 -39.955 ;
        RECT -5.605 -41.645 -5.275 -41.315 ;
        RECT -5.605 -43.005 -5.275 -42.675 ;
        RECT -5.605 -44.365 -5.275 -44.035 ;
        RECT -5.605 -45.725 -5.275 -45.395 ;
        RECT -5.605 -47.085 -5.275 -46.755 ;
        RECT -5.605 -48.445 -5.275 -48.115 ;
        RECT -5.605 -49.805 -5.275 -49.475 ;
        RECT -5.605 -51.165 -5.275 -50.835 ;
        RECT -5.605 -52.525 -5.275 -52.195 ;
        RECT -5.605 -53.885 -5.275 -53.555 ;
        RECT -5.605 -55.245 -5.275 -54.915 ;
        RECT -5.605 -56.605 -5.275 -56.275 ;
        RECT -5.605 -57.965 -5.275 -57.635 ;
        RECT -5.605 -59.325 -5.275 -58.995 ;
        RECT -5.605 -62.045 -5.275 -61.715 ;
        RECT -5.605 -66.125 -5.275 -65.795 ;
        RECT -5.605 -68.845 -5.275 -68.515 ;
        RECT -5.605 -70.205 -5.275 -69.875 ;
        RECT -5.605 -71.565 -5.275 -71.235 ;
        RECT -5.605 -72.925 -5.275 -72.595 ;
        RECT -5.605 -74.285 -5.275 -73.955 ;
        RECT -5.605 -75.645 -5.275 -75.315 ;
        RECT -5.605 -77.005 -5.275 -76.675 ;
        RECT -5.605 -78.365 -5.275 -78.035 ;
        RECT -5.605 -79.725 -5.275 -79.395 ;
        RECT -5.605 -81.085 -5.275 -80.755 ;
        RECT -5.605 -82.445 -5.275 -82.115 ;
        RECT -5.605 -83.805 -5.275 -83.475 ;
        RECT -5.605 -85.165 -5.275 -84.835 ;
        RECT -5.605 -86.525 -5.275 -86.195 ;
        RECT -5.605 -87.885 -5.275 -87.555 ;
        RECT -5.605 -89.245 -5.275 -88.915 ;
        RECT -5.605 -90.605 -5.275 -90.275 ;
        RECT -5.605 -91.965 -5.275 -91.635 ;
        RECT -5.605 -93.325 -5.275 -92.995 ;
        RECT -5.605 -94.685 -5.275 -94.355 ;
        RECT -5.605 -96.045 -5.275 -95.715 ;
        RECT -5.605 -97.405 -5.275 -97.075 ;
        RECT -5.605 -98.765 -5.275 -98.435 ;
        RECT -5.605 -100.125 -5.275 -99.795 ;
        RECT -5.605 -101.485 -5.275 -101.155 ;
        RECT -5.605 -102.845 -5.275 -102.515 ;
        RECT -5.605 -104.205 -5.275 -103.875 ;
        RECT -5.605 -105.565 -5.275 -105.235 ;
        RECT -5.605 -106.925 -5.275 -106.595 ;
        RECT -5.605 -108.285 -5.275 -107.955 ;
        RECT -5.605 -109.645 -5.275 -109.315 ;
        RECT -5.605 -111.005 -5.275 -110.675 ;
        RECT -5.605 -115.085 -5.275 -114.755 ;
        RECT -5.605 -116.445 -5.275 -116.115 ;
        RECT -5.605 -117.805 -5.275 -117.475 ;
        RECT -5.605 -119.165 -5.275 -118.835 ;
        RECT -5.605 -120.525 -5.275 -120.195 ;
        RECT -5.605 -121.885 -5.275 -121.555 ;
        RECT -5.605 -123.245 -5.275 -122.915 ;
        RECT -5.605 -124.605 -5.275 -124.275 ;
        RECT -5.605 -125.965 -5.275 -125.635 ;
        RECT -5.605 -127.325 -5.275 -126.995 ;
        RECT -5.605 -128.685 -5.275 -128.355 ;
        RECT -5.605 -130.045 -5.275 -129.715 ;
        RECT -5.605 -131.405 -5.275 -131.075 ;
        RECT -5.605 -132.765 -5.275 -132.435 ;
        RECT -5.605 -134.125 -5.275 -133.795 ;
        RECT -5.605 -135.485 -5.275 -135.155 ;
        RECT -5.605 -136.845 -5.275 -136.515 ;
        RECT -5.605 -138.205 -5.275 -137.875 ;
        RECT -5.605 -139.565 -5.275 -139.235 ;
        RECT -5.605 -140.925 -5.275 -140.595 ;
        RECT -5.605 -142.285 -5.275 -141.955 ;
        RECT -5.605 -143.645 -5.275 -143.315 ;
        RECT -5.605 -145.005 -5.275 -144.675 ;
        RECT -5.605 -146.365 -5.275 -146.035 ;
        RECT -5.605 -147.725 -5.275 -147.395 ;
        RECT -5.605 -149.085 -5.275 -148.755 ;
        RECT -5.605 -150.445 -5.275 -150.115 ;
        RECT -5.605 -151.805 -5.275 -151.475 ;
        RECT -5.605 -153.165 -5.275 -152.835 ;
        RECT -5.605 -154.525 -5.275 -154.195 ;
        RECT -5.605 -155.885 -5.275 -155.555 ;
        RECT -5.605 -157.245 -5.275 -156.915 ;
        RECT -5.605 -158.605 -5.275 -158.275 ;
        RECT -5.605 -159.965 -5.275 -159.635 ;
        RECT -5.605 -161.325 -5.275 -160.995 ;
        RECT -5.605 -162.685 -5.275 -162.355 ;
        RECT -5.605 -164.045 -5.275 -163.715 ;
        RECT -5.605 -165.405 -5.275 -165.075 ;
        RECT -5.605 -166.765 -5.275 -166.435 ;
        RECT -5.605 -168.125 -5.275 -167.795 ;
        RECT -5.605 -169.485 -5.275 -169.155 ;
        RECT -5.605 -170.845 -5.275 -170.515 ;
        RECT -5.605 -172.205 -5.275 -171.875 ;
        RECT -5.605 -173.565 -5.275 -173.235 ;
        RECT -5.605 -174.925 -5.275 -174.595 ;
        RECT -5.605 -176.285 -5.275 -175.955 ;
        RECT -5.605 -177.645 -5.275 -177.315 ;
        RECT -5.605 -179.005 -5.275 -178.675 ;
        RECT -5.605 -180.365 -5.275 -180.035 ;
        RECT -5.605 -181.725 -5.275 -181.395 ;
        RECT -5.605 -183.085 -5.275 -182.755 ;
        RECT -5.605 -184.445 -5.275 -184.115 ;
        RECT -5.605 -185.805 -5.275 -185.475 ;
        RECT -5.605 -187.165 -5.275 -186.835 ;
        RECT -5.605 -188.525 -5.275 -188.195 ;
        RECT -5.605 -189.885 -5.275 -189.555 ;
        RECT -5.605 -191.245 -5.275 -190.915 ;
        RECT -5.605 -192.605 -5.275 -192.275 ;
        RECT -5.605 -193.965 -5.275 -193.635 ;
        RECT -5.605 -195.325 -5.275 -194.995 ;
        RECT -5.605 -196.685 -5.275 -196.355 ;
        RECT -5.605 -198.045 -5.275 -197.715 ;
        RECT -5.605 -199.405 -5.275 -199.075 ;
        RECT -5.605 -200.765 -5.275 -200.435 ;
        RECT -5.605 -202.125 -5.275 -201.795 ;
        RECT -5.605 -203.485 -5.275 -203.155 ;
        RECT -5.605 -204.845 -5.275 -204.515 ;
        RECT -5.605 -206.205 -5.275 -205.875 ;
        RECT -5.605 -207.565 -5.275 -207.235 ;
        RECT -5.605 -208.925 -5.275 -208.595 ;
        RECT -5.605 -210.285 -5.275 -209.955 ;
        RECT -5.605 -211.645 -5.275 -211.315 ;
        RECT -5.605 -213.005 -5.275 -212.675 ;
        RECT -5.605 -214.365 -5.275 -214.035 ;
        RECT -5.605 -215.725 -5.275 -215.395 ;
        RECT -5.605 -217.085 -5.275 -216.755 ;
        RECT -5.605 -218.445 -5.275 -218.115 ;
        RECT -5.605 -224.09 -5.275 -222.96 ;
        RECT -5.6 -224.205 -5.28 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -4.245 132.52 -3.915 133.65 ;
        RECT -4.245 128.355 -3.915 128.685 ;
        RECT -4.245 126.995 -3.915 127.325 ;
        RECT -4.245 125.635 -3.915 125.965 ;
        RECT -4.245 124.275 -3.915 124.605 ;
        RECT -4.245 121.41 -3.915 121.74 ;
        RECT -4.245 119.235 -3.915 119.565 ;
        RECT -4.245 117.655 -3.915 117.985 ;
        RECT -4.245 116.805 -3.915 117.135 ;
        RECT -4.245 114.495 -3.915 114.825 ;
        RECT -4.245 113.645 -3.915 113.975 ;
        RECT -4.245 111.335 -3.915 111.665 ;
        RECT -4.245 110.485 -3.915 110.815 ;
        RECT -4.245 108.175 -3.915 108.505 ;
        RECT -4.245 107.325 -3.915 107.655 ;
        RECT -4.245 105.015 -3.915 105.345 ;
        RECT -4.245 103.435 -3.915 103.765 ;
        RECT -4.245 102.585 -3.915 102.915 ;
        RECT -4.245 100.275 -3.915 100.605 ;
        RECT -4.245 99.425 -3.915 99.755 ;
        RECT -4.245 97.115 -3.915 97.445 ;
        RECT -4.245 96.265 -3.915 96.595 ;
        RECT -4.245 93.955 -3.915 94.285 ;
        RECT -4.245 93.105 -3.915 93.435 ;
        RECT -4.245 90.795 -3.915 91.125 ;
        RECT -4.245 89.215 -3.915 89.545 ;
        RECT -4.245 88.365 -3.915 88.695 ;
        RECT -4.245 86.055 -3.915 86.385 ;
        RECT -4.245 85.205 -3.915 85.535 ;
        RECT -4.245 82.895 -3.915 83.225 ;
        RECT -4.245 82.045 -3.915 82.375 ;
        RECT -4.245 79.735 -3.915 80.065 ;
        RECT -4.245 78.885 -3.915 79.215 ;
        RECT -4.245 76.575 -3.915 76.905 ;
        RECT -4.245 74.995 -3.915 75.325 ;
        RECT -4.245 74.145 -3.915 74.475 ;
        RECT -4.245 71.835 -3.915 72.165 ;
        RECT -4.245 70.985 -3.915 71.315 ;
        RECT -4.245 68.675 -3.915 69.005 ;
        RECT -4.245 67.825 -3.915 68.155 ;
        RECT -4.245 65.515 -3.915 65.845 ;
        RECT -4.245 64.665 -3.915 64.995 ;
        RECT -4.245 62.355 -3.915 62.685 ;
        RECT -4.245 60.775 -3.915 61.105 ;
        RECT -4.245 59.925 -3.915 60.255 ;
        RECT -4.245 57.615 -3.915 57.945 ;
        RECT -4.245 56.765 -3.915 57.095 ;
        RECT -4.245 54.455 -3.915 54.785 ;
        RECT -4.245 53.605 -3.915 53.935 ;
        RECT -4.245 51.295 -3.915 51.625 ;
        RECT -4.245 50.445 -3.915 50.775 ;
        RECT -4.245 48.135 -3.915 48.465 ;
        RECT -4.245 46.555 -3.915 46.885 ;
        RECT -4.245 45.705 -3.915 46.035 ;
        RECT -4.245 43.395 -3.915 43.725 ;
        RECT -4.245 42.545 -3.915 42.875 ;
        RECT -4.245 40.235 -3.915 40.565 ;
        RECT -4.245 39.385 -3.915 39.715 ;
        RECT -4.245 37.075 -3.915 37.405 ;
        RECT -4.245 36.225 -3.915 36.555 ;
        RECT -4.245 33.915 -3.915 34.245 ;
        RECT -4.245 32.335 -3.915 32.665 ;
        RECT -4.245 31.485 -3.915 31.815 ;
        RECT -4.245 29.175 -3.915 29.505 ;
        RECT -4.245 28.325 -3.915 28.655 ;
        RECT -4.245 26.015 -3.915 26.345 ;
        RECT -4.245 25.165 -3.915 25.495 ;
        RECT -4.245 22.855 -3.915 23.185 ;
        RECT -4.245 22.005 -3.915 22.335 ;
        RECT -4.245 19.695 -3.915 20.025 ;
        RECT -4.245 18.115 -3.915 18.445 ;
        RECT -4.245 17.265 -3.915 17.595 ;
        RECT -4.245 14.955 -3.915 15.285 ;
        RECT -4.245 14.105 -3.915 14.435 ;
        RECT -4.245 11.795 -3.915 12.125 ;
        RECT -4.245 10.945 -3.915 11.275 ;
        RECT -4.245 8.635 -3.915 8.965 ;
        RECT -4.245 7.785 -3.915 8.115 ;
        RECT -4.245 5.475 -3.915 5.805 ;
        RECT -4.245 3.895 -3.915 4.225 ;
        RECT -4.245 3.045 -3.915 3.375 ;
        RECT -4.245 0.87 -3.915 1.2 ;
        RECT -4.245 -0.845 -3.915 -0.515 ;
        RECT -4.245 -2.205 -3.915 -1.875 ;
        RECT -4.245 -3.565 -3.915 -3.235 ;
        RECT -4.245 -4.925 -3.915 -4.595 ;
        RECT -4.245 -6.285 -3.915 -5.955 ;
        RECT -4.245 -7.645 -3.915 -7.315 ;
        RECT -4.245 -9.005 -3.915 -8.675 ;
        RECT -4.245 -10.365 -3.915 -10.035 ;
        RECT -4.245 -11.725 -3.915 -11.395 ;
        RECT -4.245 -13.085 -3.915 -12.755 ;
        RECT -4.245 -14.445 -3.915 -14.115 ;
        RECT -4.245 -15.805 -3.915 -15.475 ;
        RECT -4.245 -17.165 -3.915 -16.835 ;
        RECT -4.245 -18.525 -3.915 -18.195 ;
        RECT -4.245 -21.245 -3.915 -20.915 ;
        RECT -4.245 -22.605 -3.915 -22.275 ;
        RECT -4.245 -23.965 -3.915 -23.635 ;
        RECT -4.245 -25.325 -3.915 -24.995 ;
        RECT -4.245 -26.685 -3.915 -26.355 ;
        RECT -4.245 -28.045 -3.915 -27.715 ;
        RECT -4.245 -29.405 -3.915 -29.075 ;
        RECT -4.245 -30.765 -3.915 -30.435 ;
        RECT -4.245 -32.125 -3.915 -31.795 ;
        RECT -4.245 -33.485 -3.915 -33.155 ;
        RECT -4.245 -34.845 -3.915 -34.515 ;
        RECT -4.245 -36.205 -3.915 -35.875 ;
        RECT -4.245 -37.565 -3.915 -37.235 ;
        RECT -4.245 -38.925 -3.915 -38.595 ;
        RECT -4.245 -40.285 -3.915 -39.955 ;
        RECT -4.245 -41.645 -3.915 -41.315 ;
        RECT -4.245 -43.005 -3.915 -42.675 ;
        RECT -4.245 -44.365 -3.915 -44.035 ;
        RECT -4.245 -45.725 -3.915 -45.395 ;
        RECT -4.245 -47.085 -3.915 -46.755 ;
        RECT -4.245 -48.445 -3.915 -48.115 ;
        RECT -4.245 -49.805 -3.915 -49.475 ;
        RECT -4.245 -51.165 -3.915 -50.835 ;
        RECT -4.245 -52.525 -3.915 -52.195 ;
        RECT -4.245 -53.885 -3.915 -53.555 ;
        RECT -4.245 -55.245 -3.915 -54.915 ;
        RECT -4.245 -56.605 -3.915 -56.275 ;
        RECT -4.245 -57.965 -3.915 -57.635 ;
        RECT -4.245 -59.325 -3.915 -58.995 ;
        RECT -4.245 -62.045 -3.915 -61.715 ;
        RECT -4.245 -66.125 -3.915 -65.795 ;
        RECT -4.245 -68.845 -3.915 -68.515 ;
        RECT -4.245 -70.205 -3.915 -69.875 ;
        RECT -4.245 -71.565 -3.915 -71.235 ;
        RECT -4.245 -72.925 -3.915 -72.595 ;
        RECT -4.245 -74.285 -3.915 -73.955 ;
        RECT -4.245 -75.645 -3.915 -75.315 ;
        RECT -4.245 -77.005 -3.915 -76.675 ;
        RECT -4.245 -78.365 -3.915 -78.035 ;
        RECT -4.245 -79.725 -3.915 -79.395 ;
        RECT -4.245 -81.085 -3.915 -80.755 ;
        RECT -4.245 -82.445 -3.915 -82.115 ;
        RECT -4.245 -83.805 -3.915 -83.475 ;
        RECT -4.245 -85.165 -3.915 -84.835 ;
        RECT -4.245 -86.525 -3.915 -86.195 ;
        RECT -4.245 -87.885 -3.915 -87.555 ;
        RECT -4.245 -89.245 -3.915 -88.915 ;
        RECT -4.245 -90.605 -3.915 -90.275 ;
        RECT -4.245 -91.965 -3.915 -91.635 ;
        RECT -4.245 -93.325 -3.915 -92.995 ;
        RECT -4.245 -94.685 -3.915 -94.355 ;
        RECT -4.245 -96.045 -3.915 -95.715 ;
        RECT -4.245 -97.405 -3.915 -97.075 ;
        RECT -4.245 -98.765 -3.915 -98.435 ;
        RECT -4.245 -100.125 -3.915 -99.795 ;
        RECT -4.245 -101.485 -3.915 -101.155 ;
        RECT -4.245 -102.845 -3.915 -102.515 ;
        RECT -4.245 -104.205 -3.915 -103.875 ;
        RECT -4.245 -105.565 -3.915 -105.235 ;
        RECT -4.245 -106.925 -3.915 -106.595 ;
        RECT -4.245 -108.285 -3.915 -107.955 ;
        RECT -4.245 -109.645 -3.915 -109.315 ;
        RECT -4.245 -111.005 -3.915 -110.675 ;
        RECT -4.245 -115.085 -3.915 -114.755 ;
        RECT -4.245 -116.445 -3.915 -116.115 ;
        RECT -4.245 -117.805 -3.915 -117.475 ;
        RECT -4.245 -119.165 -3.915 -118.835 ;
        RECT -4.245 -120.525 -3.915 -120.195 ;
        RECT -4.245 -121.885 -3.915 -121.555 ;
        RECT -4.245 -123.245 -3.915 -122.915 ;
        RECT -4.245 -124.605 -3.915 -124.275 ;
        RECT -4.245 -125.965 -3.915 -125.635 ;
        RECT -4.245 -127.325 -3.915 -126.995 ;
        RECT -4.245 -128.685 -3.915 -128.355 ;
        RECT -4.245 -130.045 -3.915 -129.715 ;
        RECT -4.245 -131.405 -3.915 -131.075 ;
        RECT -4.245 -132.765 -3.915 -132.435 ;
        RECT -4.245 -134.125 -3.915 -133.795 ;
        RECT -4.245 -135.485 -3.915 -135.155 ;
        RECT -4.245 -136.845 -3.915 -136.515 ;
        RECT -4.245 -138.205 -3.915 -137.875 ;
        RECT -4.245 -139.565 -3.915 -139.235 ;
        RECT -4.245 -140.925 -3.915 -140.595 ;
        RECT -4.245 -142.285 -3.915 -141.955 ;
        RECT -4.245 -143.645 -3.915 -143.315 ;
        RECT -4.245 -145.005 -3.915 -144.675 ;
        RECT -4.245 -146.365 -3.915 -146.035 ;
        RECT -4.245 -147.725 -3.915 -147.395 ;
        RECT -4.245 -149.085 -3.915 -148.755 ;
        RECT -4.245 -150.445 -3.915 -150.115 ;
        RECT -4.245 -151.805 -3.915 -151.475 ;
        RECT -4.245 -153.165 -3.915 -152.835 ;
        RECT -4.245 -154.525 -3.915 -154.195 ;
        RECT -4.245 -155.885 -3.915 -155.555 ;
        RECT -4.245 -157.245 -3.915 -156.915 ;
        RECT -4.245 -158.605 -3.915 -158.275 ;
        RECT -4.245 -159.965 -3.915 -159.635 ;
        RECT -4.245 -161.325 -3.915 -160.995 ;
        RECT -4.245 -162.685 -3.915 -162.355 ;
        RECT -4.245 -164.045 -3.915 -163.715 ;
        RECT -4.245 -165.405 -3.915 -165.075 ;
        RECT -4.245 -166.765 -3.915 -166.435 ;
        RECT -4.245 -168.125 -3.915 -167.795 ;
        RECT -4.245 -169.485 -3.915 -169.155 ;
        RECT -4.245 -170.845 -3.915 -170.515 ;
        RECT -4.245 -172.205 -3.915 -171.875 ;
        RECT -4.245 -173.565 -3.915 -173.235 ;
        RECT -4.245 -174.925 -3.915 -174.595 ;
        RECT -4.245 -176.285 -3.915 -175.955 ;
        RECT -4.245 -177.645 -3.915 -177.315 ;
        RECT -4.245 -179.005 -3.915 -178.675 ;
        RECT -4.245 -180.365 -3.915 -180.035 ;
        RECT -4.245 -181.725 -3.915 -181.395 ;
        RECT -4.245 -183.085 -3.915 -182.755 ;
        RECT -4.245 -184.445 -3.915 -184.115 ;
        RECT -4.245 -185.805 -3.915 -185.475 ;
        RECT -4.245 -187.165 -3.915 -186.835 ;
        RECT -4.245 -188.525 -3.915 -188.195 ;
        RECT -4.245 -189.885 -3.915 -189.555 ;
        RECT -4.245 -191.245 -3.915 -190.915 ;
        RECT -4.245 -192.605 -3.915 -192.275 ;
        RECT -4.245 -193.965 -3.915 -193.635 ;
        RECT -4.245 -195.325 -3.915 -194.995 ;
        RECT -4.245 -196.685 -3.915 -196.355 ;
        RECT -4.245 -198.045 -3.915 -197.715 ;
        RECT -4.245 -199.405 -3.915 -199.075 ;
        RECT -4.245 -200.765 -3.915 -200.435 ;
        RECT -4.245 -202.125 -3.915 -201.795 ;
        RECT -4.245 -203.485 -3.915 -203.155 ;
        RECT -4.245 -204.845 -3.915 -204.515 ;
        RECT -4.245 -206.205 -3.915 -205.875 ;
        RECT -4.245 -207.565 -3.915 -207.235 ;
        RECT -4.245 -208.925 -3.915 -208.595 ;
        RECT -4.245 -210.285 -3.915 -209.955 ;
        RECT -4.245 -211.645 -3.915 -211.315 ;
        RECT -4.245 -213.005 -3.915 -212.675 ;
        RECT -4.245 -214.365 -3.915 -214.035 ;
        RECT -4.245 -215.725 -3.915 -215.395 ;
        RECT -4.245 -217.085 -3.915 -216.755 ;
        RECT -4.245 -218.445 -3.915 -218.115 ;
        RECT -4.245 -224.09 -3.915 -222.96 ;
        RECT -4.24 -224.205 -3.92 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -2.885 -139.565 -2.555 -139.235 ;
        RECT -2.885 -140.925 -2.555 -140.595 ;
        RECT -2.885 -142.285 -2.555 -141.955 ;
        RECT -2.885 -143.645 -2.555 -143.315 ;
        RECT -2.885 -145.005 -2.555 -144.675 ;
        RECT -2.885 -146.365 -2.555 -146.035 ;
        RECT -2.885 -147.725 -2.555 -147.395 ;
        RECT -2.885 -149.085 -2.555 -148.755 ;
        RECT -2.885 -150.445 -2.555 -150.115 ;
        RECT -2.885 -151.805 -2.555 -151.475 ;
        RECT -2.885 -153.165 -2.555 -152.835 ;
        RECT -2.885 -154.525 -2.555 -154.195 ;
        RECT -2.885 -155.885 -2.555 -155.555 ;
        RECT -2.885 -157.245 -2.555 -156.915 ;
        RECT -2.885 -158.605 -2.555 -158.275 ;
        RECT -2.885 -159.965 -2.555 -159.635 ;
        RECT -2.885 -161.325 -2.555 -160.995 ;
        RECT -2.885 -162.685 -2.555 -162.355 ;
        RECT -2.885 -164.045 -2.555 -163.715 ;
        RECT -2.885 -165.405 -2.555 -165.075 ;
        RECT -2.885 -166.765 -2.555 -166.435 ;
        RECT -2.885 -168.125 -2.555 -167.795 ;
        RECT -2.885 -169.485 -2.555 -169.155 ;
        RECT -2.885 -170.845 -2.555 -170.515 ;
        RECT -2.885 -172.205 -2.555 -171.875 ;
        RECT -2.885 -173.565 -2.555 -173.235 ;
        RECT -2.885 -174.925 -2.555 -174.595 ;
        RECT -2.885 -176.285 -2.555 -175.955 ;
        RECT -2.885 -177.645 -2.555 -177.315 ;
        RECT -2.885 -179.005 -2.555 -178.675 ;
        RECT -2.885 -180.365 -2.555 -180.035 ;
        RECT -2.885 -181.725 -2.555 -181.395 ;
        RECT -2.885 -183.085 -2.555 -182.755 ;
        RECT -2.885 -184.445 -2.555 -184.115 ;
        RECT -2.885 -185.805 -2.555 -185.475 ;
        RECT -2.885 -187.165 -2.555 -186.835 ;
        RECT -2.885 -188.525 -2.555 -188.195 ;
        RECT -2.885 -189.885 -2.555 -189.555 ;
        RECT -2.885 -191.245 -2.555 -190.915 ;
        RECT -2.885 -192.605 -2.555 -192.275 ;
        RECT -2.885 -193.965 -2.555 -193.635 ;
        RECT -2.885 -195.325 -2.555 -194.995 ;
        RECT -2.885 -196.685 -2.555 -196.355 ;
        RECT -2.885 -198.045 -2.555 -197.715 ;
        RECT -2.885 -199.405 -2.555 -199.075 ;
        RECT -2.885 -200.765 -2.555 -200.435 ;
        RECT -2.885 -202.125 -2.555 -201.795 ;
        RECT -2.885 -203.485 -2.555 -203.155 ;
        RECT -2.885 -204.845 -2.555 -204.515 ;
        RECT -2.885 -206.205 -2.555 -205.875 ;
        RECT -2.885 -207.565 -2.555 -207.235 ;
        RECT -2.885 -208.925 -2.555 -208.595 ;
        RECT -2.885 -210.285 -2.555 -209.955 ;
        RECT -2.885 -211.645 -2.555 -211.315 ;
        RECT -2.885 -213.005 -2.555 -212.675 ;
        RECT -2.885 -214.365 -2.555 -214.035 ;
        RECT -2.885 -215.725 -2.555 -215.395 ;
        RECT -2.885 -217.085 -2.555 -216.755 ;
        RECT -2.885 -218.445 -2.555 -218.115 ;
        RECT -2.885 -224.09 -2.555 -222.96 ;
        RECT -2.88 -224.205 -2.56 133.765 ;
        RECT -2.885 132.52 -2.555 133.65 ;
        RECT -2.885 128.355 -2.555 128.685 ;
        RECT -2.885 126.995 -2.555 127.325 ;
        RECT -2.885 125.635 -2.555 125.965 ;
        RECT -2.885 124.275 -2.555 124.605 ;
        RECT -2.885 121.41 -2.555 121.74 ;
        RECT -2.885 119.235 -2.555 119.565 ;
        RECT -2.885 117.655 -2.555 117.985 ;
        RECT -2.885 116.805 -2.555 117.135 ;
        RECT -2.885 114.495 -2.555 114.825 ;
        RECT -2.885 113.645 -2.555 113.975 ;
        RECT -2.885 111.335 -2.555 111.665 ;
        RECT -2.885 110.485 -2.555 110.815 ;
        RECT -2.885 108.175 -2.555 108.505 ;
        RECT -2.885 107.325 -2.555 107.655 ;
        RECT -2.885 105.015 -2.555 105.345 ;
        RECT -2.885 103.435 -2.555 103.765 ;
        RECT -2.885 102.585 -2.555 102.915 ;
        RECT -2.885 100.275 -2.555 100.605 ;
        RECT -2.885 99.425 -2.555 99.755 ;
        RECT -2.885 97.115 -2.555 97.445 ;
        RECT -2.885 96.265 -2.555 96.595 ;
        RECT -2.885 93.955 -2.555 94.285 ;
        RECT -2.885 93.105 -2.555 93.435 ;
        RECT -2.885 90.795 -2.555 91.125 ;
        RECT -2.885 89.215 -2.555 89.545 ;
        RECT -2.885 88.365 -2.555 88.695 ;
        RECT -2.885 86.055 -2.555 86.385 ;
        RECT -2.885 85.205 -2.555 85.535 ;
        RECT -2.885 82.895 -2.555 83.225 ;
        RECT -2.885 82.045 -2.555 82.375 ;
        RECT -2.885 79.735 -2.555 80.065 ;
        RECT -2.885 78.885 -2.555 79.215 ;
        RECT -2.885 76.575 -2.555 76.905 ;
        RECT -2.885 74.995 -2.555 75.325 ;
        RECT -2.885 74.145 -2.555 74.475 ;
        RECT -2.885 71.835 -2.555 72.165 ;
        RECT -2.885 70.985 -2.555 71.315 ;
        RECT -2.885 68.675 -2.555 69.005 ;
        RECT -2.885 67.825 -2.555 68.155 ;
        RECT -2.885 65.515 -2.555 65.845 ;
        RECT -2.885 64.665 -2.555 64.995 ;
        RECT -2.885 62.355 -2.555 62.685 ;
        RECT -2.885 60.775 -2.555 61.105 ;
        RECT -2.885 59.925 -2.555 60.255 ;
        RECT -2.885 57.615 -2.555 57.945 ;
        RECT -2.885 56.765 -2.555 57.095 ;
        RECT -2.885 54.455 -2.555 54.785 ;
        RECT -2.885 53.605 -2.555 53.935 ;
        RECT -2.885 51.295 -2.555 51.625 ;
        RECT -2.885 50.445 -2.555 50.775 ;
        RECT -2.885 48.135 -2.555 48.465 ;
        RECT -2.885 46.555 -2.555 46.885 ;
        RECT -2.885 45.705 -2.555 46.035 ;
        RECT -2.885 43.395 -2.555 43.725 ;
        RECT -2.885 42.545 -2.555 42.875 ;
        RECT -2.885 40.235 -2.555 40.565 ;
        RECT -2.885 39.385 -2.555 39.715 ;
        RECT -2.885 37.075 -2.555 37.405 ;
        RECT -2.885 36.225 -2.555 36.555 ;
        RECT -2.885 33.915 -2.555 34.245 ;
        RECT -2.885 32.335 -2.555 32.665 ;
        RECT -2.885 31.485 -2.555 31.815 ;
        RECT -2.885 29.175 -2.555 29.505 ;
        RECT -2.885 28.325 -2.555 28.655 ;
        RECT -2.885 26.015 -2.555 26.345 ;
        RECT -2.885 25.165 -2.555 25.495 ;
        RECT -2.885 22.855 -2.555 23.185 ;
        RECT -2.885 22.005 -2.555 22.335 ;
        RECT -2.885 19.695 -2.555 20.025 ;
        RECT -2.885 18.115 -2.555 18.445 ;
        RECT -2.885 17.265 -2.555 17.595 ;
        RECT -2.885 14.955 -2.555 15.285 ;
        RECT -2.885 14.105 -2.555 14.435 ;
        RECT -2.885 11.795 -2.555 12.125 ;
        RECT -2.885 10.945 -2.555 11.275 ;
        RECT -2.885 8.635 -2.555 8.965 ;
        RECT -2.885 7.785 -2.555 8.115 ;
        RECT -2.885 5.475 -2.555 5.805 ;
        RECT -2.885 3.895 -2.555 4.225 ;
        RECT -2.885 3.045 -2.555 3.375 ;
        RECT -2.885 0.87 -2.555 1.2 ;
        RECT -2.885 -0.845 -2.555 -0.515 ;
        RECT -2.885 -2.205 -2.555 -1.875 ;
        RECT -2.885 -3.565 -2.555 -3.235 ;
        RECT -2.885 -4.925 -2.555 -4.595 ;
        RECT -2.885 -6.285 -2.555 -5.955 ;
        RECT -2.885 -7.645 -2.555 -7.315 ;
        RECT -2.885 -9.005 -2.555 -8.675 ;
        RECT -2.885 -10.365 -2.555 -10.035 ;
        RECT -2.885 -11.725 -2.555 -11.395 ;
        RECT -2.885 -13.085 -2.555 -12.755 ;
        RECT -2.885 -14.445 -2.555 -14.115 ;
        RECT -2.885 -15.805 -2.555 -15.475 ;
        RECT -2.885 -17.165 -2.555 -16.835 ;
        RECT -2.885 -18.525 -2.555 -18.195 ;
        RECT -2.885 -21.245 -2.555 -20.915 ;
        RECT -2.885 -22.605 -2.555 -22.275 ;
        RECT -2.885 -23.965 -2.555 -23.635 ;
        RECT -2.885 -25.325 -2.555 -24.995 ;
        RECT -2.885 -26.685 -2.555 -26.355 ;
        RECT -2.885 -28.045 -2.555 -27.715 ;
        RECT -2.885 -29.405 -2.555 -29.075 ;
        RECT -2.885 -30.765 -2.555 -30.435 ;
        RECT -2.885 -32.125 -2.555 -31.795 ;
        RECT -2.885 -33.485 -2.555 -33.155 ;
        RECT -2.885 -34.845 -2.555 -34.515 ;
        RECT -2.885 -36.205 -2.555 -35.875 ;
        RECT -2.885 -37.565 -2.555 -37.235 ;
        RECT -2.885 -38.925 -2.555 -38.595 ;
        RECT -2.885 -40.285 -2.555 -39.955 ;
        RECT -2.885 -41.645 -2.555 -41.315 ;
        RECT -2.885 -43.005 -2.555 -42.675 ;
        RECT -2.885 -44.365 -2.555 -44.035 ;
        RECT -2.885 -45.725 -2.555 -45.395 ;
        RECT -2.885 -47.085 -2.555 -46.755 ;
        RECT -2.885 -48.445 -2.555 -48.115 ;
        RECT -2.885 -49.805 -2.555 -49.475 ;
        RECT -2.885 -51.165 -2.555 -50.835 ;
        RECT -2.885 -52.525 -2.555 -52.195 ;
        RECT -2.885 -53.885 -2.555 -53.555 ;
        RECT -2.885 -55.245 -2.555 -54.915 ;
        RECT -2.885 -56.605 -2.555 -56.275 ;
        RECT -2.885 -57.965 -2.555 -57.635 ;
        RECT -2.885 -59.325 -2.555 -58.995 ;
        RECT -2.885 -62.045 -2.555 -61.715 ;
        RECT -2.885 -66.125 -2.555 -65.795 ;
        RECT -2.885 -68.845 -2.555 -68.515 ;
        RECT -2.885 -70.205 -2.555 -69.875 ;
        RECT -2.885 -71.565 -2.555 -71.235 ;
        RECT -2.885 -72.925 -2.555 -72.595 ;
        RECT -2.885 -74.285 -2.555 -73.955 ;
        RECT -2.885 -75.645 -2.555 -75.315 ;
        RECT -2.885 -77.005 -2.555 -76.675 ;
        RECT -2.885 -78.365 -2.555 -78.035 ;
        RECT -2.885 -79.725 -2.555 -79.395 ;
        RECT -2.885 -81.085 -2.555 -80.755 ;
        RECT -2.885 -82.445 -2.555 -82.115 ;
        RECT -2.885 -83.805 -2.555 -83.475 ;
        RECT -2.885 -85.165 -2.555 -84.835 ;
        RECT -2.885 -86.525 -2.555 -86.195 ;
        RECT -2.885 -87.885 -2.555 -87.555 ;
        RECT -2.885 -89.245 -2.555 -88.915 ;
        RECT -2.885 -90.605 -2.555 -90.275 ;
        RECT -2.885 -91.965 -2.555 -91.635 ;
        RECT -2.885 -93.325 -2.555 -92.995 ;
        RECT -2.885 -94.685 -2.555 -94.355 ;
        RECT -2.885 -96.045 -2.555 -95.715 ;
        RECT -2.885 -97.405 -2.555 -97.075 ;
        RECT -2.885 -98.765 -2.555 -98.435 ;
        RECT -2.885 -100.125 -2.555 -99.795 ;
        RECT -2.885 -101.485 -2.555 -101.155 ;
        RECT -2.885 -102.845 -2.555 -102.515 ;
        RECT -2.885 -104.205 -2.555 -103.875 ;
        RECT -2.885 -105.565 -2.555 -105.235 ;
        RECT -2.885 -106.925 -2.555 -106.595 ;
        RECT -2.885 -108.285 -2.555 -107.955 ;
        RECT -2.885 -109.645 -2.555 -109.315 ;
        RECT -2.885 -111.005 -2.555 -110.675 ;
        RECT -2.885 -115.085 -2.555 -114.755 ;
        RECT -2.885 -116.445 -2.555 -116.115 ;
        RECT -2.885 -117.805 -2.555 -117.475 ;
        RECT -2.885 -119.165 -2.555 -118.835 ;
        RECT -2.885 -120.525 -2.555 -120.195 ;
        RECT -2.885 -121.885 -2.555 -121.555 ;
        RECT -2.885 -123.245 -2.555 -122.915 ;
        RECT -2.885 -124.605 -2.555 -124.275 ;
        RECT -2.885 -125.965 -2.555 -125.635 ;
        RECT -2.885 -127.325 -2.555 -126.995 ;
        RECT -2.885 -128.685 -2.555 -128.355 ;
        RECT -2.885 -130.045 -2.555 -129.715 ;
        RECT -2.885 -131.405 -2.555 -131.075 ;
        RECT -2.885 -132.765 -2.555 -132.435 ;
        RECT -2.885 -134.125 -2.555 -133.795 ;
        RECT -2.885 -135.485 -2.555 -135.155 ;
        RECT -2.885 -136.845 -2.555 -136.515 ;
        RECT -2.885 -138.205 -2.555 -137.875 ;
    END
    PORT
      LAYER met3 ;
        RECT -16.485 132.52 -16.155 133.65 ;
        RECT -16.485 128.355 -16.155 128.685 ;
        RECT -16.485 126.995 -16.155 127.325 ;
        RECT -16.485 125.635 -16.155 125.965 ;
        RECT -16.485 124.275 -16.155 124.605 ;
        RECT -16.485 122.915 -16.155 123.245 ;
        RECT -16.485 121.555 -16.155 121.885 ;
        RECT -16.485 120.195 -16.155 120.525 ;
        RECT -16.485 118.835 -16.155 119.165 ;
        RECT -16.485 117.475 -16.155 117.805 ;
        RECT -16.485 116.115 -16.155 116.445 ;
        RECT -16.485 114.755 -16.155 115.085 ;
        RECT -16.485 113.395 -16.155 113.725 ;
        RECT -16.485 112.035 -16.155 112.365 ;
        RECT -16.485 110.675 -16.155 111.005 ;
        RECT -16.485 109.315 -16.155 109.645 ;
        RECT -16.485 107.955 -16.155 108.285 ;
        RECT -16.485 106.595 -16.155 106.925 ;
        RECT -16.485 105.235 -16.155 105.565 ;
        RECT -16.485 103.875 -16.155 104.205 ;
        RECT -16.485 102.515 -16.155 102.845 ;
        RECT -16.485 101.155 -16.155 101.485 ;
        RECT -16.485 99.795 -16.155 100.125 ;
        RECT -16.485 98.435 -16.155 98.765 ;
        RECT -16.485 97.075 -16.155 97.405 ;
        RECT -16.485 95.715 -16.155 96.045 ;
        RECT -16.485 94.355 -16.155 94.685 ;
        RECT -16.485 92.995 -16.155 93.325 ;
        RECT -16.485 91.635 -16.155 91.965 ;
        RECT -16.485 90.275 -16.155 90.605 ;
        RECT -16.485 88.915 -16.155 89.245 ;
        RECT -16.485 87.555 -16.155 87.885 ;
        RECT -16.485 86.195 -16.155 86.525 ;
        RECT -16.485 84.835 -16.155 85.165 ;
        RECT -16.485 83.475 -16.155 83.805 ;
        RECT -16.485 82.115 -16.155 82.445 ;
        RECT -16.485 80.755 -16.155 81.085 ;
        RECT -16.485 79.395 -16.155 79.725 ;
        RECT -16.485 78.035 -16.155 78.365 ;
        RECT -16.485 76.675 -16.155 77.005 ;
        RECT -16.485 75.315 -16.155 75.645 ;
        RECT -16.485 73.955 -16.155 74.285 ;
        RECT -16.485 72.595 -16.155 72.925 ;
        RECT -16.485 71.235 -16.155 71.565 ;
        RECT -16.485 69.875 -16.155 70.205 ;
        RECT -16.485 68.515 -16.155 68.845 ;
        RECT -16.485 67.155 -16.155 67.485 ;
        RECT -16.485 65.795 -16.155 66.125 ;
        RECT -16.485 64.435 -16.155 64.765 ;
        RECT -16.485 63.075 -16.155 63.405 ;
        RECT -16.485 61.715 -16.155 62.045 ;
        RECT -16.485 60.355 -16.155 60.685 ;
        RECT -16.485 58.995 -16.155 59.325 ;
        RECT -16.485 57.635 -16.155 57.965 ;
        RECT -16.485 56.275 -16.155 56.605 ;
        RECT -16.485 54.915 -16.155 55.245 ;
        RECT -16.485 53.555 -16.155 53.885 ;
        RECT -16.485 52.195 -16.155 52.525 ;
        RECT -16.485 50.835 -16.155 51.165 ;
        RECT -16.485 49.475 -16.155 49.805 ;
        RECT -16.485 48.115 -16.155 48.445 ;
        RECT -16.485 46.755 -16.155 47.085 ;
        RECT -16.485 45.395 -16.155 45.725 ;
        RECT -16.485 44.035 -16.155 44.365 ;
        RECT -16.485 42.675 -16.155 43.005 ;
        RECT -16.485 41.315 -16.155 41.645 ;
        RECT -16.485 39.955 -16.155 40.285 ;
        RECT -16.485 38.595 -16.155 38.925 ;
        RECT -16.485 37.235 -16.155 37.565 ;
        RECT -16.485 35.875 -16.155 36.205 ;
        RECT -16.485 34.515 -16.155 34.845 ;
        RECT -16.485 33.155 -16.155 33.485 ;
        RECT -16.485 31.795 -16.155 32.125 ;
        RECT -16.485 30.435 -16.155 30.765 ;
        RECT -16.485 29.075 -16.155 29.405 ;
        RECT -16.485 27.715 -16.155 28.045 ;
        RECT -16.485 26.355 -16.155 26.685 ;
        RECT -16.485 24.995 -16.155 25.325 ;
        RECT -16.485 23.635 -16.155 23.965 ;
        RECT -16.485 22.275 -16.155 22.605 ;
        RECT -16.485 20.915 -16.155 21.245 ;
        RECT -16.485 19.555 -16.155 19.885 ;
        RECT -16.485 18.195 -16.155 18.525 ;
        RECT -16.485 16.835 -16.155 17.165 ;
        RECT -16.485 15.475 -16.155 15.805 ;
        RECT -16.485 14.115 -16.155 14.445 ;
        RECT -16.485 12.755 -16.155 13.085 ;
        RECT -16.485 11.395 -16.155 11.725 ;
        RECT -16.485 10.035 -16.155 10.365 ;
        RECT -16.485 8.675 -16.155 9.005 ;
        RECT -16.485 7.315 -16.155 7.645 ;
        RECT -16.485 5.955 -16.155 6.285 ;
        RECT -16.485 4.595 -16.155 4.925 ;
        RECT -16.485 3.235 -16.155 3.565 ;
        RECT -16.485 1.875 -16.155 2.205 ;
        RECT -16.485 0.515 -16.155 0.845 ;
        RECT -16.485 -0.845 -16.155 -0.515 ;
        RECT -16.485 -2.205 -16.155 -1.875 ;
        RECT -16.485 -3.565 -16.155 -3.235 ;
        RECT -16.485 -6.94 -16.155 -6.61 ;
        RECT -16.485 -7.645 -16.155 -7.315 ;
        RECT -16.485 -9.005 -16.155 -8.675 ;
        RECT -16.485 -13.085 -16.155 -12.755 ;
        RECT -16.485 -14.13 -16.155 -13.8 ;
        RECT -16.485 -17.165 -16.155 -16.835 ;
        RECT -16.485 -21.245 -16.155 -20.915 ;
        RECT -16.485 -22.605 -16.155 -22.275 ;
        RECT -16.485 -23.965 -16.155 -23.635 ;
        RECT -16.485 -26.685 -16.155 -26.355 ;
        RECT -16.485 -28.12 -16.155 -27.79 ;
        RECT -16.485 -29.405 -16.155 -29.075 ;
        RECT -16.485 -30.765 -16.155 -30.435 ;
        RECT -16.485 -33.485 -16.155 -33.155 ;
        RECT -16.485 -35.31 -16.155 -34.98 ;
        RECT -16.485 -36.205 -16.155 -35.875 ;
        RECT -16.485 -43.005 -16.155 -42.675 ;
        RECT -16.485 -44.365 -16.155 -44.035 ;
        RECT -16.485 -45.725 -16.155 -45.395 ;
        RECT -16.485 -47.085 -16.155 -46.755 ;
        RECT -16.485 -48.445 -16.155 -48.115 ;
        RECT -16.485 -49.805 -16.155 -49.475 ;
        RECT -16.485 -51.165 -16.155 -50.835 ;
        RECT -16.485 -52.15 -16.155 -51.82 ;
        RECT -16.485 -53.885 -16.155 -53.555 ;
        RECT -16.485 -55.245 -16.155 -54.915 ;
        RECT -16.485 -56.605 -16.155 -56.275 ;
        RECT -16.485 -57.965 -16.155 -57.635 ;
        RECT -16.485 -59.325 -16.155 -58.995 ;
        RECT -16.485 -60.685 -16.155 -60.355 ;
        RECT -16.485 -64.765 -16.155 -64.435 ;
        RECT -16.485 -66.125 -16.155 -65.795 ;
        RECT -16.485 -67.485 -16.155 -67.155 ;
        RECT -16.485 -68.845 -16.155 -68.515 ;
        RECT -16.485 -70.69 -16.155 -70.36 ;
        RECT -16.485 -71.565 -16.155 -71.235 ;
        RECT -16.485 -72.925 -16.155 -72.595 ;
        RECT -16.485 -74.285 -16.155 -73.955 ;
        RECT -16.485 -75.645 -16.155 -75.315 ;
        RECT -16.485 -77.005 -16.155 -76.675 ;
        RECT -16.485 -78.365 -16.155 -78.035 ;
        RECT -16.485 -81.085 -16.155 -80.755 ;
        RECT -16.485 -82.445 -16.155 -82.115 ;
        RECT -16.485 -83.805 -16.155 -83.475 ;
        RECT -16.485 -85.165 -16.155 -84.835 ;
        RECT -16.485 -87.885 -16.155 -87.555 ;
        RECT -16.485 -89.245 -16.155 -88.915 ;
        RECT -16.485 -90.605 -16.155 -90.275 ;
        RECT -16.485 -91.965 -16.155 -91.635 ;
        RECT -16.485 -93.325 -16.155 -92.995 ;
        RECT -16.485 -94.685 -16.155 -94.355 ;
        RECT -16.485 -96.33 -16.155 -96 ;
        RECT -16.485 -97.405 -16.155 -97.075 ;
        RECT -16.485 -98.765 -16.155 -98.435 ;
        RECT -16.485 -100.125 -16.155 -99.795 ;
        RECT -16.485 -101.485 -16.155 -101.155 ;
        RECT -16.485 -102.845 -16.155 -102.515 ;
        RECT -16.485 -104.205 -16.155 -103.875 ;
        RECT -16.485 -106.925 -16.155 -106.595 ;
        RECT -16.485 -108.285 -16.155 -107.955 ;
        RECT -16.485 -109.645 -16.155 -109.315 ;
        RECT -16.485 -111.005 -16.155 -110.675 ;
        RECT -16.485 -113.725 -16.155 -113.395 ;
        RECT -16.485 -114.87 -16.155 -114.54 ;
        RECT -16.485 -116.445 -16.155 -116.115 ;
        RECT -16.485 -117.805 -16.155 -117.475 ;
        RECT -16.485 -119.165 -16.155 -118.835 ;
        RECT -16.485 -120.525 -16.155 -120.195 ;
        RECT -16.485 -121.885 -16.155 -121.555 ;
        RECT -16.485 -123.245 -16.155 -122.915 ;
        RECT -16.485 -125.965 -16.155 -125.635 ;
        RECT -16.485 -127.325 -16.155 -126.995 ;
        RECT -16.485 -128.685 -16.155 -128.355 ;
        RECT -16.48 -130.72 -16.16 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -16.485 -211.645 -16.155 -211.315 ;
        RECT -16.485 -214.365 -16.155 -214.035 ;
        RECT -16.485 -215.725 -16.155 -215.395 ;
        RECT -16.485 -217.085 -16.155 -216.755 ;
        RECT -16.485 -218.445 -16.155 -218.115 ;
        RECT -16.485 -224.09 -16.155 -222.96 ;
        RECT -16.48 -224.205 -16.16 -210.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.125 132.52 -14.795 133.65 ;
        RECT -15.125 128.355 -14.795 128.685 ;
        RECT -15.125 126.995 -14.795 127.325 ;
        RECT -15.125 125.635 -14.795 125.965 ;
        RECT -15.125 124.275 -14.795 124.605 ;
        RECT -15.125 122.915 -14.795 123.245 ;
        RECT -15.125 121.555 -14.795 121.885 ;
        RECT -15.125 120.195 -14.795 120.525 ;
        RECT -15.125 118.835 -14.795 119.165 ;
        RECT -15.125 117.475 -14.795 117.805 ;
        RECT -15.125 116.115 -14.795 116.445 ;
        RECT -15.125 114.755 -14.795 115.085 ;
        RECT -15.125 113.395 -14.795 113.725 ;
        RECT -15.125 112.035 -14.795 112.365 ;
        RECT -15.125 110.675 -14.795 111.005 ;
        RECT -15.125 109.315 -14.795 109.645 ;
        RECT -15.125 107.955 -14.795 108.285 ;
        RECT -15.125 106.595 -14.795 106.925 ;
        RECT -15.125 105.235 -14.795 105.565 ;
        RECT -15.125 103.875 -14.795 104.205 ;
        RECT -15.125 102.515 -14.795 102.845 ;
        RECT -15.125 101.155 -14.795 101.485 ;
        RECT -15.125 99.795 -14.795 100.125 ;
        RECT -15.125 98.435 -14.795 98.765 ;
        RECT -15.125 97.075 -14.795 97.405 ;
        RECT -15.125 95.715 -14.795 96.045 ;
        RECT -15.125 94.355 -14.795 94.685 ;
        RECT -15.125 92.995 -14.795 93.325 ;
        RECT -15.125 91.635 -14.795 91.965 ;
        RECT -15.125 90.275 -14.795 90.605 ;
        RECT -15.125 88.915 -14.795 89.245 ;
        RECT -15.125 87.555 -14.795 87.885 ;
        RECT -15.125 86.195 -14.795 86.525 ;
        RECT -15.125 84.835 -14.795 85.165 ;
        RECT -15.125 83.475 -14.795 83.805 ;
        RECT -15.125 82.115 -14.795 82.445 ;
        RECT -15.125 80.755 -14.795 81.085 ;
        RECT -15.125 79.395 -14.795 79.725 ;
        RECT -15.125 78.035 -14.795 78.365 ;
        RECT -15.125 76.675 -14.795 77.005 ;
        RECT -15.125 75.315 -14.795 75.645 ;
        RECT -15.125 73.955 -14.795 74.285 ;
        RECT -15.125 72.595 -14.795 72.925 ;
        RECT -15.125 71.235 -14.795 71.565 ;
        RECT -15.125 69.875 -14.795 70.205 ;
        RECT -15.125 68.515 -14.795 68.845 ;
        RECT -15.125 67.155 -14.795 67.485 ;
        RECT -15.125 65.795 -14.795 66.125 ;
        RECT -15.125 64.435 -14.795 64.765 ;
        RECT -15.125 63.075 -14.795 63.405 ;
        RECT -15.125 61.715 -14.795 62.045 ;
        RECT -15.125 60.355 -14.795 60.685 ;
        RECT -15.125 58.995 -14.795 59.325 ;
        RECT -15.125 57.635 -14.795 57.965 ;
        RECT -15.125 56.275 -14.795 56.605 ;
        RECT -15.125 54.915 -14.795 55.245 ;
        RECT -15.125 53.555 -14.795 53.885 ;
        RECT -15.125 52.195 -14.795 52.525 ;
        RECT -15.125 50.835 -14.795 51.165 ;
        RECT -15.125 49.475 -14.795 49.805 ;
        RECT -15.125 48.115 -14.795 48.445 ;
        RECT -15.125 46.755 -14.795 47.085 ;
        RECT -15.125 45.395 -14.795 45.725 ;
        RECT -15.125 44.035 -14.795 44.365 ;
        RECT -15.125 42.675 -14.795 43.005 ;
        RECT -15.125 41.315 -14.795 41.645 ;
        RECT -15.125 39.955 -14.795 40.285 ;
        RECT -15.125 38.595 -14.795 38.925 ;
        RECT -15.125 37.235 -14.795 37.565 ;
        RECT -15.125 35.875 -14.795 36.205 ;
        RECT -15.125 34.515 -14.795 34.845 ;
        RECT -15.125 33.155 -14.795 33.485 ;
        RECT -15.125 31.795 -14.795 32.125 ;
        RECT -15.125 30.435 -14.795 30.765 ;
        RECT -15.125 29.075 -14.795 29.405 ;
        RECT -15.125 27.715 -14.795 28.045 ;
        RECT -15.125 26.355 -14.795 26.685 ;
        RECT -15.125 24.995 -14.795 25.325 ;
        RECT -15.125 23.635 -14.795 23.965 ;
        RECT -15.125 22.275 -14.795 22.605 ;
        RECT -15.125 20.915 -14.795 21.245 ;
        RECT -15.125 19.555 -14.795 19.885 ;
        RECT -15.125 18.195 -14.795 18.525 ;
        RECT -15.125 16.835 -14.795 17.165 ;
        RECT -15.125 15.475 -14.795 15.805 ;
        RECT -15.125 14.115 -14.795 14.445 ;
        RECT -15.125 12.755 -14.795 13.085 ;
        RECT -15.125 11.395 -14.795 11.725 ;
        RECT -15.125 10.035 -14.795 10.365 ;
        RECT -15.125 8.675 -14.795 9.005 ;
        RECT -15.125 7.315 -14.795 7.645 ;
        RECT -15.125 5.955 -14.795 6.285 ;
        RECT -15.125 4.595 -14.795 4.925 ;
        RECT -15.125 3.235 -14.795 3.565 ;
        RECT -15.125 1.875 -14.795 2.205 ;
        RECT -15.125 0.515 -14.795 0.845 ;
        RECT -15.125 -0.845 -14.795 -0.515 ;
        RECT -15.125 -2.205 -14.795 -1.875 ;
        RECT -15.125 -3.565 -14.795 -3.235 ;
        RECT -15.125 -6.94 -14.795 -6.61 ;
        RECT -15.125 -7.645 -14.795 -7.315 ;
        RECT -15.125 -9.005 -14.795 -8.675 ;
        RECT -15.125 -13.085 -14.795 -12.755 ;
        RECT -15.125 -14.13 -14.795 -13.8 ;
        RECT -15.125 -17.165 -14.795 -16.835 ;
        RECT -15.125 -21.245 -14.795 -20.915 ;
        RECT -15.125 -22.605 -14.795 -22.275 ;
        RECT -15.125 -23.965 -14.795 -23.635 ;
        RECT -15.125 -26.685 -14.795 -26.355 ;
        RECT -15.125 -28.12 -14.795 -27.79 ;
        RECT -15.125 -29.405 -14.795 -29.075 ;
        RECT -15.125 -30.765 -14.795 -30.435 ;
        RECT -15.125 -33.485 -14.795 -33.155 ;
        RECT -15.125 -35.31 -14.795 -34.98 ;
        RECT -15.125 -36.205 -14.795 -35.875 ;
        RECT -15.125 -43.005 -14.795 -42.675 ;
        RECT -15.125 -44.365 -14.795 -44.035 ;
        RECT -15.125 -45.725 -14.795 -45.395 ;
        RECT -15.125 -47.085 -14.795 -46.755 ;
        RECT -15.125 -48.445 -14.795 -48.115 ;
        RECT -15.125 -49.805 -14.795 -49.475 ;
        RECT -15.125 -51.165 -14.795 -50.835 ;
        RECT -15.125 -52.15 -14.795 -51.82 ;
        RECT -15.125 -53.885 -14.795 -53.555 ;
        RECT -15.125 -55.245 -14.795 -54.915 ;
        RECT -15.125 -56.605 -14.795 -56.275 ;
        RECT -15.125 -57.965 -14.795 -57.635 ;
        RECT -15.125 -59.325 -14.795 -58.995 ;
        RECT -15.125 -60.685 -14.795 -60.355 ;
        RECT -15.125 -64.765 -14.795 -64.435 ;
        RECT -15.125 -66.125 -14.795 -65.795 ;
        RECT -15.125 -67.485 -14.795 -67.155 ;
        RECT -15.125 -68.845 -14.795 -68.515 ;
        RECT -15.125 -70.69 -14.795 -70.36 ;
        RECT -15.125 -71.565 -14.795 -71.235 ;
        RECT -15.125 -72.925 -14.795 -72.595 ;
        RECT -15.125 -74.285 -14.795 -73.955 ;
        RECT -15.125 -75.645 -14.795 -75.315 ;
        RECT -15.125 -77.005 -14.795 -76.675 ;
        RECT -15.125 -78.365 -14.795 -78.035 ;
        RECT -15.125 -81.085 -14.795 -80.755 ;
        RECT -15.125 -82.445 -14.795 -82.115 ;
        RECT -15.125 -83.805 -14.795 -83.475 ;
        RECT -15.125 -85.165 -14.795 -84.835 ;
        RECT -15.125 -87.885 -14.795 -87.555 ;
        RECT -15.125 -89.245 -14.795 -88.915 ;
        RECT -15.125 -90.605 -14.795 -90.275 ;
        RECT -15.125 -91.965 -14.795 -91.635 ;
        RECT -15.125 -93.325 -14.795 -92.995 ;
        RECT -15.125 -94.685 -14.795 -94.355 ;
        RECT -15.125 -96.33 -14.795 -96 ;
        RECT -15.125 -97.405 -14.795 -97.075 ;
        RECT -15.125 -98.765 -14.795 -98.435 ;
        RECT -15.125 -100.125 -14.795 -99.795 ;
        RECT -15.125 -101.485 -14.795 -101.155 ;
        RECT -15.125 -102.845 -14.795 -102.515 ;
        RECT -15.125 -104.205 -14.795 -103.875 ;
        RECT -15.125 -106.925 -14.795 -106.595 ;
        RECT -15.125 -108.285 -14.795 -107.955 ;
        RECT -15.125 -109.645 -14.795 -109.315 ;
        RECT -15.125 -111.005 -14.795 -110.675 ;
        RECT -15.125 -113.725 -14.795 -113.395 ;
        RECT -15.125 -114.87 -14.795 -114.54 ;
        RECT -15.125 -116.445 -14.795 -116.115 ;
        RECT -15.125 -117.805 -14.795 -117.475 ;
        RECT -15.125 -119.165 -14.795 -118.835 ;
        RECT -15.125 -120.525 -14.795 -120.195 ;
        RECT -15.125 -121.885 -14.795 -121.555 ;
        RECT -15.125 -123.245 -14.795 -122.915 ;
        RECT -15.125 -125.965 -14.795 -125.635 ;
        RECT -15.125 -127.325 -14.795 -126.995 ;
        RECT -15.125 -128.685 -14.795 -128.355 ;
        RECT -15.12 -129.36 -14.8 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -13.765 132.52 -13.435 133.65 ;
        RECT -13.765 128.355 -13.435 128.685 ;
        RECT -13.765 126.995 -13.435 127.325 ;
        RECT -13.765 125.635 -13.435 125.965 ;
        RECT -13.765 124.275 -13.435 124.605 ;
        RECT -13.765 122.915 -13.435 123.245 ;
        RECT -13.765 121.555 -13.435 121.885 ;
        RECT -13.765 120.195 -13.435 120.525 ;
        RECT -13.765 118.835 -13.435 119.165 ;
        RECT -13.765 117.475 -13.435 117.805 ;
        RECT -13.765 116.115 -13.435 116.445 ;
        RECT -13.765 114.755 -13.435 115.085 ;
        RECT -13.765 113.395 -13.435 113.725 ;
        RECT -13.765 112.035 -13.435 112.365 ;
        RECT -13.765 110.675 -13.435 111.005 ;
        RECT -13.765 109.315 -13.435 109.645 ;
        RECT -13.765 107.955 -13.435 108.285 ;
        RECT -13.765 106.595 -13.435 106.925 ;
        RECT -13.765 105.235 -13.435 105.565 ;
        RECT -13.765 103.875 -13.435 104.205 ;
        RECT -13.765 102.515 -13.435 102.845 ;
        RECT -13.765 101.155 -13.435 101.485 ;
        RECT -13.765 99.795 -13.435 100.125 ;
        RECT -13.765 98.435 -13.435 98.765 ;
        RECT -13.765 97.075 -13.435 97.405 ;
        RECT -13.765 95.715 -13.435 96.045 ;
        RECT -13.765 94.355 -13.435 94.685 ;
        RECT -13.765 92.995 -13.435 93.325 ;
        RECT -13.765 91.635 -13.435 91.965 ;
        RECT -13.765 90.275 -13.435 90.605 ;
        RECT -13.765 88.915 -13.435 89.245 ;
        RECT -13.765 87.555 -13.435 87.885 ;
        RECT -13.765 86.195 -13.435 86.525 ;
        RECT -13.765 84.835 -13.435 85.165 ;
        RECT -13.765 83.475 -13.435 83.805 ;
        RECT -13.765 82.115 -13.435 82.445 ;
        RECT -13.765 80.755 -13.435 81.085 ;
        RECT -13.765 79.395 -13.435 79.725 ;
        RECT -13.765 78.035 -13.435 78.365 ;
        RECT -13.765 76.675 -13.435 77.005 ;
        RECT -13.765 75.315 -13.435 75.645 ;
        RECT -13.765 73.955 -13.435 74.285 ;
        RECT -13.765 72.595 -13.435 72.925 ;
        RECT -13.765 71.235 -13.435 71.565 ;
        RECT -13.765 69.875 -13.435 70.205 ;
        RECT -13.765 68.515 -13.435 68.845 ;
        RECT -13.765 67.155 -13.435 67.485 ;
        RECT -13.765 65.795 -13.435 66.125 ;
        RECT -13.765 64.435 -13.435 64.765 ;
        RECT -13.765 63.075 -13.435 63.405 ;
        RECT -13.765 61.715 -13.435 62.045 ;
        RECT -13.765 60.355 -13.435 60.685 ;
        RECT -13.765 58.995 -13.435 59.325 ;
        RECT -13.765 57.635 -13.435 57.965 ;
        RECT -13.765 56.275 -13.435 56.605 ;
        RECT -13.765 54.915 -13.435 55.245 ;
        RECT -13.765 53.555 -13.435 53.885 ;
        RECT -13.765 52.195 -13.435 52.525 ;
        RECT -13.765 50.835 -13.435 51.165 ;
        RECT -13.765 49.475 -13.435 49.805 ;
        RECT -13.765 48.115 -13.435 48.445 ;
        RECT -13.765 46.755 -13.435 47.085 ;
        RECT -13.765 45.395 -13.435 45.725 ;
        RECT -13.765 44.035 -13.435 44.365 ;
        RECT -13.765 42.675 -13.435 43.005 ;
        RECT -13.765 41.315 -13.435 41.645 ;
        RECT -13.765 39.955 -13.435 40.285 ;
        RECT -13.765 38.595 -13.435 38.925 ;
        RECT -13.765 37.235 -13.435 37.565 ;
        RECT -13.765 35.875 -13.435 36.205 ;
        RECT -13.765 34.515 -13.435 34.845 ;
        RECT -13.765 33.155 -13.435 33.485 ;
        RECT -13.765 31.795 -13.435 32.125 ;
        RECT -13.765 30.435 -13.435 30.765 ;
        RECT -13.765 29.075 -13.435 29.405 ;
        RECT -13.765 27.715 -13.435 28.045 ;
        RECT -13.765 26.355 -13.435 26.685 ;
        RECT -13.765 24.995 -13.435 25.325 ;
        RECT -13.765 23.635 -13.435 23.965 ;
        RECT -13.765 22.275 -13.435 22.605 ;
        RECT -13.765 20.915 -13.435 21.245 ;
        RECT -13.765 19.555 -13.435 19.885 ;
        RECT -13.765 18.195 -13.435 18.525 ;
        RECT -13.765 16.835 -13.435 17.165 ;
        RECT -13.765 15.475 -13.435 15.805 ;
        RECT -13.765 14.115 -13.435 14.445 ;
        RECT -13.765 12.755 -13.435 13.085 ;
        RECT -13.765 11.395 -13.435 11.725 ;
        RECT -13.765 10.035 -13.435 10.365 ;
        RECT -13.765 8.675 -13.435 9.005 ;
        RECT -13.765 7.315 -13.435 7.645 ;
        RECT -13.765 5.955 -13.435 6.285 ;
        RECT -13.765 4.595 -13.435 4.925 ;
        RECT -13.765 3.235 -13.435 3.565 ;
        RECT -13.765 1.875 -13.435 2.205 ;
        RECT -13.765 0.515 -13.435 0.845 ;
        RECT -13.765 -0.845 -13.435 -0.515 ;
        RECT -13.765 -2.205 -13.435 -1.875 ;
        RECT -13.765 -3.565 -13.435 -3.235 ;
        RECT -13.765 -6.94 -13.435 -6.61 ;
        RECT -13.765 -7.645 -13.435 -7.315 ;
        RECT -13.765 -9.005 -13.435 -8.675 ;
        RECT -13.765 -13.085 -13.435 -12.755 ;
        RECT -13.765 -14.13 -13.435 -13.8 ;
        RECT -13.765 -17.165 -13.435 -16.835 ;
        RECT -13.765 -21.245 -13.435 -20.915 ;
        RECT -13.765 -22.605 -13.435 -22.275 ;
        RECT -13.765 -23.965 -13.435 -23.635 ;
        RECT -13.765 -26.685 -13.435 -26.355 ;
        RECT -13.765 -28.12 -13.435 -27.79 ;
        RECT -13.765 -29.405 -13.435 -29.075 ;
        RECT -13.765 -30.765 -13.435 -30.435 ;
        RECT -13.765 -33.485 -13.435 -33.155 ;
        RECT -13.765 -35.31 -13.435 -34.98 ;
        RECT -13.765 -36.205 -13.435 -35.875 ;
        RECT -13.765 -43.005 -13.435 -42.675 ;
        RECT -13.765 -44.365 -13.435 -44.035 ;
        RECT -13.765 -45.725 -13.435 -45.395 ;
        RECT -13.765 -47.085 -13.435 -46.755 ;
        RECT -13.765 -48.445 -13.435 -48.115 ;
        RECT -13.765 -49.805 -13.435 -49.475 ;
        RECT -13.765 -51.165 -13.435 -50.835 ;
        RECT -13.765 -52.15 -13.435 -51.82 ;
        RECT -13.765 -53.885 -13.435 -53.555 ;
        RECT -13.765 -55.245 -13.435 -54.915 ;
        RECT -13.765 -56.605 -13.435 -56.275 ;
        RECT -13.765 -57.965 -13.435 -57.635 ;
        RECT -13.765 -59.325 -13.435 -58.995 ;
        RECT -13.765 -60.685 -13.435 -60.355 ;
        RECT -13.765 -64.765 -13.435 -64.435 ;
        RECT -13.765 -66.125 -13.435 -65.795 ;
        RECT -13.76 -66.8 -13.44 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -13.765 -145.005 -13.435 -144.675 ;
        RECT -13.765 -147.725 -13.435 -147.395 ;
        RECT -13.765 -149.085 -13.435 -148.755 ;
        RECT -13.765 -150.445 -13.435 -150.115 ;
        RECT -13.765 -151.805 -13.435 -151.475 ;
        RECT -13.765 -155.885 -13.435 -155.555 ;
        RECT -13.765 -157.245 -13.435 -156.915 ;
        RECT -13.765 -158.605 -13.435 -158.275 ;
        RECT -13.765 -159.965 -13.435 -159.635 ;
        RECT -13.765 -161.325 -13.435 -160.995 ;
        RECT -13.765 -162.685 -13.435 -162.355 ;
        RECT -13.765 -169.485 -13.435 -169.155 ;
        RECT -13.765 -170.845 -13.435 -170.515 ;
        RECT -13.765 -172.205 -13.435 -171.875 ;
        RECT -13.765 -174.925 -13.435 -174.595 ;
        RECT -13.765 -176.285 -13.435 -175.955 ;
        RECT -13.765 -177.645 -13.435 -177.315 ;
        RECT -13.765 -179.005 -13.435 -178.675 ;
        RECT -13.765 -184.445 -13.435 -184.115 ;
        RECT -13.765 -187.165 -13.435 -186.835 ;
        RECT -13.765 -189.885 -13.435 -189.555 ;
        RECT -13.765 -192.605 -13.435 -192.275 ;
        RECT -13.765 -195.325 -13.435 -194.995 ;
        RECT -13.765 -196.685 -13.435 -196.355 ;
        RECT -13.765 -198.045 -13.435 -197.715 ;
        RECT -13.765 -199.405 -13.435 -199.075 ;
        RECT -13.765 -200.765 -13.435 -200.435 ;
        RECT -13.765 -202.125 -13.435 -201.795 ;
        RECT -13.765 -203.485 -13.435 -203.155 ;
        RECT -13.765 -206.555 -13.435 -206.225 ;
        RECT -13.765 -207.565 -13.435 -207.235 ;
        RECT -13.765 -208.925 -13.435 -208.595 ;
        RECT -13.765 -211.645 -13.435 -211.315 ;
        RECT -13.765 -214.365 -13.435 -214.035 ;
        RECT -13.765 -215.725 -13.435 -215.395 ;
        RECT -13.765 -217.085 -13.435 -216.755 ;
        RECT -13.765 -218.445 -13.435 -218.115 ;
        RECT -13.765 -224.09 -13.435 -222.96 ;
        RECT -13.76 -224.205 -13.44 -141.96 ;
    END
    PORT
      LAYER met3 ;
        RECT -12.405 132.52 -12.075 133.65 ;
        RECT -12.405 128.355 -12.075 128.685 ;
        RECT -12.405 126.995 -12.075 127.325 ;
        RECT -12.405 125.635 -12.075 125.965 ;
        RECT -12.405 124.275 -12.075 124.605 ;
        RECT -12.405 122.915 -12.075 123.245 ;
        RECT -12.405 121.555 -12.075 121.885 ;
        RECT -12.405 120.195 -12.075 120.525 ;
        RECT -12.405 118.835 -12.075 119.165 ;
        RECT -12.405 117.475 -12.075 117.805 ;
        RECT -12.405 116.115 -12.075 116.445 ;
        RECT -12.405 114.755 -12.075 115.085 ;
        RECT -12.405 113.395 -12.075 113.725 ;
        RECT -12.405 112.035 -12.075 112.365 ;
        RECT -12.405 110.675 -12.075 111.005 ;
        RECT -12.405 109.315 -12.075 109.645 ;
        RECT -12.405 107.955 -12.075 108.285 ;
        RECT -12.405 106.595 -12.075 106.925 ;
        RECT -12.405 105.235 -12.075 105.565 ;
        RECT -12.405 103.875 -12.075 104.205 ;
        RECT -12.405 102.515 -12.075 102.845 ;
        RECT -12.405 101.155 -12.075 101.485 ;
        RECT -12.405 99.795 -12.075 100.125 ;
        RECT -12.405 98.435 -12.075 98.765 ;
        RECT -12.405 97.075 -12.075 97.405 ;
        RECT -12.405 95.715 -12.075 96.045 ;
        RECT -12.405 94.355 -12.075 94.685 ;
        RECT -12.405 92.995 -12.075 93.325 ;
        RECT -12.405 91.635 -12.075 91.965 ;
        RECT -12.405 90.275 -12.075 90.605 ;
        RECT -12.405 88.915 -12.075 89.245 ;
        RECT -12.405 87.555 -12.075 87.885 ;
        RECT -12.405 86.195 -12.075 86.525 ;
        RECT -12.405 84.835 -12.075 85.165 ;
        RECT -12.405 83.475 -12.075 83.805 ;
        RECT -12.405 82.115 -12.075 82.445 ;
        RECT -12.405 80.755 -12.075 81.085 ;
        RECT -12.405 79.395 -12.075 79.725 ;
        RECT -12.405 78.035 -12.075 78.365 ;
        RECT -12.405 76.675 -12.075 77.005 ;
        RECT -12.405 75.315 -12.075 75.645 ;
        RECT -12.405 73.955 -12.075 74.285 ;
        RECT -12.405 72.595 -12.075 72.925 ;
        RECT -12.405 71.235 -12.075 71.565 ;
        RECT -12.405 69.875 -12.075 70.205 ;
        RECT -12.405 68.515 -12.075 68.845 ;
        RECT -12.405 67.155 -12.075 67.485 ;
        RECT -12.405 65.795 -12.075 66.125 ;
        RECT -12.405 64.435 -12.075 64.765 ;
        RECT -12.405 63.075 -12.075 63.405 ;
        RECT -12.405 61.715 -12.075 62.045 ;
        RECT -12.405 60.355 -12.075 60.685 ;
        RECT -12.405 58.995 -12.075 59.325 ;
        RECT -12.405 57.635 -12.075 57.965 ;
        RECT -12.405 56.275 -12.075 56.605 ;
        RECT -12.405 54.915 -12.075 55.245 ;
        RECT -12.405 53.555 -12.075 53.885 ;
        RECT -12.405 52.195 -12.075 52.525 ;
        RECT -12.405 50.835 -12.075 51.165 ;
        RECT -12.405 49.475 -12.075 49.805 ;
        RECT -12.405 48.115 -12.075 48.445 ;
        RECT -12.405 46.755 -12.075 47.085 ;
        RECT -12.405 45.395 -12.075 45.725 ;
        RECT -12.405 44.035 -12.075 44.365 ;
        RECT -12.405 42.675 -12.075 43.005 ;
        RECT -12.405 41.315 -12.075 41.645 ;
        RECT -12.405 39.955 -12.075 40.285 ;
        RECT -12.405 38.595 -12.075 38.925 ;
        RECT -12.405 37.235 -12.075 37.565 ;
        RECT -12.405 35.875 -12.075 36.205 ;
        RECT -12.405 34.515 -12.075 34.845 ;
        RECT -12.405 33.155 -12.075 33.485 ;
        RECT -12.405 31.795 -12.075 32.125 ;
        RECT -12.405 30.435 -12.075 30.765 ;
        RECT -12.405 29.075 -12.075 29.405 ;
        RECT -12.405 27.715 -12.075 28.045 ;
        RECT -12.405 26.355 -12.075 26.685 ;
        RECT -12.405 24.995 -12.075 25.325 ;
        RECT -12.405 23.635 -12.075 23.965 ;
        RECT -12.405 22.275 -12.075 22.605 ;
        RECT -12.405 20.915 -12.075 21.245 ;
        RECT -12.405 19.555 -12.075 19.885 ;
        RECT -12.405 18.195 -12.075 18.525 ;
        RECT -12.405 16.835 -12.075 17.165 ;
        RECT -12.405 15.475 -12.075 15.805 ;
        RECT -12.405 14.115 -12.075 14.445 ;
        RECT -12.405 12.755 -12.075 13.085 ;
        RECT -12.405 11.395 -12.075 11.725 ;
        RECT -12.405 10.035 -12.075 10.365 ;
        RECT -12.405 8.675 -12.075 9.005 ;
        RECT -12.405 7.315 -12.075 7.645 ;
        RECT -12.405 5.955 -12.075 6.285 ;
        RECT -12.405 4.595 -12.075 4.925 ;
        RECT -12.405 3.235 -12.075 3.565 ;
        RECT -12.405 1.875 -12.075 2.205 ;
        RECT -12.405 0.515 -12.075 0.845 ;
        RECT -12.405 -0.845 -12.075 -0.515 ;
        RECT -12.405 -2.205 -12.075 -1.875 ;
        RECT -12.405 -3.565 -12.075 -3.235 ;
        RECT -12.405 -4.925 -12.075 -4.595 ;
        RECT -12.405 -6.94 -12.075 -6.61 ;
        RECT -12.405 -7.645 -12.075 -7.315 ;
        RECT -12.405 -9.005 -12.075 -8.675 ;
        RECT -12.405 -13.085 -12.075 -12.755 ;
        RECT -12.405 -14.13 -12.075 -13.8 ;
        RECT -12.405 -17.165 -12.075 -16.835 ;
        RECT -12.405 -21.245 -12.075 -20.915 ;
        RECT -12.405 -22.605 -12.075 -22.275 ;
        RECT -12.405 -23.965 -12.075 -23.635 ;
        RECT -12.405 -25.325 -12.075 -24.995 ;
        RECT -12.405 -26.685 -12.075 -26.355 ;
        RECT -12.405 -28.12 -12.075 -27.79 ;
        RECT -12.405 -29.405 -12.075 -29.075 ;
        RECT -12.405 -30.765 -12.075 -30.435 ;
        RECT -12.405 -33.485 -12.075 -33.155 ;
        RECT -12.405 -35.31 -12.075 -34.98 ;
        RECT -12.405 -36.205 -12.075 -35.875 ;
        RECT -12.405 -43.005 -12.075 -42.675 ;
        RECT -12.405 -44.365 -12.075 -44.035 ;
        RECT -12.405 -45.725 -12.075 -45.395 ;
        RECT -12.405 -47.085 -12.075 -46.755 ;
        RECT -12.405 -48.445 -12.075 -48.115 ;
        RECT -12.405 -49.805 -12.075 -49.475 ;
        RECT -12.405 -51.165 -12.075 -50.835 ;
        RECT -12.405 -52.15 -12.075 -51.82 ;
        RECT -12.405 -53.885 -12.075 -53.555 ;
        RECT -12.405 -55.245 -12.075 -54.915 ;
        RECT -12.405 -56.605 -12.075 -56.275 ;
        RECT -12.405 -57.965 -12.075 -57.635 ;
        RECT -12.405 -59.325 -12.075 -58.995 ;
        RECT -12.405 -66.125 -12.075 -65.795 ;
        RECT -12.405 -68.845 -12.075 -68.515 ;
        RECT -12.405 -70.69 -12.075 -70.36 ;
        RECT -12.405 -71.565 -12.075 -71.235 ;
        RECT -12.405 -72.925 -12.075 -72.595 ;
        RECT -12.405 -74.285 -12.075 -73.955 ;
        RECT -12.405 -75.645 -12.075 -75.315 ;
        RECT -12.405 -77.005 -12.075 -76.675 ;
        RECT -12.405 -78.365 -12.075 -78.035 ;
        RECT -12.405 -81.085 -12.075 -80.755 ;
        RECT -12.405 -82.445 -12.075 -82.115 ;
        RECT -12.405 -83.805 -12.075 -83.475 ;
        RECT -12.405 -85.165 -12.075 -84.835 ;
        RECT -12.405 -87.885 -12.075 -87.555 ;
        RECT -12.405 -89.245 -12.075 -88.915 ;
        RECT -12.405 -90.605 -12.075 -90.275 ;
        RECT -12.405 -91.965 -12.075 -91.635 ;
        RECT -12.405 -93.325 -12.075 -92.995 ;
        RECT -12.405 -94.685 -12.075 -94.355 ;
        RECT -12.405 -96.33 -12.075 -96 ;
        RECT -12.405 -97.405 -12.075 -97.075 ;
        RECT -12.405 -98.765 -12.075 -98.435 ;
        RECT -12.405 -100.125 -12.075 -99.795 ;
        RECT -12.405 -101.485 -12.075 -101.155 ;
        RECT -12.405 -102.845 -12.075 -102.515 ;
        RECT -12.405 -104.205 -12.075 -103.875 ;
        RECT -12.405 -106.925 -12.075 -106.595 ;
        RECT -12.405 -108.285 -12.075 -107.955 ;
        RECT -12.405 -109.645 -12.075 -109.315 ;
        RECT -12.405 -111.005 -12.075 -110.675 ;
        RECT -12.4 -113.04 -12.08 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -12.405 -198.045 -12.075 -197.715 ;
        RECT -12.405 -199.405 -12.075 -199.075 ;
        RECT -12.405 -200.765 -12.075 -200.435 ;
        RECT -12.405 -202.125 -12.075 -201.795 ;
        RECT -12.405 -203.485 -12.075 -203.155 ;
        RECT -12.405 -206.555 -12.075 -206.225 ;
        RECT -12.405 -207.565 -12.075 -207.235 ;
        RECT -12.405 -208.925 -12.075 -208.595 ;
        RECT -12.405 -210.285 -12.075 -209.955 ;
        RECT -12.405 -211.645 -12.075 -211.315 ;
        RECT -12.405 -214.365 -12.075 -214.035 ;
        RECT -12.405 -215.725 -12.075 -215.395 ;
        RECT -12.405 -217.085 -12.075 -216.755 ;
        RECT -12.405 -218.445 -12.075 -218.115 ;
        RECT -12.405 -224.09 -12.075 -222.96 ;
        RECT -12.4 -224.205 -12.08 -197.04 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.045 132.52 -10.715 133.65 ;
        RECT -11.045 128.355 -10.715 128.685 ;
        RECT -11.045 126.995 -10.715 127.325 ;
        RECT -11.045 125.635 -10.715 125.965 ;
        RECT -11.045 124.275 -10.715 124.605 ;
        RECT -11.045 122.915 -10.715 123.245 ;
        RECT -11.045 121.555 -10.715 121.885 ;
        RECT -11.045 120.195 -10.715 120.525 ;
        RECT -11.045 118.835 -10.715 119.165 ;
        RECT -11.045 117.475 -10.715 117.805 ;
        RECT -11.045 110.675 -10.715 111.005 ;
        RECT -11.045 107.955 -10.715 108.285 ;
        RECT -11.045 103.875 -10.715 104.205 ;
        RECT -11.045 99.795 -10.715 100.125 ;
        RECT -11.045 97.075 -10.715 97.405 ;
        RECT -11.045 90.275 -10.715 90.605 ;
        RECT -11.045 88.915 -10.715 89.245 ;
        RECT -11.045 82.115 -10.715 82.445 ;
        RECT -11.045 79.395 -10.715 79.725 ;
        RECT -11.045 75.315 -10.715 75.645 ;
        RECT -11.045 71.235 -10.715 71.565 ;
        RECT -11.045 68.515 -10.715 68.845 ;
        RECT -11.045 61.715 -10.715 62.045 ;
        RECT -11.045 60.355 -10.715 60.685 ;
        RECT -11.045 50.835 -10.715 51.165 ;
        RECT -11.045 46.755 -10.715 47.085 ;
        RECT -11.045 42.675 -10.715 43.005 ;
        RECT -11.045 39.955 -10.715 40.285 ;
        RECT -11.045 33.155 -10.715 33.485 ;
        RECT -11.045 31.795 -10.715 32.125 ;
        RECT -11.045 29.075 -10.715 29.405 ;
        RECT -11.045 22.275 -10.715 22.605 ;
        RECT -11.045 19.555 -10.715 19.885 ;
        RECT -11.045 18.195 -10.715 18.525 ;
        RECT -11.045 11.395 -10.715 11.725 ;
        RECT -11.045 4.595 -10.715 4.925 ;
        RECT -11.045 3.235 -10.715 3.565 ;
        RECT -11.045 1.875 -10.715 2.205 ;
        RECT -11.045 0.515 -10.715 0.845 ;
        RECT -11.045 -0.845 -10.715 -0.515 ;
        RECT -11.045 -2.205 -10.715 -1.875 ;
        RECT -11.045 -3.565 -10.715 -3.235 ;
        RECT -11.045 -4.925 -10.715 -4.595 ;
        RECT -11.045 -6.94 -10.715 -6.61 ;
        RECT -11.045 -7.645 -10.715 -7.315 ;
        RECT -11.045 -9.005 -10.715 -8.675 ;
        RECT -11.045 -13.085 -10.715 -12.755 ;
        RECT -11.045 -14.13 -10.715 -13.8 ;
        RECT -11.045 -17.165 -10.715 -16.835 ;
        RECT -11.045 -21.245 -10.715 -20.915 ;
        RECT -11.045 -22.605 -10.715 -22.275 ;
        RECT -11.045 -23.965 -10.715 -23.635 ;
        RECT -11.045 -25.325 -10.715 -24.995 ;
        RECT -11.045 -26.685 -10.715 -26.355 ;
        RECT -11.045 -28.12 -10.715 -27.79 ;
        RECT -11.045 -29.405 -10.715 -29.075 ;
        RECT -11.045 -30.765 -10.715 -30.435 ;
        RECT -11.045 -33.485 -10.715 -33.155 ;
        RECT -11.045 -35.31 -10.715 -34.98 ;
        RECT -11.045 -36.205 -10.715 -35.875 ;
        RECT -11.045 -43.005 -10.715 -42.675 ;
        RECT -11.045 -44.365 -10.715 -44.035 ;
        RECT -11.045 -45.725 -10.715 -45.395 ;
        RECT -11.045 -47.085 -10.715 -46.755 ;
        RECT -11.045 -48.445 -10.715 -48.115 ;
        RECT -11.045 -49.805 -10.715 -49.475 ;
        RECT -11.045 -51.165 -10.715 -50.835 ;
        RECT -11.045 -52.15 -10.715 -51.82 ;
        RECT -11.045 -53.885 -10.715 -53.555 ;
        RECT -11.045 -55.245 -10.715 -54.915 ;
        RECT -11.045 -56.605 -10.715 -56.275 ;
        RECT -11.045 -57.965 -10.715 -57.635 ;
        RECT -11.045 -59.325 -10.715 -58.995 ;
        RECT -11.045 -66.125 -10.715 -65.795 ;
        RECT -11.045 -68.845 -10.715 -68.515 ;
        RECT -11.045 -70.69 -10.715 -70.36 ;
        RECT -11.045 -71.565 -10.715 -71.235 ;
        RECT -11.045 -72.925 -10.715 -72.595 ;
        RECT -11.045 -74.285 -10.715 -73.955 ;
        RECT -11.045 -75.645 -10.715 -75.315 ;
        RECT -11.045 -77.005 -10.715 -76.675 ;
        RECT -11.045 -78.365 -10.715 -78.035 ;
        RECT -11.045 -81.085 -10.715 -80.755 ;
        RECT -11.045 -82.445 -10.715 -82.115 ;
        RECT -11.045 -83.805 -10.715 -83.475 ;
        RECT -11.045 -85.165 -10.715 -84.835 ;
        RECT -11.045 -87.885 -10.715 -87.555 ;
        RECT -11.045 -89.245 -10.715 -88.915 ;
        RECT -11.045 -90.605 -10.715 -90.275 ;
        RECT -11.045 -91.965 -10.715 -91.635 ;
        RECT -11.045 -93.325 -10.715 -92.995 ;
        RECT -11.045 -94.685 -10.715 -94.355 ;
        RECT -11.045 -96.33 -10.715 -96 ;
        RECT -11.045 -97.405 -10.715 -97.075 ;
        RECT -11.045 -98.765 -10.715 -98.435 ;
        RECT -11.045 -100.125 -10.715 -99.795 ;
        RECT -11.045 -101.485 -10.715 -101.155 ;
        RECT -11.045 -102.845 -10.715 -102.515 ;
        RECT -11.045 -104.205 -10.715 -103.875 ;
        RECT -11.045 -106.925 -10.715 -106.595 ;
        RECT -11.045 -108.285 -10.715 -107.955 ;
        RECT -11.045 -109.645 -10.715 -109.315 ;
        RECT -11.045 -111.005 -10.715 -110.675 ;
        RECT -11.045 -114.87 -10.715 -114.54 ;
        RECT -11.045 -116.445 -10.715 -116.115 ;
        RECT -11.045 -117.805 -10.715 -117.475 ;
        RECT -11.045 -119.165 -10.715 -118.835 ;
        RECT -11.045 -120.525 -10.715 -120.195 ;
        RECT -11.045 -121.885 -10.715 -121.555 ;
        RECT -11.045 -123.245 -10.715 -122.915 ;
        RECT -11.045 -125.965 -10.715 -125.635 ;
        RECT -11.045 -127.325 -10.715 -126.995 ;
        RECT -11.045 -128.685 -10.715 -128.355 ;
        RECT -11.045 -132.765 -10.715 -132.435 ;
        RECT -11.045 -134.125 -10.715 -133.795 ;
        RECT -11.045 -135.485 -10.715 -135.155 ;
        RECT -11.045 -136.845 -10.715 -136.515 ;
        RECT -11.045 -138.205 -10.715 -137.875 ;
        RECT -11.045 -140.925 -10.715 -140.595 ;
        RECT -11.045 -142.285 -10.715 -141.955 ;
        RECT -11.045 -145.005 -10.715 -144.675 ;
        RECT -11.045 -147.725 -10.715 -147.395 ;
        RECT -11.045 -149.085 -10.715 -148.755 ;
        RECT -11.045 -151.805 -10.715 -151.475 ;
        RECT -11.045 -153.165 -10.715 -152.835 ;
        RECT -11.045 -154.525 -10.715 -154.195 ;
        RECT -11.045 -155.885 -10.715 -155.555 ;
        RECT -11.045 -157.245 -10.715 -156.915 ;
        RECT -11.045 -158.605 -10.715 -158.275 ;
        RECT -11.045 -159.965 -10.715 -159.635 ;
        RECT -11.045 -161.325 -10.715 -160.995 ;
        RECT -11.045 -162.685 -10.715 -162.355 ;
        RECT -11.045 -164.045 -10.715 -163.715 ;
        RECT -11.045 -165.405 -10.715 -165.075 ;
        RECT -11.045 -166.765 -10.715 -166.435 ;
        RECT -11.045 -168.125 -10.715 -167.795 ;
        RECT -11.045 -169.485 -10.715 -169.155 ;
        RECT -11.045 -170.845 -10.715 -170.515 ;
        RECT -11.045 -172.205 -10.715 -171.875 ;
        RECT -11.045 -173.565 -10.715 -173.235 ;
        RECT -11.045 -174.925 -10.715 -174.595 ;
        RECT -11.045 -176.285 -10.715 -175.955 ;
        RECT -11.045 -177.645 -10.715 -177.315 ;
        RECT -11.045 -179.005 -10.715 -178.675 ;
        RECT -11.045 -181.725 -10.715 -181.395 ;
        RECT -11.045 -184.445 -10.715 -184.115 ;
        RECT -11.045 -185.805 -10.715 -185.475 ;
        RECT -11.045 -187.165 -10.715 -186.835 ;
        RECT -11.045 -188.525 -10.715 -188.195 ;
        RECT -11.045 -189.885 -10.715 -189.555 ;
        RECT -11.045 -191.245 -10.715 -190.915 ;
        RECT -11.045 -192.605 -10.715 -192.275 ;
        RECT -11.045 -193.965 -10.715 -193.635 ;
        RECT -11.045 -195.325 -10.715 -194.995 ;
        RECT -11.045 -196.685 -10.715 -196.355 ;
        RECT -11.045 -198.045 -10.715 -197.715 ;
        RECT -11.045 -199.405 -10.715 -199.075 ;
        RECT -11.045 -200.765 -10.715 -200.435 ;
        RECT -11.045 -202.125 -10.715 -201.795 ;
        RECT -11.045 -203.485 -10.715 -203.155 ;
        RECT -11.045 -206.555 -10.715 -206.225 ;
        RECT -11.045 -207.565 -10.715 -207.235 ;
        RECT -11.045 -208.925 -10.715 -208.595 ;
        RECT -11.045 -214.365 -10.715 -214.035 ;
        RECT -11.045 -215.725 -10.715 -215.395 ;
        RECT -11.045 -217.085 -10.715 -216.755 ;
        RECT -11.045 -218.445 -10.715 -218.115 ;
        RECT -11.045 -224.09 -10.715 -222.96 ;
        RECT -11.04 -224.205 -10.72 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.685 -75.645 -9.355 -75.315 ;
        RECT -9.685 -77.005 -9.355 -76.675 ;
        RECT -9.685 -78.365 -9.355 -78.035 ;
        RECT -9.685 -81.085 -9.355 -80.755 ;
        RECT -9.685 -82.445 -9.355 -82.115 ;
        RECT -9.685 -83.805 -9.355 -83.475 ;
        RECT -9.685 -85.165 -9.355 -84.835 ;
        RECT -9.685 -87.885 -9.355 -87.555 ;
        RECT -9.685 -89.245 -9.355 -88.915 ;
        RECT -9.685 -90.605 -9.355 -90.275 ;
        RECT -9.685 -91.965 -9.355 -91.635 ;
        RECT -9.685 -93.325 -9.355 -92.995 ;
        RECT -9.685 -94.685 -9.355 -94.355 ;
        RECT -9.685 -97.405 -9.355 -97.075 ;
        RECT -9.685 -98.765 -9.355 -98.435 ;
        RECT -9.685 -100.125 -9.355 -99.795 ;
        RECT -9.685 -101.485 -9.355 -101.155 ;
        RECT -9.685 -102.845 -9.355 -102.515 ;
        RECT -9.685 -104.205 -9.355 -103.875 ;
        RECT -9.685 -106.925 -9.355 -106.595 ;
        RECT -9.685 -108.285 -9.355 -107.955 ;
        RECT -9.685 -109.645 -9.355 -109.315 ;
        RECT -9.685 -111.005 -9.355 -110.675 ;
        RECT -9.685 -116.445 -9.355 -116.115 ;
        RECT -9.685 -117.805 -9.355 -117.475 ;
        RECT -9.685 -119.165 -9.355 -118.835 ;
        RECT -9.685 -120.525 -9.355 -120.195 ;
        RECT -9.685 -121.885 -9.355 -121.555 ;
        RECT -9.685 -123.245 -9.355 -122.915 ;
        RECT -9.685 -125.965 -9.355 -125.635 ;
        RECT -9.685 -127.325 -9.355 -126.995 ;
        RECT -9.685 -128.685 -9.355 -128.355 ;
        RECT -9.685 -132.765 -9.355 -132.435 ;
        RECT -9.685 -134.125 -9.355 -133.795 ;
        RECT -9.685 -135.485 -9.355 -135.155 ;
        RECT -9.685 -136.845 -9.355 -136.515 ;
        RECT -9.685 -138.205 -9.355 -137.875 ;
        RECT -9.685 -140.925 -9.355 -140.595 ;
        RECT -9.685 -142.285 -9.355 -141.955 ;
        RECT -9.685 -145.005 -9.355 -144.675 ;
        RECT -9.685 -146.365 -9.355 -146.035 ;
        RECT -9.685 -147.725 -9.355 -147.395 ;
        RECT -9.685 -149.085 -9.355 -148.755 ;
        RECT -9.685 -150.445 -9.355 -150.115 ;
        RECT -9.685 -151.805 -9.355 -151.475 ;
        RECT -9.685 -153.165 -9.355 -152.835 ;
        RECT -9.685 -154.525 -9.355 -154.195 ;
        RECT -9.685 -155.885 -9.355 -155.555 ;
        RECT -9.685 -157.245 -9.355 -156.915 ;
        RECT -9.685 -158.605 -9.355 -158.275 ;
        RECT -9.685 -159.965 -9.355 -159.635 ;
        RECT -9.685 -161.325 -9.355 -160.995 ;
        RECT -9.685 -162.685 -9.355 -162.355 ;
        RECT -9.685 -164.045 -9.355 -163.715 ;
        RECT -9.685 -165.405 -9.355 -165.075 ;
        RECT -9.685 -166.765 -9.355 -166.435 ;
        RECT -9.685 -168.125 -9.355 -167.795 ;
        RECT -9.685 -169.485 -9.355 -169.155 ;
        RECT -9.685 -170.845 -9.355 -170.515 ;
        RECT -9.685 -172.205 -9.355 -171.875 ;
        RECT -9.685 -173.565 -9.355 -173.235 ;
        RECT -9.685 -174.925 -9.355 -174.595 ;
        RECT -9.685 -176.285 -9.355 -175.955 ;
        RECT -9.685 -177.645 -9.355 -177.315 ;
        RECT -9.685 -179.005 -9.355 -178.675 ;
        RECT -9.685 -181.725 -9.355 -181.395 ;
        RECT -9.685 -183.085 -9.355 -182.755 ;
        RECT -9.685 -184.445 -9.355 -184.115 ;
        RECT -9.685 -185.805 -9.355 -185.475 ;
        RECT -9.685 -187.165 -9.355 -186.835 ;
        RECT -9.685 -188.525 -9.355 -188.195 ;
        RECT -9.685 -189.885 -9.355 -189.555 ;
        RECT -9.685 -191.245 -9.355 -190.915 ;
        RECT -9.685 -192.605 -9.355 -192.275 ;
        RECT -9.685 -193.965 -9.355 -193.635 ;
        RECT -9.685 -195.325 -9.355 -194.995 ;
        RECT -9.685 -196.685 -9.355 -196.355 ;
        RECT -9.685 -198.045 -9.355 -197.715 ;
        RECT -9.685 -199.405 -9.355 -199.075 ;
        RECT -9.685 -200.765 -9.355 -200.435 ;
        RECT -9.685 -202.125 -9.355 -201.795 ;
        RECT -9.685 -203.485 -9.355 -203.155 ;
        RECT -9.68 -204.16 -9.36 133.765 ;
        RECT -9.685 132.52 -9.355 133.65 ;
        RECT -9.685 128.355 -9.355 128.685 ;
        RECT -9.685 126.995 -9.355 127.325 ;
        RECT -9.685 125.635 -9.355 125.965 ;
        RECT -9.685 124.275 -9.355 124.605 ;
        RECT -9.685 122.915 -9.355 123.245 ;
        RECT -9.685 121.555 -9.355 121.885 ;
        RECT -9.685 120.195 -9.355 120.525 ;
        RECT -9.685 118.835 -9.355 119.165 ;
        RECT -9.685 117.475 -9.355 117.805 ;
        RECT -9.685 110.675 -9.355 111.005 ;
        RECT -9.685 107.955 -9.355 108.285 ;
        RECT -9.685 103.875 -9.355 104.205 ;
        RECT -9.685 99.795 -9.355 100.125 ;
        RECT -9.685 97.075 -9.355 97.405 ;
        RECT -9.685 90.275 -9.355 90.605 ;
        RECT -9.685 88.915 -9.355 89.245 ;
        RECT -9.685 82.115 -9.355 82.445 ;
        RECT -9.685 79.395 -9.355 79.725 ;
        RECT -9.685 75.315 -9.355 75.645 ;
        RECT -9.685 71.235 -9.355 71.565 ;
        RECT -9.685 68.515 -9.355 68.845 ;
        RECT -9.685 61.715 -9.355 62.045 ;
        RECT -9.685 60.355 -9.355 60.685 ;
        RECT -9.685 50.835 -9.355 51.165 ;
        RECT -9.685 46.755 -9.355 47.085 ;
        RECT -9.685 42.675 -9.355 43.005 ;
        RECT -9.685 39.955 -9.355 40.285 ;
        RECT -9.685 33.155 -9.355 33.485 ;
        RECT -9.685 31.795 -9.355 32.125 ;
        RECT -9.685 29.075 -9.355 29.405 ;
        RECT -9.685 22.275 -9.355 22.605 ;
        RECT -9.685 19.555 -9.355 19.885 ;
        RECT -9.685 18.195 -9.355 18.525 ;
        RECT -9.685 11.395 -9.355 11.725 ;
        RECT -9.685 4.595 -9.355 4.925 ;
        RECT -9.685 3.235 -9.355 3.565 ;
        RECT -9.685 1.875 -9.355 2.205 ;
        RECT -9.685 0.515 -9.355 0.845 ;
        RECT -9.685 -0.845 -9.355 -0.515 ;
        RECT -9.685 -2.205 -9.355 -1.875 ;
        RECT -9.685 -3.565 -9.355 -3.235 ;
        RECT -9.685 -4.925 -9.355 -4.595 ;
        RECT -9.685 -7.645 -9.355 -7.315 ;
        RECT -9.685 -9.005 -9.355 -8.675 ;
        RECT -9.685 -13.085 -9.355 -12.755 ;
        RECT -9.685 -17.165 -9.355 -16.835 ;
        RECT -9.685 -21.245 -9.355 -20.915 ;
        RECT -9.685 -22.605 -9.355 -22.275 ;
        RECT -9.685 -23.965 -9.355 -23.635 ;
        RECT -9.685 -25.325 -9.355 -24.995 ;
        RECT -9.685 -26.685 -9.355 -26.355 ;
        RECT -9.685 -29.405 -9.355 -29.075 ;
        RECT -9.685 -30.765 -9.355 -30.435 ;
        RECT -9.685 -33.485 -9.355 -33.155 ;
        RECT -9.685 -36.205 -9.355 -35.875 ;
        RECT -9.685 -43.005 -9.355 -42.675 ;
        RECT -9.685 -44.365 -9.355 -44.035 ;
        RECT -9.685 -45.725 -9.355 -45.395 ;
        RECT -9.685 -47.085 -9.355 -46.755 ;
        RECT -9.685 -48.445 -9.355 -48.115 ;
        RECT -9.685 -49.805 -9.355 -49.475 ;
        RECT -9.685 -51.165 -9.355 -50.835 ;
        RECT -9.685 -53.885 -9.355 -53.555 ;
        RECT -9.685 -55.245 -9.355 -54.915 ;
        RECT -9.685 -56.605 -9.355 -56.275 ;
        RECT -9.685 -57.965 -9.355 -57.635 ;
        RECT -9.685 -59.325 -9.355 -58.995 ;
        RECT -9.685 -66.125 -9.355 -65.795 ;
        RECT -9.685 -68.845 -9.355 -68.515 ;
        RECT -9.685 -71.565 -9.355 -71.235 ;
        RECT -9.685 -72.925 -9.355 -72.595 ;
        RECT -9.685 -74.285 -9.355 -73.955 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.285 132.52 -22.955 133.65 ;
        RECT -23.285 128.355 -22.955 128.685 ;
        RECT -23.285 126.995 -22.955 127.325 ;
        RECT -23.285 125.635 -22.955 125.965 ;
        RECT -23.285 124.275 -22.955 124.605 ;
        RECT -23.285 122.915 -22.955 123.245 ;
        RECT -23.285 121.555 -22.955 121.885 ;
        RECT -23.285 120.195 -22.955 120.525 ;
        RECT -23.285 118.835 -22.955 119.165 ;
        RECT -23.285 117.475 -22.955 117.805 ;
        RECT -23.285 116.115 -22.955 116.445 ;
        RECT -23.285 114.755 -22.955 115.085 ;
        RECT -23.285 113.395 -22.955 113.725 ;
        RECT -23.285 112.035 -22.955 112.365 ;
        RECT -23.285 110.675 -22.955 111.005 ;
        RECT -23.285 109.315 -22.955 109.645 ;
        RECT -23.285 107.955 -22.955 108.285 ;
        RECT -23.285 106.595 -22.955 106.925 ;
        RECT -23.285 105.235 -22.955 105.565 ;
        RECT -23.285 103.875 -22.955 104.205 ;
        RECT -23.285 102.515 -22.955 102.845 ;
        RECT -23.285 101.155 -22.955 101.485 ;
        RECT -23.285 99.795 -22.955 100.125 ;
        RECT -23.285 98.435 -22.955 98.765 ;
        RECT -23.285 97.075 -22.955 97.405 ;
        RECT -23.285 95.715 -22.955 96.045 ;
        RECT -23.285 94.355 -22.955 94.685 ;
        RECT -23.285 92.995 -22.955 93.325 ;
        RECT -23.285 91.635 -22.955 91.965 ;
        RECT -23.285 90.275 -22.955 90.605 ;
        RECT -23.285 88.915 -22.955 89.245 ;
        RECT -23.285 87.555 -22.955 87.885 ;
        RECT -23.285 86.195 -22.955 86.525 ;
        RECT -23.285 84.835 -22.955 85.165 ;
        RECT -23.285 83.475 -22.955 83.805 ;
        RECT -23.285 82.115 -22.955 82.445 ;
        RECT -23.285 80.755 -22.955 81.085 ;
        RECT -23.285 79.395 -22.955 79.725 ;
        RECT -23.285 78.035 -22.955 78.365 ;
        RECT -23.285 76.675 -22.955 77.005 ;
        RECT -23.285 75.315 -22.955 75.645 ;
        RECT -23.285 73.955 -22.955 74.285 ;
        RECT -23.285 72.595 -22.955 72.925 ;
        RECT -23.285 71.235 -22.955 71.565 ;
        RECT -23.285 69.875 -22.955 70.205 ;
        RECT -23.285 68.515 -22.955 68.845 ;
        RECT -23.285 67.155 -22.955 67.485 ;
        RECT -23.285 65.795 -22.955 66.125 ;
        RECT -23.285 64.435 -22.955 64.765 ;
        RECT -23.285 63.075 -22.955 63.405 ;
        RECT -23.285 61.715 -22.955 62.045 ;
        RECT -23.285 60.355 -22.955 60.685 ;
        RECT -23.285 58.995 -22.955 59.325 ;
        RECT -23.285 57.635 -22.955 57.965 ;
        RECT -23.285 56.275 -22.955 56.605 ;
        RECT -23.285 54.915 -22.955 55.245 ;
        RECT -23.285 53.555 -22.955 53.885 ;
        RECT -23.285 52.195 -22.955 52.525 ;
        RECT -23.285 50.835 -22.955 51.165 ;
        RECT -23.285 49.475 -22.955 49.805 ;
        RECT -23.285 48.115 -22.955 48.445 ;
        RECT -23.285 46.755 -22.955 47.085 ;
        RECT -23.285 45.395 -22.955 45.725 ;
        RECT -23.285 44.035 -22.955 44.365 ;
        RECT -23.285 42.675 -22.955 43.005 ;
        RECT -23.285 41.315 -22.955 41.645 ;
        RECT -23.285 39.955 -22.955 40.285 ;
        RECT -23.285 38.595 -22.955 38.925 ;
        RECT -23.285 37.235 -22.955 37.565 ;
        RECT -23.285 35.875 -22.955 36.205 ;
        RECT -23.285 34.515 -22.955 34.845 ;
        RECT -23.285 33.155 -22.955 33.485 ;
        RECT -23.285 31.795 -22.955 32.125 ;
        RECT -23.285 30.435 -22.955 30.765 ;
        RECT -23.285 29.075 -22.955 29.405 ;
        RECT -23.285 27.715 -22.955 28.045 ;
        RECT -23.285 26.355 -22.955 26.685 ;
        RECT -23.285 24.995 -22.955 25.325 ;
        RECT -23.285 23.635 -22.955 23.965 ;
        RECT -23.285 22.275 -22.955 22.605 ;
        RECT -23.285 20.915 -22.955 21.245 ;
        RECT -23.285 19.555 -22.955 19.885 ;
        RECT -23.285 18.195 -22.955 18.525 ;
        RECT -23.285 16.835 -22.955 17.165 ;
        RECT -23.285 15.475 -22.955 15.805 ;
        RECT -23.285 14.115 -22.955 14.445 ;
        RECT -23.285 12.755 -22.955 13.085 ;
        RECT -23.285 11.395 -22.955 11.725 ;
        RECT -23.285 10.035 -22.955 10.365 ;
        RECT -23.285 8.675 -22.955 9.005 ;
        RECT -23.285 7.315 -22.955 7.645 ;
        RECT -23.285 5.955 -22.955 6.285 ;
        RECT -23.285 4.595 -22.955 4.925 ;
        RECT -23.285 3.235 -22.955 3.565 ;
        RECT -23.285 1.875 -22.955 2.205 ;
        RECT -23.285 0.515 -22.955 0.845 ;
        RECT -23.285 -0.845 -22.955 -0.515 ;
        RECT -23.285 -6.94 -22.955 -6.61 ;
        RECT -23.285 -7.645 -22.955 -7.315 ;
        RECT -23.285 -9.005 -22.955 -8.675 ;
        RECT -23.285 -13.085 -22.955 -12.755 ;
        RECT -23.285 -14.13 -22.955 -13.8 ;
        RECT -23.285 -17.165 -22.955 -16.835 ;
        RECT -23.285 -21.245 -22.955 -20.915 ;
        RECT -23.285 -26.685 -22.955 -26.355 ;
        RECT -23.285 -28.12 -22.955 -27.79 ;
        RECT -23.285 -29.405 -22.955 -29.075 ;
        RECT -23.285 -35.31 -22.955 -34.98 ;
        RECT -23.285 -43.005 -22.955 -42.675 ;
        RECT -23.285 -44.365 -22.955 -44.035 ;
        RECT -23.285 -45.725 -22.955 -45.395 ;
        RECT -23.285 -47.085 -22.955 -46.755 ;
        RECT -23.285 -48.445 -22.955 -48.115 ;
        RECT -23.285 -49.805 -22.955 -49.475 ;
        RECT -23.285 -51.165 -22.955 -50.835 ;
        RECT -23.285 -52.525 -22.955 -52.195 ;
        RECT -23.285 -53.885 -22.955 -53.555 ;
        RECT -23.285 -55.245 -22.955 -54.915 ;
        RECT -23.285 -56.605 -22.955 -56.275 ;
        RECT -23.285 -57.965 -22.955 -57.635 ;
        RECT -23.285 -59.325 -22.955 -58.995 ;
        RECT -23.285 -60.685 -22.955 -60.355 ;
        RECT -23.285 -62.045 -22.955 -61.715 ;
        RECT -23.285 -63.405 -22.955 -63.075 ;
        RECT -23.285 -64.765 -22.955 -64.435 ;
        RECT -23.285 -66.125 -22.955 -65.795 ;
        RECT -23.285 -67.485 -22.955 -67.155 ;
        RECT -23.285 -68.845 -22.955 -68.515 ;
        RECT -23.285 -70.205 -22.955 -69.875 ;
        RECT -23.285 -71.565 -22.955 -71.235 ;
        RECT -23.285 -72.925 -22.955 -72.595 ;
        RECT -23.285 -74.285 -22.955 -73.955 ;
        RECT -23.285 -75.645 -22.955 -75.315 ;
        RECT -23.285 -77.005 -22.955 -76.675 ;
        RECT -23.285 -78.365 -22.955 -78.035 ;
        RECT -23.285 -79.725 -22.955 -79.395 ;
        RECT -23.285 -81.085 -22.955 -80.755 ;
        RECT -23.285 -82.445 -22.955 -82.115 ;
        RECT -23.285 -83.805 -22.955 -83.475 ;
        RECT -23.285 -85.165 -22.955 -84.835 ;
        RECT -23.285 -86.525 -22.955 -86.195 ;
        RECT -23.285 -87.885 -22.955 -87.555 ;
        RECT -23.285 -89.245 -22.955 -88.915 ;
        RECT -23.285 -90.605 -22.955 -90.275 ;
        RECT -23.285 -91.965 -22.955 -91.635 ;
        RECT -23.285 -93.325 -22.955 -92.995 ;
        RECT -23.285 -94.685 -22.955 -94.355 ;
        RECT -23.285 -96.045 -22.955 -95.715 ;
        RECT -23.285 -97.405 -22.955 -97.075 ;
        RECT -23.285 -98.765 -22.955 -98.435 ;
        RECT -23.285 -100.125 -22.955 -99.795 ;
        RECT -23.285 -101.485 -22.955 -101.155 ;
        RECT -23.285 -102.845 -22.955 -102.515 ;
        RECT -23.285 -104.205 -22.955 -103.875 ;
        RECT -23.285 -109.645 -22.955 -109.315 ;
        RECT -23.285 -111.005 -22.955 -110.675 ;
        RECT -23.285 -112.365 -22.955 -112.035 ;
        RECT -23.285 -113.725 -22.955 -113.395 ;
        RECT -23.285 -115.085 -22.955 -114.755 ;
        RECT -23.285 -116.445 -22.955 -116.115 ;
        RECT -23.285 -117.805 -22.955 -117.475 ;
        RECT -23.285 -119.165 -22.955 -118.835 ;
        RECT -23.285 -120.525 -22.955 -120.195 ;
        RECT -23.285 -121.885 -22.955 -121.555 ;
        RECT -23.285 -123.245 -22.955 -122.915 ;
        RECT -23.285 -124.605 -22.955 -124.275 ;
        RECT -23.285 -125.965 -22.955 -125.635 ;
        RECT -23.285 -127.325 -22.955 -126.995 ;
        RECT -23.285 -128.685 -22.955 -128.355 ;
        RECT -23.285 -130.045 -22.955 -129.715 ;
        RECT -23.285 -131.405 -22.955 -131.075 ;
        RECT -23.285 -132.765 -22.955 -132.435 ;
        RECT -23.285 -134.125 -22.955 -133.795 ;
        RECT -23.285 -135.485 -22.955 -135.155 ;
        RECT -23.285 -136.845 -22.955 -136.515 ;
        RECT -23.285 -138.205 -22.955 -137.875 ;
        RECT -23.285 -139.565 -22.955 -139.235 ;
        RECT -23.285 -142.285 -22.955 -141.955 ;
        RECT -23.285 -143.645 -22.955 -143.315 ;
        RECT -23.285 -145.005 -22.955 -144.675 ;
        RECT -23.285 -146.365 -22.955 -146.035 ;
        RECT -23.285 -147.725 -22.955 -147.395 ;
        RECT -23.285 -149.085 -22.955 -148.755 ;
        RECT -23.285 -150.445 -22.955 -150.115 ;
        RECT -23.285 -151.805 -22.955 -151.475 ;
        RECT -23.285 -154.525 -22.955 -154.195 ;
        RECT -23.285 -155.885 -22.955 -155.555 ;
        RECT -23.285 -157.245 -22.955 -156.915 ;
        RECT -23.285 -158.605 -22.955 -158.275 ;
        RECT -23.285 -159.965 -22.955 -159.635 ;
        RECT -23.285 -161.325 -22.955 -160.995 ;
        RECT -23.285 -162.685 -22.955 -162.355 ;
        RECT -23.285 -165.405 -22.955 -165.075 ;
        RECT -23.285 -172.205 -22.955 -171.875 ;
        RECT -23.285 -173.565 -22.955 -173.235 ;
        RECT -23.285 -174.925 -22.955 -174.595 ;
        RECT -23.285 -176.285 -22.955 -175.955 ;
        RECT -23.285 -179.005 -22.955 -178.675 ;
        RECT -23.285 -180.365 -22.955 -180.035 ;
        RECT -23.285 -183.085 -22.955 -182.755 ;
        RECT -23.285 -184.445 -22.955 -184.115 ;
        RECT -23.285 -185.805 -22.955 -185.475 ;
        RECT -23.285 -189.885 -22.955 -189.555 ;
        RECT -23.285 -195.325 -22.955 -194.995 ;
        RECT -23.285 -196.685 -22.955 -196.355 ;
        RECT -23.285 -198.045 -22.955 -197.715 ;
        RECT -23.285 -199.405 -22.955 -199.075 ;
        RECT -23.285 -200.765 -22.955 -200.435 ;
        RECT -23.285 -202.125 -22.955 -201.795 ;
        RECT -23.285 -203.485 -22.955 -203.155 ;
        RECT -23.285 -204.845 -22.955 -204.515 ;
        RECT -23.285 -206.555 -22.955 -206.225 ;
        RECT -23.285 -207.565 -22.955 -207.235 ;
        RECT -23.28 -208.24 -22.96 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.285 -214.365 -22.955 -214.035 ;
        RECT -23.285 -215.725 -22.955 -215.395 ;
        RECT -23.285 -217.085 -22.955 -216.755 ;
        RECT -23.285 -218.445 -22.955 -218.115 ;
        RECT -23.285 -224.09 -22.955 -222.96 ;
        RECT -23.28 -224.205 -22.96 -210.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.925 132.52 -21.595 133.65 ;
        RECT -21.925 128.355 -21.595 128.685 ;
        RECT -21.925 126.995 -21.595 127.325 ;
        RECT -21.925 125.635 -21.595 125.965 ;
        RECT -21.925 124.275 -21.595 124.605 ;
        RECT -21.925 122.915 -21.595 123.245 ;
        RECT -21.925 121.555 -21.595 121.885 ;
        RECT -21.925 120.195 -21.595 120.525 ;
        RECT -21.925 118.835 -21.595 119.165 ;
        RECT -21.925 117.475 -21.595 117.805 ;
        RECT -21.925 116.115 -21.595 116.445 ;
        RECT -21.925 114.755 -21.595 115.085 ;
        RECT -21.925 113.395 -21.595 113.725 ;
        RECT -21.925 112.035 -21.595 112.365 ;
        RECT -21.925 110.675 -21.595 111.005 ;
        RECT -21.925 109.315 -21.595 109.645 ;
        RECT -21.925 107.955 -21.595 108.285 ;
        RECT -21.925 106.595 -21.595 106.925 ;
        RECT -21.925 105.235 -21.595 105.565 ;
        RECT -21.925 103.875 -21.595 104.205 ;
        RECT -21.925 102.515 -21.595 102.845 ;
        RECT -21.925 101.155 -21.595 101.485 ;
        RECT -21.925 99.795 -21.595 100.125 ;
        RECT -21.925 98.435 -21.595 98.765 ;
        RECT -21.925 97.075 -21.595 97.405 ;
        RECT -21.925 95.715 -21.595 96.045 ;
        RECT -21.925 94.355 -21.595 94.685 ;
        RECT -21.925 92.995 -21.595 93.325 ;
        RECT -21.925 91.635 -21.595 91.965 ;
        RECT -21.925 90.275 -21.595 90.605 ;
        RECT -21.925 88.915 -21.595 89.245 ;
        RECT -21.925 87.555 -21.595 87.885 ;
        RECT -21.925 86.195 -21.595 86.525 ;
        RECT -21.925 84.835 -21.595 85.165 ;
        RECT -21.925 83.475 -21.595 83.805 ;
        RECT -21.925 82.115 -21.595 82.445 ;
        RECT -21.925 80.755 -21.595 81.085 ;
        RECT -21.925 79.395 -21.595 79.725 ;
        RECT -21.925 78.035 -21.595 78.365 ;
        RECT -21.925 76.675 -21.595 77.005 ;
        RECT -21.925 75.315 -21.595 75.645 ;
        RECT -21.925 73.955 -21.595 74.285 ;
        RECT -21.925 72.595 -21.595 72.925 ;
        RECT -21.925 71.235 -21.595 71.565 ;
        RECT -21.925 69.875 -21.595 70.205 ;
        RECT -21.925 68.515 -21.595 68.845 ;
        RECT -21.925 67.155 -21.595 67.485 ;
        RECT -21.925 65.795 -21.595 66.125 ;
        RECT -21.925 64.435 -21.595 64.765 ;
        RECT -21.925 63.075 -21.595 63.405 ;
        RECT -21.925 61.715 -21.595 62.045 ;
        RECT -21.925 60.355 -21.595 60.685 ;
        RECT -21.925 58.995 -21.595 59.325 ;
        RECT -21.925 57.635 -21.595 57.965 ;
        RECT -21.925 56.275 -21.595 56.605 ;
        RECT -21.925 54.915 -21.595 55.245 ;
        RECT -21.925 53.555 -21.595 53.885 ;
        RECT -21.925 52.195 -21.595 52.525 ;
        RECT -21.925 50.835 -21.595 51.165 ;
        RECT -21.925 49.475 -21.595 49.805 ;
        RECT -21.925 48.115 -21.595 48.445 ;
        RECT -21.925 46.755 -21.595 47.085 ;
        RECT -21.925 45.395 -21.595 45.725 ;
        RECT -21.925 44.035 -21.595 44.365 ;
        RECT -21.925 42.675 -21.595 43.005 ;
        RECT -21.925 41.315 -21.595 41.645 ;
        RECT -21.925 39.955 -21.595 40.285 ;
        RECT -21.925 38.595 -21.595 38.925 ;
        RECT -21.925 37.235 -21.595 37.565 ;
        RECT -21.925 35.875 -21.595 36.205 ;
        RECT -21.925 34.515 -21.595 34.845 ;
        RECT -21.925 33.155 -21.595 33.485 ;
        RECT -21.925 31.795 -21.595 32.125 ;
        RECT -21.925 30.435 -21.595 30.765 ;
        RECT -21.925 29.075 -21.595 29.405 ;
        RECT -21.925 27.715 -21.595 28.045 ;
        RECT -21.925 26.355 -21.595 26.685 ;
        RECT -21.925 24.995 -21.595 25.325 ;
        RECT -21.925 23.635 -21.595 23.965 ;
        RECT -21.925 22.275 -21.595 22.605 ;
        RECT -21.925 20.915 -21.595 21.245 ;
        RECT -21.925 19.555 -21.595 19.885 ;
        RECT -21.925 18.195 -21.595 18.525 ;
        RECT -21.925 16.835 -21.595 17.165 ;
        RECT -21.925 15.475 -21.595 15.805 ;
        RECT -21.925 14.115 -21.595 14.445 ;
        RECT -21.925 12.755 -21.595 13.085 ;
        RECT -21.925 11.395 -21.595 11.725 ;
        RECT -21.925 10.035 -21.595 10.365 ;
        RECT -21.925 8.675 -21.595 9.005 ;
        RECT -21.925 7.315 -21.595 7.645 ;
        RECT -21.925 5.955 -21.595 6.285 ;
        RECT -21.925 4.595 -21.595 4.925 ;
        RECT -21.925 3.235 -21.595 3.565 ;
        RECT -21.925 1.875 -21.595 2.205 ;
        RECT -21.925 0.515 -21.595 0.845 ;
        RECT -21.925 -0.845 -21.595 -0.515 ;
        RECT -21.925 -2.205 -21.595 -1.875 ;
        RECT -21.925 -6.94 -21.595 -6.61 ;
        RECT -21.925 -7.645 -21.595 -7.315 ;
        RECT -21.925 -9.005 -21.595 -8.675 ;
        RECT -21.925 -13.085 -21.595 -12.755 ;
        RECT -21.925 -14.13 -21.595 -13.8 ;
        RECT -21.925 -17.165 -21.595 -16.835 ;
        RECT -21.92 -19.2 -21.6 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.925 -35.31 -21.595 -34.98 ;
        RECT -21.92 -40.96 -21.6 -31.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.925 -109.645 -21.595 -109.315 ;
        RECT -21.925 -111.005 -21.595 -110.675 ;
        RECT -21.925 -112.365 -21.595 -112.035 ;
        RECT -21.925 -113.725 -21.595 -113.395 ;
        RECT -21.925 -115.085 -21.595 -114.755 ;
        RECT -21.925 -116.445 -21.595 -116.115 ;
        RECT -21.925 -117.805 -21.595 -117.475 ;
        RECT -21.925 -119.165 -21.595 -118.835 ;
        RECT -21.925 -120.525 -21.595 -120.195 ;
        RECT -21.925 -121.885 -21.595 -121.555 ;
        RECT -21.925 -123.245 -21.595 -122.915 ;
        RECT -21.925 -124.605 -21.595 -124.275 ;
        RECT -21.925 -125.965 -21.595 -125.635 ;
        RECT -21.925 -127.325 -21.595 -126.995 ;
        RECT -21.925 -128.685 -21.595 -128.355 ;
        RECT -21.925 -130.045 -21.595 -129.715 ;
        RECT -21.925 -131.405 -21.595 -131.075 ;
        RECT -21.925 -132.765 -21.595 -132.435 ;
        RECT -21.925 -134.125 -21.595 -133.795 ;
        RECT -21.925 -135.485 -21.595 -135.155 ;
        RECT -21.925 -136.845 -21.595 -136.515 ;
        RECT -21.925 -138.205 -21.595 -137.875 ;
        RECT -21.925 -139.565 -21.595 -139.235 ;
        RECT -21.925 -142.285 -21.595 -141.955 ;
        RECT -21.925 -143.645 -21.595 -143.315 ;
        RECT -21.925 -145.005 -21.595 -144.675 ;
        RECT -21.925 -146.365 -21.595 -146.035 ;
        RECT -21.925 -147.725 -21.595 -147.395 ;
        RECT -21.925 -149.085 -21.595 -148.755 ;
        RECT -21.925 -150.445 -21.595 -150.115 ;
        RECT -21.925 -151.805 -21.595 -151.475 ;
        RECT -21.925 -154.525 -21.595 -154.195 ;
        RECT -21.925 -155.885 -21.595 -155.555 ;
        RECT -21.925 -157.245 -21.595 -156.915 ;
        RECT -21.925 -158.605 -21.595 -158.275 ;
        RECT -21.925 -159.965 -21.595 -159.635 ;
        RECT -21.925 -161.325 -21.595 -160.995 ;
        RECT -21.925 -162.685 -21.595 -162.355 ;
        RECT -21.925 -165.405 -21.595 -165.075 ;
        RECT -21.925 -172.205 -21.595 -171.875 ;
        RECT -21.925 -173.565 -21.595 -173.235 ;
        RECT -21.925 -174.925 -21.595 -174.595 ;
        RECT -21.925 -176.285 -21.595 -175.955 ;
        RECT -21.925 -179.005 -21.595 -178.675 ;
        RECT -21.925 -180.365 -21.595 -180.035 ;
        RECT -21.925 -183.085 -21.595 -182.755 ;
        RECT -21.925 -184.445 -21.595 -184.115 ;
        RECT -21.925 -185.805 -21.595 -185.475 ;
        RECT -21.925 -189.885 -21.595 -189.555 ;
        RECT -21.925 -195.325 -21.595 -194.995 ;
        RECT -21.925 -196.685 -21.595 -196.355 ;
        RECT -21.925 -198.045 -21.595 -197.715 ;
        RECT -21.925 -199.405 -21.595 -199.075 ;
        RECT -21.925 -200.765 -21.595 -200.435 ;
        RECT -21.925 -202.125 -21.595 -201.795 ;
        RECT -21.925 -203.485 -21.595 -203.155 ;
        RECT -21.925 -204.845 -21.595 -204.515 ;
        RECT -21.925 -206.555 -21.595 -206.225 ;
        RECT -21.925 -207.565 -21.595 -207.235 ;
        RECT -21.925 -214.365 -21.595 -214.035 ;
        RECT -21.925 -215.725 -21.595 -215.395 ;
        RECT -21.925 -217.085 -21.595 -216.755 ;
        RECT -21.925 -218.445 -21.595 -218.115 ;
        RECT -21.925 -224.09 -21.595 -222.96 ;
        RECT -21.92 -224.205 -21.6 -105.92 ;
    END
    PORT
      LAYER met3 ;
        RECT -20.565 132.52 -20.235 133.65 ;
        RECT -20.565 128.355 -20.235 128.685 ;
        RECT -20.565 126.995 -20.235 127.325 ;
        RECT -20.565 125.635 -20.235 125.965 ;
        RECT -20.565 124.275 -20.235 124.605 ;
        RECT -20.565 122.915 -20.235 123.245 ;
        RECT -20.565 121.555 -20.235 121.885 ;
        RECT -20.565 120.195 -20.235 120.525 ;
        RECT -20.565 118.835 -20.235 119.165 ;
        RECT -20.565 117.475 -20.235 117.805 ;
        RECT -20.565 116.115 -20.235 116.445 ;
        RECT -20.565 114.755 -20.235 115.085 ;
        RECT -20.565 113.395 -20.235 113.725 ;
        RECT -20.565 112.035 -20.235 112.365 ;
        RECT -20.565 110.675 -20.235 111.005 ;
        RECT -20.565 109.315 -20.235 109.645 ;
        RECT -20.565 107.955 -20.235 108.285 ;
        RECT -20.565 106.595 -20.235 106.925 ;
        RECT -20.565 105.235 -20.235 105.565 ;
        RECT -20.565 103.875 -20.235 104.205 ;
        RECT -20.565 102.515 -20.235 102.845 ;
        RECT -20.565 101.155 -20.235 101.485 ;
        RECT -20.565 99.795 -20.235 100.125 ;
        RECT -20.565 98.435 -20.235 98.765 ;
        RECT -20.565 97.075 -20.235 97.405 ;
        RECT -20.565 95.715 -20.235 96.045 ;
        RECT -20.565 94.355 -20.235 94.685 ;
        RECT -20.565 92.995 -20.235 93.325 ;
        RECT -20.565 91.635 -20.235 91.965 ;
        RECT -20.565 90.275 -20.235 90.605 ;
        RECT -20.565 88.915 -20.235 89.245 ;
        RECT -20.565 87.555 -20.235 87.885 ;
        RECT -20.565 86.195 -20.235 86.525 ;
        RECT -20.565 84.835 -20.235 85.165 ;
        RECT -20.565 83.475 -20.235 83.805 ;
        RECT -20.565 82.115 -20.235 82.445 ;
        RECT -20.565 80.755 -20.235 81.085 ;
        RECT -20.565 79.395 -20.235 79.725 ;
        RECT -20.565 78.035 -20.235 78.365 ;
        RECT -20.565 76.675 -20.235 77.005 ;
        RECT -20.565 75.315 -20.235 75.645 ;
        RECT -20.565 73.955 -20.235 74.285 ;
        RECT -20.565 72.595 -20.235 72.925 ;
        RECT -20.565 71.235 -20.235 71.565 ;
        RECT -20.565 69.875 -20.235 70.205 ;
        RECT -20.565 68.515 -20.235 68.845 ;
        RECT -20.565 67.155 -20.235 67.485 ;
        RECT -20.565 65.795 -20.235 66.125 ;
        RECT -20.565 64.435 -20.235 64.765 ;
        RECT -20.565 63.075 -20.235 63.405 ;
        RECT -20.565 61.715 -20.235 62.045 ;
        RECT -20.565 60.355 -20.235 60.685 ;
        RECT -20.565 58.995 -20.235 59.325 ;
        RECT -20.565 57.635 -20.235 57.965 ;
        RECT -20.565 56.275 -20.235 56.605 ;
        RECT -20.565 54.915 -20.235 55.245 ;
        RECT -20.565 53.555 -20.235 53.885 ;
        RECT -20.565 52.195 -20.235 52.525 ;
        RECT -20.565 50.835 -20.235 51.165 ;
        RECT -20.565 49.475 -20.235 49.805 ;
        RECT -20.565 48.115 -20.235 48.445 ;
        RECT -20.565 46.755 -20.235 47.085 ;
        RECT -20.565 45.395 -20.235 45.725 ;
        RECT -20.565 44.035 -20.235 44.365 ;
        RECT -20.565 42.675 -20.235 43.005 ;
        RECT -20.565 41.315 -20.235 41.645 ;
        RECT -20.565 39.955 -20.235 40.285 ;
        RECT -20.565 38.595 -20.235 38.925 ;
        RECT -20.565 37.235 -20.235 37.565 ;
        RECT -20.565 35.875 -20.235 36.205 ;
        RECT -20.565 34.515 -20.235 34.845 ;
        RECT -20.565 33.155 -20.235 33.485 ;
        RECT -20.565 31.795 -20.235 32.125 ;
        RECT -20.565 30.435 -20.235 30.765 ;
        RECT -20.565 29.075 -20.235 29.405 ;
        RECT -20.565 27.715 -20.235 28.045 ;
        RECT -20.565 26.355 -20.235 26.685 ;
        RECT -20.565 24.995 -20.235 25.325 ;
        RECT -20.565 23.635 -20.235 23.965 ;
        RECT -20.565 22.275 -20.235 22.605 ;
        RECT -20.565 20.915 -20.235 21.245 ;
        RECT -20.565 19.555 -20.235 19.885 ;
        RECT -20.565 18.195 -20.235 18.525 ;
        RECT -20.565 16.835 -20.235 17.165 ;
        RECT -20.565 15.475 -20.235 15.805 ;
        RECT -20.565 14.115 -20.235 14.445 ;
        RECT -20.565 12.755 -20.235 13.085 ;
        RECT -20.565 11.395 -20.235 11.725 ;
        RECT -20.565 10.035 -20.235 10.365 ;
        RECT -20.565 8.675 -20.235 9.005 ;
        RECT -20.565 7.315 -20.235 7.645 ;
        RECT -20.565 5.955 -20.235 6.285 ;
        RECT -20.565 4.595 -20.235 4.925 ;
        RECT -20.565 3.235 -20.235 3.565 ;
        RECT -20.565 1.875 -20.235 2.205 ;
        RECT -20.565 0.515 -20.235 0.845 ;
        RECT -20.565 -0.845 -20.235 -0.515 ;
        RECT -20.565 -2.205 -20.235 -1.875 ;
        RECT -20.565 -6.94 -20.235 -6.61 ;
        RECT -20.565 -7.645 -20.235 -7.315 ;
        RECT -20.565 -9.005 -20.235 -8.675 ;
        RECT -20.565 -13.085 -20.235 -12.755 ;
        RECT -20.565 -14.13 -20.235 -13.8 ;
        RECT -20.565 -17.165 -20.235 -16.835 ;
        RECT -20.56 -18.52 -20.24 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -20.565 -35.31 -20.235 -34.98 ;
        RECT -20.56 -39.6 -20.24 -33.84 ;
    END
    PORT
      LAYER met3 ;
        RECT -20.565 -109.645 -20.235 -109.315 ;
        RECT -20.565 -111.005 -20.235 -110.675 ;
        RECT -20.565 -112.365 -20.235 -112.035 ;
        RECT -20.565 -113.725 -20.235 -113.395 ;
        RECT -20.565 -116.445 -20.235 -116.115 ;
        RECT -20.565 -117.805 -20.235 -117.475 ;
        RECT -20.565 -119.165 -20.235 -118.835 ;
        RECT -20.565 -120.525 -20.235 -120.195 ;
        RECT -20.565 -121.885 -20.235 -121.555 ;
        RECT -20.565 -123.245 -20.235 -122.915 ;
        RECT -20.565 -125.965 -20.235 -125.635 ;
        RECT -20.565 -127.325 -20.235 -126.995 ;
        RECT -20.565 -128.685 -20.235 -128.355 ;
        RECT -20.565 -132.765 -20.235 -132.435 ;
        RECT -20.565 -134.125 -20.235 -133.795 ;
        RECT -20.565 -135.485 -20.235 -135.155 ;
        RECT -20.565 -136.845 -20.235 -136.515 ;
        RECT -20.565 -138.205 -20.235 -137.875 ;
        RECT -20.565 -139.565 -20.235 -139.235 ;
        RECT -20.565 -143.645 -20.235 -143.315 ;
        RECT -20.565 -145.005 -20.235 -144.675 ;
        RECT -20.565 -147.725 -20.235 -147.395 ;
        RECT -20.565 -149.085 -20.235 -148.755 ;
        RECT -20.565 -150.445 -20.235 -150.115 ;
        RECT -20.565 -151.805 -20.235 -151.475 ;
        RECT -20.565 -154.525 -20.235 -154.195 ;
        RECT -20.565 -155.885 -20.235 -155.555 ;
        RECT -20.565 -157.245 -20.235 -156.915 ;
        RECT -20.565 -158.605 -20.235 -158.275 ;
        RECT -20.565 -159.965 -20.235 -159.635 ;
        RECT -20.565 -161.325 -20.235 -160.995 ;
        RECT -20.565 -162.685 -20.235 -162.355 ;
        RECT -20.565 -165.405 -20.235 -165.075 ;
        RECT -20.565 -174.925 -20.235 -174.595 ;
        RECT -20.565 -176.285 -20.235 -175.955 ;
        RECT -20.565 -179.005 -20.235 -178.675 ;
        RECT -20.565 -184.445 -20.235 -184.115 ;
        RECT -20.565 -189.885 -20.235 -189.555 ;
        RECT -20.565 -193.965 -20.235 -193.635 ;
        RECT -20.565 -195.325 -20.235 -194.995 ;
        RECT -20.565 -196.685 -20.235 -196.355 ;
        RECT -20.565 -198.045 -20.235 -197.715 ;
        RECT -20.565 -199.405 -20.235 -199.075 ;
        RECT -20.565 -200.765 -20.235 -200.435 ;
        RECT -20.565 -202.125 -20.235 -201.795 ;
        RECT -20.565 -203.485 -20.235 -203.155 ;
        RECT -20.565 -204.845 -20.235 -204.515 ;
        RECT -20.565 -206.555 -20.235 -206.225 ;
        RECT -20.565 -207.565 -20.235 -207.235 ;
        RECT -20.565 -214.365 -20.235 -214.035 ;
        RECT -20.565 -215.725 -20.235 -215.395 ;
        RECT -20.565 -217.085 -20.235 -216.755 ;
        RECT -20.565 -218.445 -20.235 -218.115 ;
        RECT -20.565 -224.09 -20.235 -222.96 ;
        RECT -20.56 -224.205 -20.24 -105.24 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.205 132.52 -18.875 133.65 ;
        RECT -19.205 128.355 -18.875 128.685 ;
        RECT -19.205 126.995 -18.875 127.325 ;
        RECT -19.205 125.635 -18.875 125.965 ;
        RECT -19.205 124.275 -18.875 124.605 ;
        RECT -19.205 122.915 -18.875 123.245 ;
        RECT -19.205 121.555 -18.875 121.885 ;
        RECT -19.205 120.195 -18.875 120.525 ;
        RECT -19.205 118.835 -18.875 119.165 ;
        RECT -19.205 117.475 -18.875 117.805 ;
        RECT -19.205 116.115 -18.875 116.445 ;
        RECT -19.205 114.755 -18.875 115.085 ;
        RECT -19.205 113.395 -18.875 113.725 ;
        RECT -19.205 112.035 -18.875 112.365 ;
        RECT -19.205 110.675 -18.875 111.005 ;
        RECT -19.205 109.315 -18.875 109.645 ;
        RECT -19.205 107.955 -18.875 108.285 ;
        RECT -19.205 106.595 -18.875 106.925 ;
        RECT -19.205 105.235 -18.875 105.565 ;
        RECT -19.205 103.875 -18.875 104.205 ;
        RECT -19.205 102.515 -18.875 102.845 ;
        RECT -19.205 101.155 -18.875 101.485 ;
        RECT -19.205 99.795 -18.875 100.125 ;
        RECT -19.205 98.435 -18.875 98.765 ;
        RECT -19.205 97.075 -18.875 97.405 ;
        RECT -19.205 95.715 -18.875 96.045 ;
        RECT -19.205 94.355 -18.875 94.685 ;
        RECT -19.205 92.995 -18.875 93.325 ;
        RECT -19.205 91.635 -18.875 91.965 ;
        RECT -19.205 90.275 -18.875 90.605 ;
        RECT -19.205 88.915 -18.875 89.245 ;
        RECT -19.205 87.555 -18.875 87.885 ;
        RECT -19.205 86.195 -18.875 86.525 ;
        RECT -19.205 84.835 -18.875 85.165 ;
        RECT -19.205 83.475 -18.875 83.805 ;
        RECT -19.205 82.115 -18.875 82.445 ;
        RECT -19.205 80.755 -18.875 81.085 ;
        RECT -19.205 79.395 -18.875 79.725 ;
        RECT -19.205 78.035 -18.875 78.365 ;
        RECT -19.205 76.675 -18.875 77.005 ;
        RECT -19.205 75.315 -18.875 75.645 ;
        RECT -19.205 73.955 -18.875 74.285 ;
        RECT -19.205 72.595 -18.875 72.925 ;
        RECT -19.205 71.235 -18.875 71.565 ;
        RECT -19.205 69.875 -18.875 70.205 ;
        RECT -19.205 68.515 -18.875 68.845 ;
        RECT -19.205 67.155 -18.875 67.485 ;
        RECT -19.205 65.795 -18.875 66.125 ;
        RECT -19.205 64.435 -18.875 64.765 ;
        RECT -19.205 63.075 -18.875 63.405 ;
        RECT -19.205 61.715 -18.875 62.045 ;
        RECT -19.205 60.355 -18.875 60.685 ;
        RECT -19.205 58.995 -18.875 59.325 ;
        RECT -19.205 57.635 -18.875 57.965 ;
        RECT -19.205 56.275 -18.875 56.605 ;
        RECT -19.205 54.915 -18.875 55.245 ;
        RECT -19.205 53.555 -18.875 53.885 ;
        RECT -19.205 52.195 -18.875 52.525 ;
        RECT -19.205 50.835 -18.875 51.165 ;
        RECT -19.205 49.475 -18.875 49.805 ;
        RECT -19.205 48.115 -18.875 48.445 ;
        RECT -19.205 46.755 -18.875 47.085 ;
        RECT -19.205 45.395 -18.875 45.725 ;
        RECT -19.205 44.035 -18.875 44.365 ;
        RECT -19.205 42.675 -18.875 43.005 ;
        RECT -19.205 41.315 -18.875 41.645 ;
        RECT -19.205 39.955 -18.875 40.285 ;
        RECT -19.205 38.595 -18.875 38.925 ;
        RECT -19.205 37.235 -18.875 37.565 ;
        RECT -19.205 35.875 -18.875 36.205 ;
        RECT -19.205 34.515 -18.875 34.845 ;
        RECT -19.205 33.155 -18.875 33.485 ;
        RECT -19.205 31.795 -18.875 32.125 ;
        RECT -19.205 30.435 -18.875 30.765 ;
        RECT -19.205 29.075 -18.875 29.405 ;
        RECT -19.205 27.715 -18.875 28.045 ;
        RECT -19.205 26.355 -18.875 26.685 ;
        RECT -19.205 24.995 -18.875 25.325 ;
        RECT -19.205 23.635 -18.875 23.965 ;
        RECT -19.205 22.275 -18.875 22.605 ;
        RECT -19.205 20.915 -18.875 21.245 ;
        RECT -19.205 19.555 -18.875 19.885 ;
        RECT -19.205 18.195 -18.875 18.525 ;
        RECT -19.205 16.835 -18.875 17.165 ;
        RECT -19.205 15.475 -18.875 15.805 ;
        RECT -19.205 14.115 -18.875 14.445 ;
        RECT -19.205 12.755 -18.875 13.085 ;
        RECT -19.205 11.395 -18.875 11.725 ;
        RECT -19.205 10.035 -18.875 10.365 ;
        RECT -19.205 8.675 -18.875 9.005 ;
        RECT -19.205 7.315 -18.875 7.645 ;
        RECT -19.205 5.955 -18.875 6.285 ;
        RECT -19.205 4.595 -18.875 4.925 ;
        RECT -19.205 3.235 -18.875 3.565 ;
        RECT -19.205 1.875 -18.875 2.205 ;
        RECT -19.205 0.515 -18.875 0.845 ;
        RECT -19.205 -0.845 -18.875 -0.515 ;
        RECT -19.205 -2.205 -18.875 -1.875 ;
        RECT -19.205 -6.94 -18.875 -6.61 ;
        RECT -19.205 -7.645 -18.875 -7.315 ;
        RECT -19.205 -9.005 -18.875 -8.675 ;
        RECT -19.205 -13.085 -18.875 -12.755 ;
        RECT -19.205 -14.13 -18.875 -13.8 ;
        RECT -19.205 -17.165 -18.875 -16.835 ;
        RECT -19.2 -17.84 -18.88 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.205 -109.645 -18.875 -109.315 ;
        RECT -19.205 -111.005 -18.875 -110.675 ;
        RECT -19.205 -112.365 -18.875 -112.035 ;
        RECT -19.205 -113.725 -18.875 -113.395 ;
        RECT -19.205 -114.87 -18.875 -114.54 ;
        RECT -19.205 -116.445 -18.875 -116.115 ;
        RECT -19.205 -117.805 -18.875 -117.475 ;
        RECT -19.205 -119.165 -18.875 -118.835 ;
        RECT -19.205 -120.525 -18.875 -120.195 ;
        RECT -19.205 -121.885 -18.875 -121.555 ;
        RECT -19.205 -123.245 -18.875 -122.915 ;
        RECT -19.205 -125.965 -18.875 -125.635 ;
        RECT -19.205 -127.325 -18.875 -126.995 ;
        RECT -19.205 -128.685 -18.875 -128.355 ;
        RECT -19.205 -132.765 -18.875 -132.435 ;
        RECT -19.205 -134.125 -18.875 -133.795 ;
        RECT -19.205 -135.485 -18.875 -135.155 ;
        RECT -19.205 -136.845 -18.875 -136.515 ;
        RECT -19.205 -138.205 -18.875 -137.875 ;
        RECT -19.205 -139.565 -18.875 -139.235 ;
        RECT -19.205 -145.005 -18.875 -144.675 ;
        RECT -19.205 -147.725 -18.875 -147.395 ;
        RECT -19.205 -149.085 -18.875 -148.755 ;
        RECT -19.205 -150.445 -18.875 -150.115 ;
        RECT -19.205 -151.805 -18.875 -151.475 ;
        RECT -19.205 -154.525 -18.875 -154.195 ;
        RECT -19.205 -155.885 -18.875 -155.555 ;
        RECT -19.205 -157.245 -18.875 -156.915 ;
        RECT -19.205 -158.605 -18.875 -158.275 ;
        RECT -19.205 -159.965 -18.875 -159.635 ;
        RECT -19.205 -161.325 -18.875 -160.995 ;
        RECT -19.205 -162.685 -18.875 -162.355 ;
        RECT -19.205 -165.405 -18.875 -165.075 ;
        RECT -19.205 -174.925 -18.875 -174.595 ;
        RECT -19.205 -176.285 -18.875 -175.955 ;
        RECT -19.205 -181.725 -18.875 -181.395 ;
        RECT -19.205 -189.885 -18.875 -189.555 ;
        RECT -19.205 -195.325 -18.875 -194.995 ;
        RECT -19.205 -196.685 -18.875 -196.355 ;
        RECT -19.205 -198.045 -18.875 -197.715 ;
        RECT -19.205 -199.405 -18.875 -199.075 ;
        RECT -19.205 -200.765 -18.875 -200.435 ;
        RECT -19.205 -202.125 -18.875 -201.795 ;
        RECT -19.205 -203.485 -18.875 -203.155 ;
        RECT -19.205 -206.555 -18.875 -206.225 ;
        RECT -19.205 -207.565 -18.875 -207.235 ;
        RECT -19.2 -208.92 -18.88 -107.96 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.205 -214.365 -18.875 -214.035 ;
        RECT -19.205 -215.725 -18.875 -215.395 ;
        RECT -19.205 -217.085 -18.875 -216.755 ;
        RECT -19.205 -218.445 -18.875 -218.115 ;
        RECT -19.205 -224.09 -18.875 -222.96 ;
        RECT -19.2 -224.205 -18.88 -212 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.845 65.795 -17.515 66.125 ;
        RECT -17.845 64.435 -17.515 64.765 ;
        RECT -17.845 63.075 -17.515 63.405 ;
        RECT -17.845 61.715 -17.515 62.045 ;
        RECT -17.845 60.355 -17.515 60.685 ;
        RECT -17.845 58.995 -17.515 59.325 ;
        RECT -17.845 57.635 -17.515 57.965 ;
        RECT -17.845 56.275 -17.515 56.605 ;
        RECT -17.845 54.915 -17.515 55.245 ;
        RECT -17.845 53.555 -17.515 53.885 ;
        RECT -17.845 52.195 -17.515 52.525 ;
        RECT -17.845 50.835 -17.515 51.165 ;
        RECT -17.845 49.475 -17.515 49.805 ;
        RECT -17.845 48.115 -17.515 48.445 ;
        RECT -17.845 46.755 -17.515 47.085 ;
        RECT -17.845 45.395 -17.515 45.725 ;
        RECT -17.845 44.035 -17.515 44.365 ;
        RECT -17.845 42.675 -17.515 43.005 ;
        RECT -17.845 41.315 -17.515 41.645 ;
        RECT -17.845 39.955 -17.515 40.285 ;
        RECT -17.845 38.595 -17.515 38.925 ;
        RECT -17.845 37.235 -17.515 37.565 ;
        RECT -17.845 35.875 -17.515 36.205 ;
        RECT -17.845 34.515 -17.515 34.845 ;
        RECT -17.845 33.155 -17.515 33.485 ;
        RECT -17.845 31.795 -17.515 32.125 ;
        RECT -17.845 30.435 -17.515 30.765 ;
        RECT -17.845 29.075 -17.515 29.405 ;
        RECT -17.845 27.715 -17.515 28.045 ;
        RECT -17.845 26.355 -17.515 26.685 ;
        RECT -17.845 24.995 -17.515 25.325 ;
        RECT -17.845 23.635 -17.515 23.965 ;
        RECT -17.845 22.275 -17.515 22.605 ;
        RECT -17.845 20.915 -17.515 21.245 ;
        RECT -17.845 19.555 -17.515 19.885 ;
        RECT -17.845 18.195 -17.515 18.525 ;
        RECT -17.845 16.835 -17.515 17.165 ;
        RECT -17.845 15.475 -17.515 15.805 ;
        RECT -17.845 14.115 -17.515 14.445 ;
        RECT -17.845 12.755 -17.515 13.085 ;
        RECT -17.845 11.395 -17.515 11.725 ;
        RECT -17.845 10.035 -17.515 10.365 ;
        RECT -17.845 8.675 -17.515 9.005 ;
        RECT -17.845 7.315 -17.515 7.645 ;
        RECT -17.845 5.955 -17.515 6.285 ;
        RECT -17.845 4.595 -17.515 4.925 ;
        RECT -17.845 3.235 -17.515 3.565 ;
        RECT -17.845 1.875 -17.515 2.205 ;
        RECT -17.845 0.515 -17.515 0.845 ;
        RECT -17.845 -0.845 -17.515 -0.515 ;
        RECT -17.845 -2.205 -17.515 -1.875 ;
        RECT -17.845 -6.94 -17.515 -6.61 ;
        RECT -17.845 -7.645 -17.515 -7.315 ;
        RECT -17.845 -9.005 -17.515 -8.675 ;
        RECT -17.845 -13.085 -17.515 -12.755 ;
        RECT -17.845 -14.13 -17.515 -13.8 ;
        RECT -17.845 -17.165 -17.515 -16.835 ;
        RECT -17.845 -21.245 -17.515 -20.915 ;
        RECT -17.845 -22.605 -17.515 -22.275 ;
        RECT -17.845 -26.685 -17.515 -26.355 ;
        RECT -17.845 -28.12 -17.515 -27.79 ;
        RECT -17.845 -29.405 -17.515 -29.075 ;
        RECT -17.845 -30.765 -17.515 -30.435 ;
        RECT -17.845 -33.485 -17.515 -33.155 ;
        RECT -17.845 -35.31 -17.515 -34.98 ;
        RECT -17.845 -36.205 -17.515 -35.875 ;
        RECT -17.845 -43.005 -17.515 -42.675 ;
        RECT -17.845 -44.365 -17.515 -44.035 ;
        RECT -17.845 -45.725 -17.515 -45.395 ;
        RECT -17.845 -47.085 -17.515 -46.755 ;
        RECT -17.845 -48.445 -17.515 -48.115 ;
        RECT -17.845 -49.805 -17.515 -49.475 ;
        RECT -17.845 -51.165 -17.515 -50.835 ;
        RECT -17.845 -52.15 -17.515 -51.82 ;
        RECT -17.845 -53.885 -17.515 -53.555 ;
        RECT -17.845 -55.245 -17.515 -54.915 ;
        RECT -17.845 -56.605 -17.515 -56.275 ;
        RECT -17.845 -57.965 -17.515 -57.635 ;
        RECT -17.845 -59.325 -17.515 -58.995 ;
        RECT -17.845 -60.685 -17.515 -60.355 ;
        RECT -17.845 -64.765 -17.515 -64.435 ;
        RECT -17.845 -66.125 -17.515 -65.795 ;
        RECT -17.845 -67.485 -17.515 -67.155 ;
        RECT -17.845 -68.845 -17.515 -68.515 ;
        RECT -17.845 -70.69 -17.515 -70.36 ;
        RECT -17.845 -71.565 -17.515 -71.235 ;
        RECT -17.845 -72.925 -17.515 -72.595 ;
        RECT -17.845 -74.285 -17.515 -73.955 ;
        RECT -17.845 -75.645 -17.515 -75.315 ;
        RECT -17.845 -77.005 -17.515 -76.675 ;
        RECT -17.845 -78.365 -17.515 -78.035 ;
        RECT -17.845 -81.085 -17.515 -80.755 ;
        RECT -17.845 -82.445 -17.515 -82.115 ;
        RECT -17.845 -83.805 -17.515 -83.475 ;
        RECT -17.845 -85.165 -17.515 -84.835 ;
        RECT -17.845 -87.885 -17.515 -87.555 ;
        RECT -17.845 -89.245 -17.515 -88.915 ;
        RECT -17.845 -90.605 -17.515 -90.275 ;
        RECT -17.845 -91.965 -17.515 -91.635 ;
        RECT -17.845 -93.325 -17.515 -92.995 ;
        RECT -17.845 -94.685 -17.515 -94.355 ;
        RECT -17.845 -96.33 -17.515 -96 ;
        RECT -17.845 -97.405 -17.515 -97.075 ;
        RECT -17.845 -98.765 -17.515 -98.435 ;
        RECT -17.845 -100.125 -17.515 -99.795 ;
        RECT -17.845 -101.485 -17.515 -101.155 ;
        RECT -17.845 -102.845 -17.515 -102.515 ;
        RECT -17.845 -104.205 -17.515 -103.875 ;
        RECT -17.845 -106.925 -17.515 -106.595 ;
        RECT -17.845 -108.285 -17.515 -107.955 ;
        RECT -17.845 -109.645 -17.515 -109.315 ;
        RECT -17.845 -111.005 -17.515 -110.675 ;
        RECT -17.845 -113.725 -17.515 -113.395 ;
        RECT -17.845 -114.87 -17.515 -114.54 ;
        RECT -17.845 -116.445 -17.515 -116.115 ;
        RECT -17.845 -117.805 -17.515 -117.475 ;
        RECT -17.845 -119.165 -17.515 -118.835 ;
        RECT -17.845 -120.525 -17.515 -120.195 ;
        RECT -17.845 -121.885 -17.515 -121.555 ;
        RECT -17.845 -123.245 -17.515 -122.915 ;
        RECT -17.845 -125.965 -17.515 -125.635 ;
        RECT -17.845 -127.325 -17.515 -126.995 ;
        RECT -17.845 -128.685 -17.515 -128.355 ;
        RECT -17.845 -132.765 -17.515 -132.435 ;
        RECT -17.845 -134.125 -17.515 -133.795 ;
        RECT -17.845 -135.485 -17.515 -135.155 ;
        RECT -17.845 -136.845 -17.515 -136.515 ;
        RECT -17.845 -138.205 -17.515 -137.875 ;
        RECT -17.845 -145.005 -17.515 -144.675 ;
        RECT -17.845 -147.725 -17.515 -147.395 ;
        RECT -17.845 -149.085 -17.515 -148.755 ;
        RECT -17.845 -150.445 -17.515 -150.115 ;
        RECT -17.845 -151.805 -17.515 -151.475 ;
        RECT -17.845 -155.885 -17.515 -155.555 ;
        RECT -17.845 -157.245 -17.515 -156.915 ;
        RECT -17.845 -158.605 -17.515 -158.275 ;
        RECT -17.845 -159.965 -17.515 -159.635 ;
        RECT -17.845 -161.325 -17.515 -160.995 ;
        RECT -17.845 -162.685 -17.515 -162.355 ;
        RECT -17.845 -165.405 -17.515 -165.075 ;
        RECT -17.845 -174.925 -17.515 -174.595 ;
        RECT -17.845 -176.285 -17.515 -175.955 ;
        RECT -17.845 -181.725 -17.515 -181.395 ;
        RECT -17.845 -183.085 -17.515 -182.755 ;
        RECT -17.845 -189.885 -17.515 -189.555 ;
        RECT -17.845 -195.325 -17.515 -194.995 ;
        RECT -17.845 -196.685 -17.515 -196.355 ;
        RECT -17.845 -198.045 -17.515 -197.715 ;
        RECT -17.845 -199.405 -17.515 -199.075 ;
        RECT -17.845 -200.765 -17.515 -200.435 ;
        RECT -17.845 -202.125 -17.515 -201.795 ;
        RECT -17.845 -203.485 -17.515 -203.155 ;
        RECT -17.845 -206.555 -17.515 -206.225 ;
        RECT -17.845 -207.565 -17.515 -207.235 ;
        RECT -17.845 -210.285 -17.515 -209.955 ;
        RECT -17.845 -214.365 -17.515 -214.035 ;
        RECT -17.845 -215.725 -17.515 -215.395 ;
        RECT -17.845 -217.085 -17.515 -216.755 ;
        RECT -17.845 -218.445 -17.515 -218.115 ;
        RECT -17.845 -224.09 -17.515 -222.96 ;
        RECT -17.84 -224.205 -17.52 133.765 ;
        RECT -17.845 132.52 -17.515 133.65 ;
        RECT -17.845 128.355 -17.515 128.685 ;
        RECT -17.845 126.995 -17.515 127.325 ;
        RECT -17.845 125.635 -17.515 125.965 ;
        RECT -17.845 124.275 -17.515 124.605 ;
        RECT -17.845 122.915 -17.515 123.245 ;
        RECT -17.845 121.555 -17.515 121.885 ;
        RECT -17.845 120.195 -17.515 120.525 ;
        RECT -17.845 118.835 -17.515 119.165 ;
        RECT -17.845 117.475 -17.515 117.805 ;
        RECT -17.845 116.115 -17.515 116.445 ;
        RECT -17.845 114.755 -17.515 115.085 ;
        RECT -17.845 113.395 -17.515 113.725 ;
        RECT -17.845 112.035 -17.515 112.365 ;
        RECT -17.845 110.675 -17.515 111.005 ;
        RECT -17.845 109.315 -17.515 109.645 ;
        RECT -17.845 107.955 -17.515 108.285 ;
        RECT -17.845 106.595 -17.515 106.925 ;
        RECT -17.845 105.235 -17.515 105.565 ;
        RECT -17.845 103.875 -17.515 104.205 ;
        RECT -17.845 102.515 -17.515 102.845 ;
        RECT -17.845 101.155 -17.515 101.485 ;
        RECT -17.845 99.795 -17.515 100.125 ;
        RECT -17.845 98.435 -17.515 98.765 ;
        RECT -17.845 97.075 -17.515 97.405 ;
        RECT -17.845 95.715 -17.515 96.045 ;
        RECT -17.845 94.355 -17.515 94.685 ;
        RECT -17.845 92.995 -17.515 93.325 ;
        RECT -17.845 91.635 -17.515 91.965 ;
        RECT -17.845 90.275 -17.515 90.605 ;
        RECT -17.845 88.915 -17.515 89.245 ;
        RECT -17.845 87.555 -17.515 87.885 ;
        RECT -17.845 86.195 -17.515 86.525 ;
        RECT -17.845 84.835 -17.515 85.165 ;
        RECT -17.845 83.475 -17.515 83.805 ;
        RECT -17.845 82.115 -17.515 82.445 ;
        RECT -17.845 80.755 -17.515 81.085 ;
        RECT -17.845 79.395 -17.515 79.725 ;
        RECT -17.845 78.035 -17.515 78.365 ;
        RECT -17.845 76.675 -17.515 77.005 ;
        RECT -17.845 75.315 -17.515 75.645 ;
        RECT -17.845 73.955 -17.515 74.285 ;
        RECT -17.845 72.595 -17.515 72.925 ;
        RECT -17.845 71.235 -17.515 71.565 ;
        RECT -17.845 69.875 -17.515 70.205 ;
        RECT -17.845 68.515 -17.515 68.845 ;
        RECT -17.845 67.155 -17.515 67.485 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.085 132.52 -29.755 133.65 ;
        RECT -30.085 128.355 -29.755 128.685 ;
        RECT -30.085 126.995 -29.755 127.325 ;
        RECT -30.085 125.635 -29.755 125.965 ;
        RECT -30.085 124.275 -29.755 124.605 ;
        RECT -30.085 122.915 -29.755 123.245 ;
        RECT -30.085 121.555 -29.755 121.885 ;
        RECT -30.085 120.195 -29.755 120.525 ;
        RECT -30.085 118.835 -29.755 119.165 ;
        RECT -30.085 117.475 -29.755 117.805 ;
        RECT -30.085 116.115 -29.755 116.445 ;
        RECT -30.085 114.755 -29.755 115.085 ;
        RECT -30.085 113.395 -29.755 113.725 ;
        RECT -30.085 112.035 -29.755 112.365 ;
        RECT -30.085 110.675 -29.755 111.005 ;
        RECT -30.085 109.315 -29.755 109.645 ;
        RECT -30.085 107.955 -29.755 108.285 ;
        RECT -30.085 106.595 -29.755 106.925 ;
        RECT -30.085 105.235 -29.755 105.565 ;
        RECT -30.085 103.875 -29.755 104.205 ;
        RECT -30.085 102.515 -29.755 102.845 ;
        RECT -30.085 101.155 -29.755 101.485 ;
        RECT -30.085 99.795 -29.755 100.125 ;
        RECT -30.085 98.435 -29.755 98.765 ;
        RECT -30.085 97.075 -29.755 97.405 ;
        RECT -30.085 95.715 -29.755 96.045 ;
        RECT -30.085 94.355 -29.755 94.685 ;
        RECT -30.085 92.995 -29.755 93.325 ;
        RECT -30.085 91.635 -29.755 91.965 ;
        RECT -30.085 90.275 -29.755 90.605 ;
        RECT -30.085 88.915 -29.755 89.245 ;
        RECT -30.085 87.555 -29.755 87.885 ;
        RECT -30.085 86.195 -29.755 86.525 ;
        RECT -30.085 84.835 -29.755 85.165 ;
        RECT -30.085 83.475 -29.755 83.805 ;
        RECT -30.085 82.115 -29.755 82.445 ;
        RECT -30.085 80.755 -29.755 81.085 ;
        RECT -30.085 79.395 -29.755 79.725 ;
        RECT -30.085 78.035 -29.755 78.365 ;
        RECT -30.085 76.675 -29.755 77.005 ;
        RECT -30.085 75.315 -29.755 75.645 ;
        RECT -30.085 73.955 -29.755 74.285 ;
        RECT -30.085 72.595 -29.755 72.925 ;
        RECT -30.085 71.235 -29.755 71.565 ;
        RECT -30.085 69.875 -29.755 70.205 ;
        RECT -30.085 68.515 -29.755 68.845 ;
        RECT -30.085 67.155 -29.755 67.485 ;
        RECT -30.085 65.795 -29.755 66.125 ;
        RECT -30.085 64.435 -29.755 64.765 ;
        RECT -30.085 63.075 -29.755 63.405 ;
        RECT -30.085 61.715 -29.755 62.045 ;
        RECT -30.085 60.355 -29.755 60.685 ;
        RECT -30.085 58.995 -29.755 59.325 ;
        RECT -30.085 57.635 -29.755 57.965 ;
        RECT -30.085 56.275 -29.755 56.605 ;
        RECT -30.085 54.915 -29.755 55.245 ;
        RECT -30.085 53.555 -29.755 53.885 ;
        RECT -30.085 52.195 -29.755 52.525 ;
        RECT -30.085 50.835 -29.755 51.165 ;
        RECT -30.085 49.475 -29.755 49.805 ;
        RECT -30.085 48.115 -29.755 48.445 ;
        RECT -30.085 46.755 -29.755 47.085 ;
        RECT -30.085 45.395 -29.755 45.725 ;
        RECT -30.085 44.035 -29.755 44.365 ;
        RECT -30.085 42.675 -29.755 43.005 ;
        RECT -30.085 41.315 -29.755 41.645 ;
        RECT -30.085 39.955 -29.755 40.285 ;
        RECT -30.085 38.595 -29.755 38.925 ;
        RECT -30.085 37.235 -29.755 37.565 ;
        RECT -30.085 35.875 -29.755 36.205 ;
        RECT -30.085 34.515 -29.755 34.845 ;
        RECT -30.085 33.155 -29.755 33.485 ;
        RECT -30.085 31.795 -29.755 32.125 ;
        RECT -30.085 30.435 -29.755 30.765 ;
        RECT -30.085 29.075 -29.755 29.405 ;
        RECT -30.085 27.715 -29.755 28.045 ;
        RECT -30.085 26.355 -29.755 26.685 ;
        RECT -30.085 24.995 -29.755 25.325 ;
        RECT -30.085 23.635 -29.755 23.965 ;
        RECT -30.085 22.275 -29.755 22.605 ;
        RECT -30.085 20.915 -29.755 21.245 ;
        RECT -30.085 19.555 -29.755 19.885 ;
        RECT -30.085 18.195 -29.755 18.525 ;
        RECT -30.085 16.835 -29.755 17.165 ;
        RECT -30.085 15.475 -29.755 15.805 ;
        RECT -30.085 14.115 -29.755 14.445 ;
        RECT -30.085 12.755 -29.755 13.085 ;
        RECT -30.085 11.395 -29.755 11.725 ;
        RECT -30.085 10.035 -29.755 10.365 ;
        RECT -30.085 8.675 -29.755 9.005 ;
        RECT -30.085 7.315 -29.755 7.645 ;
        RECT -30.085 5.955 -29.755 6.285 ;
        RECT -30.085 4.595 -29.755 4.925 ;
        RECT -30.085 3.235 -29.755 3.565 ;
        RECT -30.085 1.875 -29.755 2.205 ;
        RECT -30.085 0.515 -29.755 0.845 ;
        RECT -30.085 -7.645 -29.755 -7.315 ;
        RECT -30.085 -9.005 -29.755 -8.675 ;
        RECT -30.085 -13.085 -29.755 -12.755 ;
        RECT -30.085 -17.165 -29.755 -16.835 ;
        RECT -30.085 -26.685 -29.755 -26.355 ;
        RECT -30.085 -29.405 -29.755 -29.075 ;
        RECT -30.085 -43.005 -29.755 -42.675 ;
        RECT -30.085 -44.365 -29.755 -44.035 ;
        RECT -30.085 -45.725 -29.755 -45.395 ;
        RECT -30.085 -47.085 -29.755 -46.755 ;
        RECT -30.085 -48.445 -29.755 -48.115 ;
        RECT -30.085 -49.805 -29.755 -49.475 ;
        RECT -30.085 -51.165 -29.755 -50.835 ;
        RECT -30.085 -52.525 -29.755 -52.195 ;
        RECT -30.085 -53.885 -29.755 -53.555 ;
        RECT -30.085 -55.245 -29.755 -54.915 ;
        RECT -30.085 -56.605 -29.755 -56.275 ;
        RECT -30.085 -57.965 -29.755 -57.635 ;
        RECT -30.085 -59.325 -29.755 -58.995 ;
        RECT -30.085 -60.685 -29.755 -60.355 ;
        RECT -30.085 -62.045 -29.755 -61.715 ;
        RECT -30.085 -63.405 -29.755 -63.075 ;
        RECT -30.085 -64.765 -29.755 -64.435 ;
        RECT -30.085 -66.125 -29.755 -65.795 ;
        RECT -30.085 -67.485 -29.755 -67.155 ;
        RECT -30.085 -68.845 -29.755 -68.515 ;
        RECT -30.085 -70.205 -29.755 -69.875 ;
        RECT -30.085 -71.565 -29.755 -71.235 ;
        RECT -30.085 -72.925 -29.755 -72.595 ;
        RECT -30.085 -74.285 -29.755 -73.955 ;
        RECT -30.085 -75.645 -29.755 -75.315 ;
        RECT -30.085 -77.005 -29.755 -76.675 ;
        RECT -30.085 -78.365 -29.755 -78.035 ;
        RECT -30.085 -79.725 -29.755 -79.395 ;
        RECT -30.085 -81.085 -29.755 -80.755 ;
        RECT -30.085 -82.445 -29.755 -82.115 ;
        RECT -30.085 -83.805 -29.755 -83.475 ;
        RECT -30.085 -85.165 -29.755 -84.835 ;
        RECT -30.085 -86.525 -29.755 -86.195 ;
        RECT -30.085 -87.885 -29.755 -87.555 ;
        RECT -30.085 -89.245 -29.755 -88.915 ;
        RECT -30.085 -90.605 -29.755 -90.275 ;
        RECT -30.085 -91.965 -29.755 -91.635 ;
        RECT -30.085 -93.325 -29.755 -92.995 ;
        RECT -30.085 -94.685 -29.755 -94.355 ;
        RECT -30.085 -96.045 -29.755 -95.715 ;
        RECT -30.085 -97.405 -29.755 -97.075 ;
        RECT -30.085 -98.765 -29.755 -98.435 ;
        RECT -30.085 -100.125 -29.755 -99.795 ;
        RECT -30.085 -101.485 -29.755 -101.155 ;
        RECT -30.085 -102.845 -29.755 -102.515 ;
        RECT -30.085 -104.205 -29.755 -103.875 ;
        RECT -30.085 -105.565 -29.755 -105.235 ;
        RECT -30.085 -109.645 -29.755 -109.315 ;
        RECT -30.085 -111.005 -29.755 -110.675 ;
        RECT -30.085 -111.87 -29.755 -111.54 ;
        RECT -30.085 -113.725 -29.755 -113.395 ;
        RECT -30.085 -115.085 -29.755 -114.755 ;
        RECT -30.085 -116.445 -29.755 -116.115 ;
        RECT -30.085 -117.805 -29.755 -117.475 ;
        RECT -30.085 -120.525 -29.755 -120.195 ;
        RECT -30.085 -121.885 -29.755 -121.555 ;
        RECT -30.085 -123.245 -29.755 -122.915 ;
        RECT -30.085 -124.71 -29.755 -124.38 ;
        RECT -30.085 -125.965 -29.755 -125.635 ;
        RECT -30.085 -127.325 -29.755 -126.995 ;
        RECT -30.085 -130.045 -29.755 -129.715 ;
        RECT -30.08 -132.08 -29.76 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.085 -214.365 -29.755 -214.035 ;
        RECT -30.085 -215.725 -29.755 -215.395 ;
        RECT -30.085 -217.085 -29.755 -216.755 ;
        RECT -30.085 -218.445 -29.755 -218.115 ;
        RECT -30.085 -224.09 -29.755 -222.96 ;
        RECT -30.08 -224.205 -29.76 -210.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -28.725 132.52 -28.395 133.65 ;
        RECT -28.725 128.355 -28.395 128.685 ;
        RECT -28.725 126.995 -28.395 127.325 ;
        RECT -28.725 125.635 -28.395 125.965 ;
        RECT -28.725 124.275 -28.395 124.605 ;
        RECT -28.725 122.915 -28.395 123.245 ;
        RECT -28.725 121.555 -28.395 121.885 ;
        RECT -28.725 120.195 -28.395 120.525 ;
        RECT -28.725 118.835 -28.395 119.165 ;
        RECT -28.725 117.475 -28.395 117.805 ;
        RECT -28.725 116.115 -28.395 116.445 ;
        RECT -28.725 114.755 -28.395 115.085 ;
        RECT -28.725 113.395 -28.395 113.725 ;
        RECT -28.725 112.035 -28.395 112.365 ;
        RECT -28.725 110.675 -28.395 111.005 ;
        RECT -28.725 109.315 -28.395 109.645 ;
        RECT -28.725 107.955 -28.395 108.285 ;
        RECT -28.725 106.595 -28.395 106.925 ;
        RECT -28.725 105.235 -28.395 105.565 ;
        RECT -28.725 103.875 -28.395 104.205 ;
        RECT -28.725 102.515 -28.395 102.845 ;
        RECT -28.725 101.155 -28.395 101.485 ;
        RECT -28.725 99.795 -28.395 100.125 ;
        RECT -28.725 98.435 -28.395 98.765 ;
        RECT -28.725 97.075 -28.395 97.405 ;
        RECT -28.725 95.715 -28.395 96.045 ;
        RECT -28.725 94.355 -28.395 94.685 ;
        RECT -28.725 92.995 -28.395 93.325 ;
        RECT -28.725 91.635 -28.395 91.965 ;
        RECT -28.725 90.275 -28.395 90.605 ;
        RECT -28.725 88.915 -28.395 89.245 ;
        RECT -28.725 87.555 -28.395 87.885 ;
        RECT -28.725 86.195 -28.395 86.525 ;
        RECT -28.725 84.835 -28.395 85.165 ;
        RECT -28.725 83.475 -28.395 83.805 ;
        RECT -28.725 82.115 -28.395 82.445 ;
        RECT -28.725 80.755 -28.395 81.085 ;
        RECT -28.725 79.395 -28.395 79.725 ;
        RECT -28.725 78.035 -28.395 78.365 ;
        RECT -28.725 76.675 -28.395 77.005 ;
        RECT -28.725 75.315 -28.395 75.645 ;
        RECT -28.725 73.955 -28.395 74.285 ;
        RECT -28.725 72.595 -28.395 72.925 ;
        RECT -28.725 71.235 -28.395 71.565 ;
        RECT -28.725 69.875 -28.395 70.205 ;
        RECT -28.725 68.515 -28.395 68.845 ;
        RECT -28.725 67.155 -28.395 67.485 ;
        RECT -28.725 65.795 -28.395 66.125 ;
        RECT -28.725 64.435 -28.395 64.765 ;
        RECT -28.725 63.075 -28.395 63.405 ;
        RECT -28.725 61.715 -28.395 62.045 ;
        RECT -28.725 60.355 -28.395 60.685 ;
        RECT -28.725 58.995 -28.395 59.325 ;
        RECT -28.725 57.635 -28.395 57.965 ;
        RECT -28.725 56.275 -28.395 56.605 ;
        RECT -28.725 54.915 -28.395 55.245 ;
        RECT -28.725 53.555 -28.395 53.885 ;
        RECT -28.725 52.195 -28.395 52.525 ;
        RECT -28.725 50.835 -28.395 51.165 ;
        RECT -28.725 49.475 -28.395 49.805 ;
        RECT -28.725 48.115 -28.395 48.445 ;
        RECT -28.725 46.755 -28.395 47.085 ;
        RECT -28.725 45.395 -28.395 45.725 ;
        RECT -28.725 44.035 -28.395 44.365 ;
        RECT -28.725 42.675 -28.395 43.005 ;
        RECT -28.725 41.315 -28.395 41.645 ;
        RECT -28.725 39.955 -28.395 40.285 ;
        RECT -28.725 38.595 -28.395 38.925 ;
        RECT -28.725 37.235 -28.395 37.565 ;
        RECT -28.725 35.875 -28.395 36.205 ;
        RECT -28.725 34.515 -28.395 34.845 ;
        RECT -28.725 33.155 -28.395 33.485 ;
        RECT -28.725 31.795 -28.395 32.125 ;
        RECT -28.725 30.435 -28.395 30.765 ;
        RECT -28.725 29.075 -28.395 29.405 ;
        RECT -28.725 27.715 -28.395 28.045 ;
        RECT -28.725 26.355 -28.395 26.685 ;
        RECT -28.725 24.995 -28.395 25.325 ;
        RECT -28.725 23.635 -28.395 23.965 ;
        RECT -28.725 22.275 -28.395 22.605 ;
        RECT -28.725 20.915 -28.395 21.245 ;
        RECT -28.725 19.555 -28.395 19.885 ;
        RECT -28.725 18.195 -28.395 18.525 ;
        RECT -28.725 16.835 -28.395 17.165 ;
        RECT -28.725 15.475 -28.395 15.805 ;
        RECT -28.725 14.115 -28.395 14.445 ;
        RECT -28.725 12.755 -28.395 13.085 ;
        RECT -28.725 11.395 -28.395 11.725 ;
        RECT -28.725 10.035 -28.395 10.365 ;
        RECT -28.725 8.675 -28.395 9.005 ;
        RECT -28.725 7.315 -28.395 7.645 ;
        RECT -28.725 5.955 -28.395 6.285 ;
        RECT -28.725 4.595 -28.395 4.925 ;
        RECT -28.725 3.235 -28.395 3.565 ;
        RECT -28.725 1.875 -28.395 2.205 ;
        RECT -28.725 0.515 -28.395 0.845 ;
        RECT -28.725 -6.94 -28.395 -6.61 ;
        RECT -28.725 -7.645 -28.395 -7.315 ;
        RECT -28.725 -9.005 -28.395 -8.675 ;
        RECT -28.725 -13.085 -28.395 -12.755 ;
        RECT -28.725 -14.13 -28.395 -13.8 ;
        RECT -28.725 -17.165 -28.395 -16.835 ;
        RECT -28.725 -26.685 -28.395 -26.355 ;
        RECT -28.725 -28.12 -28.395 -27.79 ;
        RECT -28.725 -29.405 -28.395 -29.075 ;
        RECT -28.725 -35.31 -28.395 -34.98 ;
        RECT -28.725 -43.005 -28.395 -42.675 ;
        RECT -28.725 -44.365 -28.395 -44.035 ;
        RECT -28.725 -45.725 -28.395 -45.395 ;
        RECT -28.725 -47.085 -28.395 -46.755 ;
        RECT -28.725 -48.445 -28.395 -48.115 ;
        RECT -28.725 -49.805 -28.395 -49.475 ;
        RECT -28.725 -51.165 -28.395 -50.835 ;
        RECT -28.725 -52.525 -28.395 -52.195 ;
        RECT -28.725 -53.885 -28.395 -53.555 ;
        RECT -28.725 -55.245 -28.395 -54.915 ;
        RECT -28.725 -56.605 -28.395 -56.275 ;
        RECT -28.725 -57.965 -28.395 -57.635 ;
        RECT -28.725 -59.325 -28.395 -58.995 ;
        RECT -28.725 -60.685 -28.395 -60.355 ;
        RECT -28.725 -62.045 -28.395 -61.715 ;
        RECT -28.725 -63.405 -28.395 -63.075 ;
        RECT -28.725 -64.765 -28.395 -64.435 ;
        RECT -28.725 -66.125 -28.395 -65.795 ;
        RECT -28.725 -67.485 -28.395 -67.155 ;
        RECT -28.725 -68.845 -28.395 -68.515 ;
        RECT -28.725 -70.205 -28.395 -69.875 ;
        RECT -28.725 -71.565 -28.395 -71.235 ;
        RECT -28.725 -72.925 -28.395 -72.595 ;
        RECT -28.725 -74.285 -28.395 -73.955 ;
        RECT -28.725 -75.645 -28.395 -75.315 ;
        RECT -28.725 -77.005 -28.395 -76.675 ;
        RECT -28.725 -78.365 -28.395 -78.035 ;
        RECT -28.725 -79.725 -28.395 -79.395 ;
        RECT -28.725 -81.085 -28.395 -80.755 ;
        RECT -28.725 -82.445 -28.395 -82.115 ;
        RECT -28.725 -83.805 -28.395 -83.475 ;
        RECT -28.725 -85.165 -28.395 -84.835 ;
        RECT -28.725 -86.525 -28.395 -86.195 ;
        RECT -28.725 -87.885 -28.395 -87.555 ;
        RECT -28.725 -89.245 -28.395 -88.915 ;
        RECT -28.725 -90.605 -28.395 -90.275 ;
        RECT -28.725 -91.965 -28.395 -91.635 ;
        RECT -28.725 -93.325 -28.395 -92.995 ;
        RECT -28.725 -94.685 -28.395 -94.355 ;
        RECT -28.725 -96.045 -28.395 -95.715 ;
        RECT -28.725 -97.405 -28.395 -97.075 ;
        RECT -28.725 -98.765 -28.395 -98.435 ;
        RECT -28.725 -100.125 -28.395 -99.795 ;
        RECT -28.725 -101.485 -28.395 -101.155 ;
        RECT -28.725 -102.845 -28.395 -102.515 ;
        RECT -28.725 -104.205 -28.395 -103.875 ;
        RECT -28.725 -109.645 -28.395 -109.315 ;
        RECT -28.725 -111.005 -28.395 -110.675 ;
        RECT -28.725 -111.87 -28.395 -111.54 ;
        RECT -28.725 -113.725 -28.395 -113.395 ;
        RECT -28.725 -115.085 -28.395 -114.755 ;
        RECT -28.725 -116.445 -28.395 -116.115 ;
        RECT -28.725 -117.805 -28.395 -117.475 ;
        RECT -28.725 -120.525 -28.395 -120.195 ;
        RECT -28.725 -121.885 -28.395 -121.555 ;
        RECT -28.725 -123.245 -28.395 -122.915 ;
        RECT -28.725 -124.71 -28.395 -124.38 ;
        RECT -28.725 -125.965 -28.395 -125.635 ;
        RECT -28.725 -127.325 -28.395 -126.995 ;
        RECT -28.725 -130.045 -28.395 -129.715 ;
        RECT -28.725 -132.765 -28.395 -132.435 ;
        RECT -28.725 -134.125 -28.395 -133.795 ;
        RECT -28.725 -135.485 -28.395 -135.155 ;
        RECT -28.725 -136.845 -28.395 -136.515 ;
        RECT -28.725 -138.205 -28.395 -137.875 ;
        RECT -28.725 -139.565 -28.395 -139.235 ;
        RECT -28.725 -142.285 -28.395 -141.955 ;
        RECT -28.725 -143.645 -28.395 -143.315 ;
        RECT -28.725 -145.005 -28.395 -144.675 ;
        RECT -28.725 -146.365 -28.395 -146.035 ;
        RECT -28.725 -147.725 -28.395 -147.395 ;
        RECT -28.725 -149.085 -28.395 -148.755 ;
        RECT -28.725 -150.445 -28.395 -150.115 ;
        RECT -28.725 -151.805 -28.395 -151.475 ;
        RECT -28.725 -153.165 -28.395 -152.835 ;
        RECT -28.725 -154.525 -28.395 -154.195 ;
        RECT -28.725 -155.885 -28.395 -155.555 ;
        RECT -28.725 -157.245 -28.395 -156.915 ;
        RECT -28.725 -158.605 -28.395 -158.275 ;
        RECT -28.725 -159.965 -28.395 -159.635 ;
        RECT -28.725 -161.325 -28.395 -160.995 ;
        RECT -28.725 -162.685 -28.395 -162.355 ;
        RECT -28.725 -164.045 -28.395 -163.715 ;
        RECT -28.725 -165.405 -28.395 -165.075 ;
        RECT -28.725 -166.765 -28.395 -166.435 ;
        RECT -28.725 -170.845 -28.395 -170.515 ;
        RECT -28.725 -172.205 -28.395 -171.875 ;
        RECT -28.725 -173.565 -28.395 -173.235 ;
        RECT -28.725 -174.925 -28.395 -174.595 ;
        RECT -28.725 -176.285 -28.395 -175.955 ;
        RECT -28.725 -179.005 -28.395 -178.675 ;
        RECT -28.725 -180.365 -28.395 -180.035 ;
        RECT -28.725 -181.725 -28.395 -181.395 ;
        RECT -28.725 -183.085 -28.395 -182.755 ;
        RECT -28.725 -184.445 -28.395 -184.115 ;
        RECT -28.725 -185.805 -28.395 -185.475 ;
        RECT -28.725 -188.525 -28.395 -188.195 ;
        RECT -28.725 -189.885 -28.395 -189.555 ;
        RECT -28.725 -195.325 -28.395 -194.995 ;
        RECT -28.725 -196.685 -28.395 -196.355 ;
        RECT -28.725 -198.045 -28.395 -197.715 ;
        RECT -28.725 -199.405 -28.395 -199.075 ;
        RECT -28.725 -200.765 -28.395 -200.435 ;
        RECT -28.725 -202.125 -28.395 -201.795 ;
        RECT -28.725 -203.485 -28.395 -203.155 ;
        RECT -28.725 -204.845 -28.395 -204.515 ;
        RECT -28.725 -207.565 -28.395 -207.235 ;
        RECT -28.725 -208.925 -28.395 -208.595 ;
        RECT -28.725 -211.645 -28.395 -211.315 ;
        RECT -28.725 -214.365 -28.395 -214.035 ;
        RECT -28.725 -215.725 -28.395 -215.395 ;
        RECT -28.725 -217.085 -28.395 -216.755 ;
        RECT -28.725 -218.445 -28.395 -218.115 ;
        RECT -28.725 -224.09 -28.395 -222.96 ;
        RECT -28.72 -224.205 -28.4 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -27.365 132.52 -27.035 133.65 ;
        RECT -27.365 128.355 -27.035 128.685 ;
        RECT -27.365 126.995 -27.035 127.325 ;
        RECT -27.365 125.635 -27.035 125.965 ;
        RECT -27.365 124.275 -27.035 124.605 ;
        RECT -27.365 122.915 -27.035 123.245 ;
        RECT -27.365 121.555 -27.035 121.885 ;
        RECT -27.365 120.195 -27.035 120.525 ;
        RECT -27.365 118.835 -27.035 119.165 ;
        RECT -27.365 117.475 -27.035 117.805 ;
        RECT -27.365 116.115 -27.035 116.445 ;
        RECT -27.365 114.755 -27.035 115.085 ;
        RECT -27.365 113.395 -27.035 113.725 ;
        RECT -27.365 112.035 -27.035 112.365 ;
        RECT -27.365 110.675 -27.035 111.005 ;
        RECT -27.365 109.315 -27.035 109.645 ;
        RECT -27.365 107.955 -27.035 108.285 ;
        RECT -27.365 106.595 -27.035 106.925 ;
        RECT -27.365 105.235 -27.035 105.565 ;
        RECT -27.365 103.875 -27.035 104.205 ;
        RECT -27.365 102.515 -27.035 102.845 ;
        RECT -27.365 101.155 -27.035 101.485 ;
        RECT -27.365 99.795 -27.035 100.125 ;
        RECT -27.365 98.435 -27.035 98.765 ;
        RECT -27.365 97.075 -27.035 97.405 ;
        RECT -27.365 95.715 -27.035 96.045 ;
        RECT -27.365 94.355 -27.035 94.685 ;
        RECT -27.365 92.995 -27.035 93.325 ;
        RECT -27.365 91.635 -27.035 91.965 ;
        RECT -27.365 90.275 -27.035 90.605 ;
        RECT -27.365 88.915 -27.035 89.245 ;
        RECT -27.365 87.555 -27.035 87.885 ;
        RECT -27.365 86.195 -27.035 86.525 ;
        RECT -27.365 84.835 -27.035 85.165 ;
        RECT -27.365 83.475 -27.035 83.805 ;
        RECT -27.365 82.115 -27.035 82.445 ;
        RECT -27.365 80.755 -27.035 81.085 ;
        RECT -27.365 79.395 -27.035 79.725 ;
        RECT -27.365 78.035 -27.035 78.365 ;
        RECT -27.365 76.675 -27.035 77.005 ;
        RECT -27.365 75.315 -27.035 75.645 ;
        RECT -27.365 73.955 -27.035 74.285 ;
        RECT -27.365 72.595 -27.035 72.925 ;
        RECT -27.365 71.235 -27.035 71.565 ;
        RECT -27.365 69.875 -27.035 70.205 ;
        RECT -27.365 68.515 -27.035 68.845 ;
        RECT -27.365 67.155 -27.035 67.485 ;
        RECT -27.365 65.795 -27.035 66.125 ;
        RECT -27.365 64.435 -27.035 64.765 ;
        RECT -27.365 63.075 -27.035 63.405 ;
        RECT -27.365 61.715 -27.035 62.045 ;
        RECT -27.365 60.355 -27.035 60.685 ;
        RECT -27.365 58.995 -27.035 59.325 ;
        RECT -27.365 57.635 -27.035 57.965 ;
        RECT -27.365 56.275 -27.035 56.605 ;
        RECT -27.365 54.915 -27.035 55.245 ;
        RECT -27.365 53.555 -27.035 53.885 ;
        RECT -27.365 52.195 -27.035 52.525 ;
        RECT -27.365 50.835 -27.035 51.165 ;
        RECT -27.365 49.475 -27.035 49.805 ;
        RECT -27.365 48.115 -27.035 48.445 ;
        RECT -27.365 46.755 -27.035 47.085 ;
        RECT -27.365 45.395 -27.035 45.725 ;
        RECT -27.365 44.035 -27.035 44.365 ;
        RECT -27.365 42.675 -27.035 43.005 ;
        RECT -27.365 41.315 -27.035 41.645 ;
        RECT -27.365 39.955 -27.035 40.285 ;
        RECT -27.365 38.595 -27.035 38.925 ;
        RECT -27.365 37.235 -27.035 37.565 ;
        RECT -27.365 35.875 -27.035 36.205 ;
        RECT -27.365 34.515 -27.035 34.845 ;
        RECT -27.365 33.155 -27.035 33.485 ;
        RECT -27.365 31.795 -27.035 32.125 ;
        RECT -27.365 30.435 -27.035 30.765 ;
        RECT -27.365 29.075 -27.035 29.405 ;
        RECT -27.365 27.715 -27.035 28.045 ;
        RECT -27.365 26.355 -27.035 26.685 ;
        RECT -27.365 24.995 -27.035 25.325 ;
        RECT -27.365 23.635 -27.035 23.965 ;
        RECT -27.365 22.275 -27.035 22.605 ;
        RECT -27.365 20.915 -27.035 21.245 ;
        RECT -27.365 19.555 -27.035 19.885 ;
        RECT -27.365 18.195 -27.035 18.525 ;
        RECT -27.365 16.835 -27.035 17.165 ;
        RECT -27.365 15.475 -27.035 15.805 ;
        RECT -27.365 14.115 -27.035 14.445 ;
        RECT -27.365 12.755 -27.035 13.085 ;
        RECT -27.365 11.395 -27.035 11.725 ;
        RECT -27.365 10.035 -27.035 10.365 ;
        RECT -27.365 8.675 -27.035 9.005 ;
        RECT -27.365 7.315 -27.035 7.645 ;
        RECT -27.365 5.955 -27.035 6.285 ;
        RECT -27.365 4.595 -27.035 4.925 ;
        RECT -27.365 3.235 -27.035 3.565 ;
        RECT -27.365 1.875 -27.035 2.205 ;
        RECT -27.365 0.515 -27.035 0.845 ;
        RECT -27.365 -6.94 -27.035 -6.61 ;
        RECT -27.365 -7.645 -27.035 -7.315 ;
        RECT -27.365 -9.005 -27.035 -8.675 ;
        RECT -27.365 -13.085 -27.035 -12.755 ;
        RECT -27.365 -14.13 -27.035 -13.8 ;
        RECT -27.365 -17.165 -27.035 -16.835 ;
        RECT -27.365 -26.685 -27.035 -26.355 ;
        RECT -27.365 -28.12 -27.035 -27.79 ;
        RECT -27.365 -29.405 -27.035 -29.075 ;
        RECT -27.365 -35.31 -27.035 -34.98 ;
        RECT -27.365 -43.005 -27.035 -42.675 ;
        RECT -27.365 -44.365 -27.035 -44.035 ;
        RECT -27.365 -45.725 -27.035 -45.395 ;
        RECT -27.365 -47.085 -27.035 -46.755 ;
        RECT -27.365 -48.445 -27.035 -48.115 ;
        RECT -27.365 -49.805 -27.035 -49.475 ;
        RECT -27.365 -51.165 -27.035 -50.835 ;
        RECT -27.365 -52.525 -27.035 -52.195 ;
        RECT -27.365 -53.885 -27.035 -53.555 ;
        RECT -27.365 -55.245 -27.035 -54.915 ;
        RECT -27.365 -56.605 -27.035 -56.275 ;
        RECT -27.365 -57.965 -27.035 -57.635 ;
        RECT -27.365 -59.325 -27.035 -58.995 ;
        RECT -27.365 -60.685 -27.035 -60.355 ;
        RECT -27.365 -62.045 -27.035 -61.715 ;
        RECT -27.365 -63.405 -27.035 -63.075 ;
        RECT -27.365 -64.765 -27.035 -64.435 ;
        RECT -27.365 -66.125 -27.035 -65.795 ;
        RECT -27.365 -67.485 -27.035 -67.155 ;
        RECT -27.365 -68.845 -27.035 -68.515 ;
        RECT -27.365 -70.205 -27.035 -69.875 ;
        RECT -27.365 -71.565 -27.035 -71.235 ;
        RECT -27.365 -72.925 -27.035 -72.595 ;
        RECT -27.365 -74.285 -27.035 -73.955 ;
        RECT -27.365 -75.645 -27.035 -75.315 ;
        RECT -27.365 -77.005 -27.035 -76.675 ;
        RECT -27.365 -78.365 -27.035 -78.035 ;
        RECT -27.365 -79.725 -27.035 -79.395 ;
        RECT -27.365 -81.085 -27.035 -80.755 ;
        RECT -27.365 -82.445 -27.035 -82.115 ;
        RECT -27.365 -83.805 -27.035 -83.475 ;
        RECT -27.365 -85.165 -27.035 -84.835 ;
        RECT -27.365 -86.525 -27.035 -86.195 ;
        RECT -27.365 -87.885 -27.035 -87.555 ;
        RECT -27.365 -89.245 -27.035 -88.915 ;
        RECT -27.365 -90.605 -27.035 -90.275 ;
        RECT -27.365 -91.965 -27.035 -91.635 ;
        RECT -27.365 -93.325 -27.035 -92.995 ;
        RECT -27.365 -94.685 -27.035 -94.355 ;
        RECT -27.365 -96.045 -27.035 -95.715 ;
        RECT -27.365 -97.405 -27.035 -97.075 ;
        RECT -27.365 -98.765 -27.035 -98.435 ;
        RECT -27.365 -100.125 -27.035 -99.795 ;
        RECT -27.365 -101.485 -27.035 -101.155 ;
        RECT -27.365 -102.845 -27.035 -102.515 ;
        RECT -27.365 -104.205 -27.035 -103.875 ;
        RECT -27.365 -109.645 -27.035 -109.315 ;
        RECT -27.365 -111.005 -27.035 -110.675 ;
        RECT -27.365 -111.87 -27.035 -111.54 ;
        RECT -27.365 -113.725 -27.035 -113.395 ;
        RECT -27.365 -115.085 -27.035 -114.755 ;
        RECT -27.365 -116.445 -27.035 -116.115 ;
        RECT -27.365 -117.805 -27.035 -117.475 ;
        RECT -27.365 -120.525 -27.035 -120.195 ;
        RECT -27.365 -121.885 -27.035 -121.555 ;
        RECT -27.365 -123.245 -27.035 -122.915 ;
        RECT -27.365 -124.71 -27.035 -124.38 ;
        RECT -27.365 -125.965 -27.035 -125.635 ;
        RECT -27.365 -127.325 -27.035 -126.995 ;
        RECT -27.365 -130.045 -27.035 -129.715 ;
        RECT -27.365 -132.765 -27.035 -132.435 ;
        RECT -27.365 -134.125 -27.035 -133.795 ;
        RECT -27.365 -135.485 -27.035 -135.155 ;
        RECT -27.365 -136.845 -27.035 -136.515 ;
        RECT -27.365 -138.205 -27.035 -137.875 ;
        RECT -27.365 -139.565 -27.035 -139.235 ;
        RECT -27.365 -142.285 -27.035 -141.955 ;
        RECT -27.365 -143.645 -27.035 -143.315 ;
        RECT -27.365 -145.005 -27.035 -144.675 ;
        RECT -27.365 -146.365 -27.035 -146.035 ;
        RECT -27.365 -147.725 -27.035 -147.395 ;
        RECT -27.365 -149.085 -27.035 -148.755 ;
        RECT -27.365 -150.445 -27.035 -150.115 ;
        RECT -27.365 -151.805 -27.035 -151.475 ;
        RECT -27.365 -153.165 -27.035 -152.835 ;
        RECT -27.365 -154.525 -27.035 -154.195 ;
        RECT -27.365 -155.885 -27.035 -155.555 ;
        RECT -27.365 -157.245 -27.035 -156.915 ;
        RECT -27.365 -158.605 -27.035 -158.275 ;
        RECT -27.365 -159.965 -27.035 -159.635 ;
        RECT -27.365 -161.325 -27.035 -160.995 ;
        RECT -27.365 -162.685 -27.035 -162.355 ;
        RECT -27.365 -165.405 -27.035 -165.075 ;
        RECT -27.365 -166.765 -27.035 -166.435 ;
        RECT -27.365 -170.845 -27.035 -170.515 ;
        RECT -27.365 -172.205 -27.035 -171.875 ;
        RECT -27.365 -173.565 -27.035 -173.235 ;
        RECT -27.365 -174.925 -27.035 -174.595 ;
        RECT -27.365 -176.285 -27.035 -175.955 ;
        RECT -27.365 -179.005 -27.035 -178.675 ;
        RECT -27.365 -180.365 -27.035 -180.035 ;
        RECT -27.365 -181.725 -27.035 -181.395 ;
        RECT -27.365 -183.085 -27.035 -182.755 ;
        RECT -27.365 -184.445 -27.035 -184.115 ;
        RECT -27.365 -185.805 -27.035 -185.475 ;
        RECT -27.365 -188.525 -27.035 -188.195 ;
        RECT -27.365 -189.885 -27.035 -189.555 ;
        RECT -27.365 -195.325 -27.035 -194.995 ;
        RECT -27.365 -196.685 -27.035 -196.355 ;
        RECT -27.365 -198.045 -27.035 -197.715 ;
        RECT -27.365 -199.405 -27.035 -199.075 ;
        RECT -27.365 -200.765 -27.035 -200.435 ;
        RECT -27.365 -202.125 -27.035 -201.795 ;
        RECT -27.365 -203.485 -27.035 -203.155 ;
        RECT -27.365 -204.845 -27.035 -204.515 ;
        RECT -27.365 -206.555 -27.035 -206.225 ;
        RECT -27.365 -207.565 -27.035 -207.235 ;
        RECT -27.365 -208.925 -27.035 -208.595 ;
        RECT -27.365 -211.645 -27.035 -211.315 ;
        RECT -27.365 -214.365 -27.035 -214.035 ;
        RECT -27.365 -215.725 -27.035 -215.395 ;
        RECT -27.365 -217.085 -27.035 -216.755 ;
        RECT -27.365 -218.445 -27.035 -218.115 ;
        RECT -27.365 -224.09 -27.035 -222.96 ;
        RECT -27.36 -224.205 -27.04 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.005 132.52 -25.675 133.65 ;
        RECT -26.005 128.355 -25.675 128.685 ;
        RECT -26.005 126.995 -25.675 127.325 ;
        RECT -26.005 125.635 -25.675 125.965 ;
        RECT -26.005 124.275 -25.675 124.605 ;
        RECT -26.005 122.915 -25.675 123.245 ;
        RECT -26.005 121.555 -25.675 121.885 ;
        RECT -26.005 120.195 -25.675 120.525 ;
        RECT -26.005 118.835 -25.675 119.165 ;
        RECT -26.005 117.475 -25.675 117.805 ;
        RECT -26.005 116.115 -25.675 116.445 ;
        RECT -26.005 114.755 -25.675 115.085 ;
        RECT -26.005 113.395 -25.675 113.725 ;
        RECT -26.005 112.035 -25.675 112.365 ;
        RECT -26.005 110.675 -25.675 111.005 ;
        RECT -26.005 109.315 -25.675 109.645 ;
        RECT -26.005 107.955 -25.675 108.285 ;
        RECT -26.005 106.595 -25.675 106.925 ;
        RECT -26.005 105.235 -25.675 105.565 ;
        RECT -26.005 103.875 -25.675 104.205 ;
        RECT -26.005 102.515 -25.675 102.845 ;
        RECT -26.005 101.155 -25.675 101.485 ;
        RECT -26.005 99.795 -25.675 100.125 ;
        RECT -26.005 98.435 -25.675 98.765 ;
        RECT -26.005 97.075 -25.675 97.405 ;
        RECT -26.005 95.715 -25.675 96.045 ;
        RECT -26.005 94.355 -25.675 94.685 ;
        RECT -26.005 92.995 -25.675 93.325 ;
        RECT -26.005 91.635 -25.675 91.965 ;
        RECT -26.005 90.275 -25.675 90.605 ;
        RECT -26.005 88.915 -25.675 89.245 ;
        RECT -26.005 87.555 -25.675 87.885 ;
        RECT -26.005 86.195 -25.675 86.525 ;
        RECT -26.005 84.835 -25.675 85.165 ;
        RECT -26.005 83.475 -25.675 83.805 ;
        RECT -26.005 82.115 -25.675 82.445 ;
        RECT -26.005 80.755 -25.675 81.085 ;
        RECT -26.005 79.395 -25.675 79.725 ;
        RECT -26.005 78.035 -25.675 78.365 ;
        RECT -26.005 76.675 -25.675 77.005 ;
        RECT -26.005 75.315 -25.675 75.645 ;
        RECT -26.005 73.955 -25.675 74.285 ;
        RECT -26.005 72.595 -25.675 72.925 ;
        RECT -26.005 71.235 -25.675 71.565 ;
        RECT -26.005 69.875 -25.675 70.205 ;
        RECT -26.005 68.515 -25.675 68.845 ;
        RECT -26.005 67.155 -25.675 67.485 ;
        RECT -26.005 65.795 -25.675 66.125 ;
        RECT -26.005 64.435 -25.675 64.765 ;
        RECT -26.005 63.075 -25.675 63.405 ;
        RECT -26.005 61.715 -25.675 62.045 ;
        RECT -26.005 60.355 -25.675 60.685 ;
        RECT -26.005 58.995 -25.675 59.325 ;
        RECT -26.005 57.635 -25.675 57.965 ;
        RECT -26.005 56.275 -25.675 56.605 ;
        RECT -26.005 54.915 -25.675 55.245 ;
        RECT -26.005 53.555 -25.675 53.885 ;
        RECT -26.005 52.195 -25.675 52.525 ;
        RECT -26.005 50.835 -25.675 51.165 ;
        RECT -26.005 49.475 -25.675 49.805 ;
        RECT -26.005 48.115 -25.675 48.445 ;
        RECT -26.005 46.755 -25.675 47.085 ;
        RECT -26.005 45.395 -25.675 45.725 ;
        RECT -26.005 44.035 -25.675 44.365 ;
        RECT -26.005 42.675 -25.675 43.005 ;
        RECT -26.005 41.315 -25.675 41.645 ;
        RECT -26.005 39.955 -25.675 40.285 ;
        RECT -26.005 38.595 -25.675 38.925 ;
        RECT -26.005 37.235 -25.675 37.565 ;
        RECT -26.005 35.875 -25.675 36.205 ;
        RECT -26.005 34.515 -25.675 34.845 ;
        RECT -26.005 33.155 -25.675 33.485 ;
        RECT -26.005 31.795 -25.675 32.125 ;
        RECT -26.005 30.435 -25.675 30.765 ;
        RECT -26.005 29.075 -25.675 29.405 ;
        RECT -26.005 27.715 -25.675 28.045 ;
        RECT -26.005 26.355 -25.675 26.685 ;
        RECT -26.005 24.995 -25.675 25.325 ;
        RECT -26.005 23.635 -25.675 23.965 ;
        RECT -26.005 22.275 -25.675 22.605 ;
        RECT -26.005 20.915 -25.675 21.245 ;
        RECT -26.005 19.555 -25.675 19.885 ;
        RECT -26.005 18.195 -25.675 18.525 ;
        RECT -26.005 16.835 -25.675 17.165 ;
        RECT -26.005 15.475 -25.675 15.805 ;
        RECT -26.005 14.115 -25.675 14.445 ;
        RECT -26.005 12.755 -25.675 13.085 ;
        RECT -26.005 11.395 -25.675 11.725 ;
        RECT -26.005 10.035 -25.675 10.365 ;
        RECT -26.005 8.675 -25.675 9.005 ;
        RECT -26.005 7.315 -25.675 7.645 ;
        RECT -26.005 5.955 -25.675 6.285 ;
        RECT -26.005 4.595 -25.675 4.925 ;
        RECT -26.005 3.235 -25.675 3.565 ;
        RECT -26.005 1.875 -25.675 2.205 ;
        RECT -26.005 0.515 -25.675 0.845 ;
        RECT -26.005 -0.845 -25.675 -0.515 ;
        RECT -26.005 -6.94 -25.675 -6.61 ;
        RECT -26.005 -7.645 -25.675 -7.315 ;
        RECT -26.005 -9.005 -25.675 -8.675 ;
        RECT -26.005 -13.085 -25.675 -12.755 ;
        RECT -26.005 -14.13 -25.675 -13.8 ;
        RECT -26.005 -17.165 -25.675 -16.835 ;
        RECT -26.005 -21.245 -25.675 -20.915 ;
        RECT -26.005 -26.685 -25.675 -26.355 ;
        RECT -26.005 -28.12 -25.675 -27.79 ;
        RECT -26.005 -29.405 -25.675 -29.075 ;
        RECT -26.005 -35.31 -25.675 -34.98 ;
        RECT -26.005 -43.005 -25.675 -42.675 ;
        RECT -26.005 -44.365 -25.675 -44.035 ;
        RECT -26.005 -45.725 -25.675 -45.395 ;
        RECT -26.005 -47.085 -25.675 -46.755 ;
        RECT -26.005 -48.445 -25.675 -48.115 ;
        RECT -26.005 -49.805 -25.675 -49.475 ;
        RECT -26.005 -51.165 -25.675 -50.835 ;
        RECT -26.005 -52.525 -25.675 -52.195 ;
        RECT -26.005 -53.885 -25.675 -53.555 ;
        RECT -26.005 -55.245 -25.675 -54.915 ;
        RECT -26.005 -56.605 -25.675 -56.275 ;
        RECT -26.005 -57.965 -25.675 -57.635 ;
        RECT -26.005 -59.325 -25.675 -58.995 ;
        RECT -26.005 -60.685 -25.675 -60.355 ;
        RECT -26.005 -62.045 -25.675 -61.715 ;
        RECT -26.005 -63.405 -25.675 -63.075 ;
        RECT -26.005 -64.765 -25.675 -64.435 ;
        RECT -26.005 -66.125 -25.675 -65.795 ;
        RECT -26.005 -67.485 -25.675 -67.155 ;
        RECT -26.005 -68.845 -25.675 -68.515 ;
        RECT -26.005 -70.205 -25.675 -69.875 ;
        RECT -26.005 -71.565 -25.675 -71.235 ;
        RECT -26.005 -72.925 -25.675 -72.595 ;
        RECT -26.005 -74.285 -25.675 -73.955 ;
        RECT -26.005 -75.645 -25.675 -75.315 ;
        RECT -26.005 -77.005 -25.675 -76.675 ;
        RECT -26.005 -78.365 -25.675 -78.035 ;
        RECT -26.005 -79.725 -25.675 -79.395 ;
        RECT -26.005 -81.085 -25.675 -80.755 ;
        RECT -26.005 -82.445 -25.675 -82.115 ;
        RECT -26.005 -83.805 -25.675 -83.475 ;
        RECT -26.005 -85.165 -25.675 -84.835 ;
        RECT -26.005 -86.525 -25.675 -86.195 ;
        RECT -26.005 -87.885 -25.675 -87.555 ;
        RECT -26.005 -89.245 -25.675 -88.915 ;
        RECT -26.005 -90.605 -25.675 -90.275 ;
        RECT -26.005 -91.965 -25.675 -91.635 ;
        RECT -26.005 -93.325 -25.675 -92.995 ;
        RECT -26.005 -94.685 -25.675 -94.355 ;
        RECT -26.005 -96.045 -25.675 -95.715 ;
        RECT -26.005 -97.405 -25.675 -97.075 ;
        RECT -26.005 -98.765 -25.675 -98.435 ;
        RECT -26.005 -100.125 -25.675 -99.795 ;
        RECT -26.005 -101.485 -25.675 -101.155 ;
        RECT -26.005 -102.845 -25.675 -102.515 ;
        RECT -26.005 -104.205 -25.675 -103.875 ;
        RECT -26.005 -109.645 -25.675 -109.315 ;
        RECT -26.005 -111.005 -25.675 -110.675 ;
        RECT -26.005 -112.365 -25.675 -112.035 ;
        RECT -26.005 -113.725 -25.675 -113.395 ;
        RECT -26.005 -115.085 -25.675 -114.755 ;
        RECT -26.005 -116.445 -25.675 -116.115 ;
        RECT -26.005 -117.805 -25.675 -117.475 ;
        RECT -26.005 -119.165 -25.675 -118.835 ;
        RECT -26.005 -120.525 -25.675 -120.195 ;
        RECT -26.005 -121.885 -25.675 -121.555 ;
        RECT -26.005 -123.245 -25.675 -122.915 ;
        RECT -26.005 -124.605 -25.675 -124.275 ;
        RECT -26.005 -125.965 -25.675 -125.635 ;
        RECT -26.005 -127.325 -25.675 -126.995 ;
        RECT -26.005 -128.685 -25.675 -128.355 ;
        RECT -26.005 -130.045 -25.675 -129.715 ;
        RECT -26.005 -131.405 -25.675 -131.075 ;
        RECT -26.005 -132.765 -25.675 -132.435 ;
        RECT -26.005 -134.125 -25.675 -133.795 ;
        RECT -26.005 -135.485 -25.675 -135.155 ;
        RECT -26.005 -136.845 -25.675 -136.515 ;
        RECT -26.005 -138.205 -25.675 -137.875 ;
        RECT -26.005 -139.565 -25.675 -139.235 ;
        RECT -26.005 -142.285 -25.675 -141.955 ;
        RECT -26.005 -143.645 -25.675 -143.315 ;
        RECT -26.005 -145.005 -25.675 -144.675 ;
        RECT -26.005 -146.365 -25.675 -146.035 ;
        RECT -26.005 -147.725 -25.675 -147.395 ;
        RECT -26.005 -149.085 -25.675 -148.755 ;
        RECT -26.005 -150.445 -25.675 -150.115 ;
        RECT -26.005 -151.805 -25.675 -151.475 ;
        RECT -26.005 -153.165 -25.675 -152.835 ;
        RECT -26.005 -154.525 -25.675 -154.195 ;
        RECT -26.005 -155.885 -25.675 -155.555 ;
        RECT -26.005 -157.245 -25.675 -156.915 ;
        RECT -26.005 -158.605 -25.675 -158.275 ;
        RECT -26.005 -159.965 -25.675 -159.635 ;
        RECT -26.005 -161.325 -25.675 -160.995 ;
        RECT -26.005 -162.685 -25.675 -162.355 ;
        RECT -26.005 -165.405 -25.675 -165.075 ;
        RECT -26.005 -166.765 -25.675 -166.435 ;
        RECT -26.005 -172.205 -25.675 -171.875 ;
        RECT -26.005 -173.565 -25.675 -173.235 ;
        RECT -26.005 -174.925 -25.675 -174.595 ;
        RECT -26.005 -176.285 -25.675 -175.955 ;
        RECT -26.005 -179.005 -25.675 -178.675 ;
        RECT -26.005 -180.365 -25.675 -180.035 ;
        RECT -26.005 -181.725 -25.675 -181.395 ;
        RECT -26.005 -184.445 -25.675 -184.115 ;
        RECT -26.005 -185.805 -25.675 -185.475 ;
        RECT -26.005 -189.885 -25.675 -189.555 ;
        RECT -26.005 -195.325 -25.675 -194.995 ;
        RECT -26.005 -196.685 -25.675 -196.355 ;
        RECT -26.005 -198.045 -25.675 -197.715 ;
        RECT -26.005 -199.405 -25.675 -199.075 ;
        RECT -26.005 -200.765 -25.675 -200.435 ;
        RECT -26.005 -202.125 -25.675 -201.795 ;
        RECT -26.005 -203.485 -25.675 -203.155 ;
        RECT -26.005 -204.845 -25.675 -204.515 ;
        RECT -26.005 -206.555 -25.675 -206.225 ;
        RECT -26.005 -207.565 -25.675 -207.235 ;
        RECT -26.005 -208.925 -25.675 -208.595 ;
        RECT -26.005 -211.645 -25.675 -211.315 ;
        RECT -26.005 -214.365 -25.675 -214.035 ;
        RECT -26.005 -215.725 -25.675 -215.395 ;
        RECT -26.005 -217.085 -25.675 -216.755 ;
        RECT -26.005 -218.445 -25.675 -218.115 ;
        RECT -26.005 -224.09 -25.675 -222.96 ;
        RECT -26 -224.205 -25.68 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -24.645 -68.845 -24.315 -68.515 ;
        RECT -24.645 -70.205 -24.315 -69.875 ;
        RECT -24.645 -71.565 -24.315 -71.235 ;
        RECT -24.645 -72.925 -24.315 -72.595 ;
        RECT -24.645 -74.285 -24.315 -73.955 ;
        RECT -24.645 -75.645 -24.315 -75.315 ;
        RECT -24.645 -77.005 -24.315 -76.675 ;
        RECT -24.645 -78.365 -24.315 -78.035 ;
        RECT -24.645 -79.725 -24.315 -79.395 ;
        RECT -24.645 -81.085 -24.315 -80.755 ;
        RECT -24.645 -82.445 -24.315 -82.115 ;
        RECT -24.645 -83.805 -24.315 -83.475 ;
        RECT -24.645 -85.165 -24.315 -84.835 ;
        RECT -24.645 -86.525 -24.315 -86.195 ;
        RECT -24.645 -87.885 -24.315 -87.555 ;
        RECT -24.645 -89.245 -24.315 -88.915 ;
        RECT -24.645 -90.605 -24.315 -90.275 ;
        RECT -24.645 -91.965 -24.315 -91.635 ;
        RECT -24.645 -93.325 -24.315 -92.995 ;
        RECT -24.645 -94.685 -24.315 -94.355 ;
        RECT -24.645 -96.045 -24.315 -95.715 ;
        RECT -24.645 -97.405 -24.315 -97.075 ;
        RECT -24.645 -98.765 -24.315 -98.435 ;
        RECT -24.645 -100.125 -24.315 -99.795 ;
        RECT -24.645 -101.485 -24.315 -101.155 ;
        RECT -24.645 -102.845 -24.315 -102.515 ;
        RECT -24.645 -104.205 -24.315 -103.875 ;
        RECT -24.645 -109.645 -24.315 -109.315 ;
        RECT -24.645 -111.005 -24.315 -110.675 ;
        RECT -24.645 -112.365 -24.315 -112.035 ;
        RECT -24.645 -113.725 -24.315 -113.395 ;
        RECT -24.645 -115.085 -24.315 -114.755 ;
        RECT -24.645 -116.445 -24.315 -116.115 ;
        RECT -24.645 -117.805 -24.315 -117.475 ;
        RECT -24.645 -119.165 -24.315 -118.835 ;
        RECT -24.645 -120.525 -24.315 -120.195 ;
        RECT -24.645 -121.885 -24.315 -121.555 ;
        RECT -24.645 -123.245 -24.315 -122.915 ;
        RECT -24.645 -124.605 -24.315 -124.275 ;
        RECT -24.645 -125.965 -24.315 -125.635 ;
        RECT -24.645 -127.325 -24.315 -126.995 ;
        RECT -24.645 -128.685 -24.315 -128.355 ;
        RECT -24.645 -130.045 -24.315 -129.715 ;
        RECT -24.645 -131.405 -24.315 -131.075 ;
        RECT -24.645 -132.765 -24.315 -132.435 ;
        RECT -24.645 -134.125 -24.315 -133.795 ;
        RECT -24.645 -135.485 -24.315 -135.155 ;
        RECT -24.645 -136.845 -24.315 -136.515 ;
        RECT -24.645 -138.205 -24.315 -137.875 ;
        RECT -24.645 -139.565 -24.315 -139.235 ;
        RECT -24.645 -142.285 -24.315 -141.955 ;
        RECT -24.645 -143.645 -24.315 -143.315 ;
        RECT -24.645 -145.005 -24.315 -144.675 ;
        RECT -24.645 -146.365 -24.315 -146.035 ;
        RECT -24.645 -147.725 -24.315 -147.395 ;
        RECT -24.645 -149.085 -24.315 -148.755 ;
        RECT -24.645 -150.445 -24.315 -150.115 ;
        RECT -24.645 -151.805 -24.315 -151.475 ;
        RECT -24.645 -153.165 -24.315 -152.835 ;
        RECT -24.645 -154.525 -24.315 -154.195 ;
        RECT -24.645 -155.885 -24.315 -155.555 ;
        RECT -24.645 -157.245 -24.315 -156.915 ;
        RECT -24.645 -158.605 -24.315 -158.275 ;
        RECT -24.645 -159.965 -24.315 -159.635 ;
        RECT -24.645 -161.325 -24.315 -160.995 ;
        RECT -24.645 -162.685 -24.315 -162.355 ;
        RECT -24.645 -165.405 -24.315 -165.075 ;
        RECT -24.645 -166.765 -24.315 -166.435 ;
        RECT -24.645 -172.205 -24.315 -171.875 ;
        RECT -24.645 -173.565 -24.315 -173.235 ;
        RECT -24.645 -174.925 -24.315 -174.595 ;
        RECT -24.645 -176.285 -24.315 -175.955 ;
        RECT -24.645 -179.005 -24.315 -178.675 ;
        RECT -24.645 -180.365 -24.315 -180.035 ;
        RECT -24.645 -181.725 -24.315 -181.395 ;
        RECT -24.645 -184.445 -24.315 -184.115 ;
        RECT -24.645 -185.805 -24.315 -185.475 ;
        RECT -24.645 -189.885 -24.315 -189.555 ;
        RECT -24.645 -195.325 -24.315 -194.995 ;
        RECT -24.645 -196.685 -24.315 -196.355 ;
        RECT -24.645 -198.045 -24.315 -197.715 ;
        RECT -24.645 -199.405 -24.315 -199.075 ;
        RECT -24.645 -200.765 -24.315 -200.435 ;
        RECT -24.645 -202.125 -24.315 -201.795 ;
        RECT -24.645 -203.485 -24.315 -203.155 ;
        RECT -24.645 -204.845 -24.315 -204.515 ;
        RECT -24.645 -206.555 -24.315 -206.225 ;
        RECT -24.645 -207.565 -24.315 -207.235 ;
        RECT -24.645 -208.925 -24.315 -208.595 ;
        RECT -24.645 -210.285 -24.315 -209.955 ;
        RECT -24.645 -211.645 -24.315 -211.315 ;
        RECT -24.645 -214.365 -24.315 -214.035 ;
        RECT -24.645 -215.725 -24.315 -215.395 ;
        RECT -24.645 -217.085 -24.315 -216.755 ;
        RECT -24.645 -218.445 -24.315 -218.115 ;
        RECT -24.645 -224.09 -24.315 -222.96 ;
        RECT -24.64 -224.205 -24.32 133.765 ;
        RECT -24.645 132.52 -24.315 133.65 ;
        RECT -24.645 128.355 -24.315 128.685 ;
        RECT -24.645 126.995 -24.315 127.325 ;
        RECT -24.645 125.635 -24.315 125.965 ;
        RECT -24.645 124.275 -24.315 124.605 ;
        RECT -24.645 122.915 -24.315 123.245 ;
        RECT -24.645 121.555 -24.315 121.885 ;
        RECT -24.645 120.195 -24.315 120.525 ;
        RECT -24.645 118.835 -24.315 119.165 ;
        RECT -24.645 117.475 -24.315 117.805 ;
        RECT -24.645 116.115 -24.315 116.445 ;
        RECT -24.645 114.755 -24.315 115.085 ;
        RECT -24.645 113.395 -24.315 113.725 ;
        RECT -24.645 112.035 -24.315 112.365 ;
        RECT -24.645 110.675 -24.315 111.005 ;
        RECT -24.645 109.315 -24.315 109.645 ;
        RECT -24.645 107.955 -24.315 108.285 ;
        RECT -24.645 106.595 -24.315 106.925 ;
        RECT -24.645 105.235 -24.315 105.565 ;
        RECT -24.645 103.875 -24.315 104.205 ;
        RECT -24.645 102.515 -24.315 102.845 ;
        RECT -24.645 101.155 -24.315 101.485 ;
        RECT -24.645 99.795 -24.315 100.125 ;
        RECT -24.645 98.435 -24.315 98.765 ;
        RECT -24.645 97.075 -24.315 97.405 ;
        RECT -24.645 95.715 -24.315 96.045 ;
        RECT -24.645 94.355 -24.315 94.685 ;
        RECT -24.645 92.995 -24.315 93.325 ;
        RECT -24.645 91.635 -24.315 91.965 ;
        RECT -24.645 90.275 -24.315 90.605 ;
        RECT -24.645 88.915 -24.315 89.245 ;
        RECT -24.645 87.555 -24.315 87.885 ;
        RECT -24.645 86.195 -24.315 86.525 ;
        RECT -24.645 84.835 -24.315 85.165 ;
        RECT -24.645 83.475 -24.315 83.805 ;
        RECT -24.645 82.115 -24.315 82.445 ;
        RECT -24.645 80.755 -24.315 81.085 ;
        RECT -24.645 79.395 -24.315 79.725 ;
        RECT -24.645 78.035 -24.315 78.365 ;
        RECT -24.645 76.675 -24.315 77.005 ;
        RECT -24.645 75.315 -24.315 75.645 ;
        RECT -24.645 73.955 -24.315 74.285 ;
        RECT -24.645 72.595 -24.315 72.925 ;
        RECT -24.645 71.235 -24.315 71.565 ;
        RECT -24.645 69.875 -24.315 70.205 ;
        RECT -24.645 68.515 -24.315 68.845 ;
        RECT -24.645 67.155 -24.315 67.485 ;
        RECT -24.645 65.795 -24.315 66.125 ;
        RECT -24.645 64.435 -24.315 64.765 ;
        RECT -24.645 63.075 -24.315 63.405 ;
        RECT -24.645 61.715 -24.315 62.045 ;
        RECT -24.645 60.355 -24.315 60.685 ;
        RECT -24.645 58.995 -24.315 59.325 ;
        RECT -24.645 57.635 -24.315 57.965 ;
        RECT -24.645 56.275 -24.315 56.605 ;
        RECT -24.645 54.915 -24.315 55.245 ;
        RECT -24.645 53.555 -24.315 53.885 ;
        RECT -24.645 52.195 -24.315 52.525 ;
        RECT -24.645 50.835 -24.315 51.165 ;
        RECT -24.645 49.475 -24.315 49.805 ;
        RECT -24.645 48.115 -24.315 48.445 ;
        RECT -24.645 46.755 -24.315 47.085 ;
        RECT -24.645 45.395 -24.315 45.725 ;
        RECT -24.645 44.035 -24.315 44.365 ;
        RECT -24.645 42.675 -24.315 43.005 ;
        RECT -24.645 41.315 -24.315 41.645 ;
        RECT -24.645 39.955 -24.315 40.285 ;
        RECT -24.645 38.595 -24.315 38.925 ;
        RECT -24.645 37.235 -24.315 37.565 ;
        RECT -24.645 35.875 -24.315 36.205 ;
        RECT -24.645 34.515 -24.315 34.845 ;
        RECT -24.645 33.155 -24.315 33.485 ;
        RECT -24.645 31.795 -24.315 32.125 ;
        RECT -24.645 30.435 -24.315 30.765 ;
        RECT -24.645 29.075 -24.315 29.405 ;
        RECT -24.645 27.715 -24.315 28.045 ;
        RECT -24.645 26.355 -24.315 26.685 ;
        RECT -24.645 24.995 -24.315 25.325 ;
        RECT -24.645 23.635 -24.315 23.965 ;
        RECT -24.645 22.275 -24.315 22.605 ;
        RECT -24.645 20.915 -24.315 21.245 ;
        RECT -24.645 19.555 -24.315 19.885 ;
        RECT -24.645 18.195 -24.315 18.525 ;
        RECT -24.645 16.835 -24.315 17.165 ;
        RECT -24.645 15.475 -24.315 15.805 ;
        RECT -24.645 14.115 -24.315 14.445 ;
        RECT -24.645 12.755 -24.315 13.085 ;
        RECT -24.645 11.395 -24.315 11.725 ;
        RECT -24.645 10.035 -24.315 10.365 ;
        RECT -24.645 8.675 -24.315 9.005 ;
        RECT -24.645 7.315 -24.315 7.645 ;
        RECT -24.645 5.955 -24.315 6.285 ;
        RECT -24.645 4.595 -24.315 4.925 ;
        RECT -24.645 3.235 -24.315 3.565 ;
        RECT -24.645 1.875 -24.315 2.205 ;
        RECT -24.645 0.515 -24.315 0.845 ;
        RECT -24.645 -0.845 -24.315 -0.515 ;
        RECT -24.645 -6.94 -24.315 -6.61 ;
        RECT -24.645 -7.645 -24.315 -7.315 ;
        RECT -24.645 -9.005 -24.315 -8.675 ;
        RECT -24.645 -13.085 -24.315 -12.755 ;
        RECT -24.645 -14.13 -24.315 -13.8 ;
        RECT -24.645 -17.165 -24.315 -16.835 ;
        RECT -24.645 -21.245 -24.315 -20.915 ;
        RECT -24.645 -26.685 -24.315 -26.355 ;
        RECT -24.645 -28.12 -24.315 -27.79 ;
        RECT -24.645 -29.405 -24.315 -29.075 ;
        RECT -24.645 -35.31 -24.315 -34.98 ;
        RECT -24.645 -43.005 -24.315 -42.675 ;
        RECT -24.645 -44.365 -24.315 -44.035 ;
        RECT -24.645 -45.725 -24.315 -45.395 ;
        RECT -24.645 -47.085 -24.315 -46.755 ;
        RECT -24.645 -48.445 -24.315 -48.115 ;
        RECT -24.645 -49.805 -24.315 -49.475 ;
        RECT -24.645 -51.165 -24.315 -50.835 ;
        RECT -24.645 -52.525 -24.315 -52.195 ;
        RECT -24.645 -53.885 -24.315 -53.555 ;
        RECT -24.645 -55.245 -24.315 -54.915 ;
        RECT -24.645 -56.605 -24.315 -56.275 ;
        RECT -24.645 -57.965 -24.315 -57.635 ;
        RECT -24.645 -59.325 -24.315 -58.995 ;
        RECT -24.645 -60.685 -24.315 -60.355 ;
        RECT -24.645 -62.045 -24.315 -61.715 ;
        RECT -24.645 -63.405 -24.315 -63.075 ;
        RECT -24.645 -64.765 -24.315 -64.435 ;
        RECT -24.645 -66.125 -24.315 -65.795 ;
        RECT -24.645 -67.485 -24.315 -67.155 ;
    END
    PORT
      LAYER met3 ;
        RECT -35.525 132.52 -35.195 133.65 ;
        RECT -35.525 128.355 -35.195 128.685 ;
        RECT -35.525 126.995 -35.195 127.325 ;
        RECT -35.525 125.635 -35.195 125.965 ;
        RECT -35.525 124.275 -35.195 124.605 ;
        RECT -35.525 122.915 -35.195 123.245 ;
        RECT -35.525 121.555 -35.195 121.885 ;
        RECT -35.525 120.195 -35.195 120.525 ;
        RECT -35.525 118.835 -35.195 119.165 ;
        RECT -35.525 117.475 -35.195 117.805 ;
        RECT -35.525 116.115 -35.195 116.445 ;
        RECT -35.525 114.755 -35.195 115.085 ;
        RECT -35.525 113.395 -35.195 113.725 ;
        RECT -35.525 112.035 -35.195 112.365 ;
        RECT -35.525 110.675 -35.195 111.005 ;
        RECT -35.525 109.315 -35.195 109.645 ;
        RECT -35.525 107.955 -35.195 108.285 ;
        RECT -35.525 106.595 -35.195 106.925 ;
        RECT -35.525 105.235 -35.195 105.565 ;
        RECT -35.525 103.875 -35.195 104.205 ;
        RECT -35.525 102.515 -35.195 102.845 ;
        RECT -35.525 101.155 -35.195 101.485 ;
        RECT -35.525 99.795 -35.195 100.125 ;
        RECT -35.525 98.435 -35.195 98.765 ;
        RECT -35.525 97.075 -35.195 97.405 ;
        RECT -35.525 95.715 -35.195 96.045 ;
        RECT -35.525 94.355 -35.195 94.685 ;
        RECT -35.525 92.995 -35.195 93.325 ;
        RECT -35.525 91.635 -35.195 91.965 ;
        RECT -35.525 90.275 -35.195 90.605 ;
        RECT -35.525 88.915 -35.195 89.245 ;
        RECT -35.525 87.555 -35.195 87.885 ;
        RECT -35.525 86.195 -35.195 86.525 ;
        RECT -35.525 84.835 -35.195 85.165 ;
        RECT -35.525 83.475 -35.195 83.805 ;
        RECT -35.525 82.115 -35.195 82.445 ;
        RECT -35.525 80.755 -35.195 81.085 ;
        RECT -35.525 79.395 -35.195 79.725 ;
        RECT -35.525 78.035 -35.195 78.365 ;
        RECT -35.525 76.675 -35.195 77.005 ;
        RECT -35.525 75.315 -35.195 75.645 ;
        RECT -35.525 73.955 -35.195 74.285 ;
        RECT -35.525 72.595 -35.195 72.925 ;
        RECT -35.525 71.235 -35.195 71.565 ;
        RECT -35.525 69.875 -35.195 70.205 ;
        RECT -35.525 68.515 -35.195 68.845 ;
        RECT -35.525 67.155 -35.195 67.485 ;
        RECT -35.525 65.795 -35.195 66.125 ;
        RECT -35.525 64.435 -35.195 64.765 ;
        RECT -35.525 63.075 -35.195 63.405 ;
        RECT -35.525 61.715 -35.195 62.045 ;
        RECT -35.525 60.355 -35.195 60.685 ;
        RECT -35.525 58.995 -35.195 59.325 ;
        RECT -35.525 57.635 -35.195 57.965 ;
        RECT -35.525 56.275 -35.195 56.605 ;
        RECT -35.525 54.915 -35.195 55.245 ;
        RECT -35.525 53.555 -35.195 53.885 ;
        RECT -35.525 52.195 -35.195 52.525 ;
        RECT -35.525 50.835 -35.195 51.165 ;
        RECT -35.525 49.475 -35.195 49.805 ;
        RECT -35.525 48.115 -35.195 48.445 ;
        RECT -35.525 46.755 -35.195 47.085 ;
        RECT -35.525 45.395 -35.195 45.725 ;
        RECT -35.525 44.035 -35.195 44.365 ;
        RECT -35.525 42.675 -35.195 43.005 ;
        RECT -35.525 41.315 -35.195 41.645 ;
        RECT -35.525 39.955 -35.195 40.285 ;
        RECT -35.525 38.595 -35.195 38.925 ;
        RECT -35.525 37.235 -35.195 37.565 ;
        RECT -35.525 35.875 -35.195 36.205 ;
        RECT -35.525 34.515 -35.195 34.845 ;
        RECT -35.525 33.155 -35.195 33.485 ;
        RECT -35.525 31.795 -35.195 32.125 ;
        RECT -35.525 30.435 -35.195 30.765 ;
        RECT -35.525 29.075 -35.195 29.405 ;
        RECT -35.525 27.715 -35.195 28.045 ;
        RECT -35.525 26.355 -35.195 26.685 ;
        RECT -35.525 24.995 -35.195 25.325 ;
        RECT -35.525 23.635 -35.195 23.965 ;
        RECT -35.525 22.275 -35.195 22.605 ;
        RECT -35.525 20.915 -35.195 21.245 ;
        RECT -35.525 19.555 -35.195 19.885 ;
        RECT -35.525 18.195 -35.195 18.525 ;
        RECT -35.525 16.835 -35.195 17.165 ;
        RECT -35.525 15.475 -35.195 15.805 ;
        RECT -35.525 14.115 -35.195 14.445 ;
        RECT -35.525 12.755 -35.195 13.085 ;
        RECT -35.525 11.395 -35.195 11.725 ;
        RECT -35.525 10.035 -35.195 10.365 ;
        RECT -35.525 8.675 -35.195 9.005 ;
        RECT -35.525 7.315 -35.195 7.645 ;
        RECT -35.525 5.955 -35.195 6.285 ;
        RECT -35.525 4.595 -35.195 4.925 ;
        RECT -35.525 3.235 -35.195 3.565 ;
        RECT -35.525 1.875 -35.195 2.205 ;
        RECT -35.525 0.515 -35.195 0.845 ;
        RECT -35.525 -0.845 -35.195 -0.515 ;
        RECT -35.525 -2.205 -35.195 -1.875 ;
        RECT -35.525 -6.285 -35.195 -5.955 ;
        RECT -35.525 -7.645 -35.195 -7.315 ;
        RECT -35.525 -9.005 -35.195 -8.675 ;
        RECT -35.525 -11.725 -35.195 -11.395 ;
        RECT -35.525 -13.085 -35.195 -12.755 ;
        RECT -35.525 -14.445 -35.195 -14.115 ;
        RECT -35.525 -15.805 -35.195 -15.475 ;
        RECT -35.525 -17.165 -35.195 -16.835 ;
        RECT -35.525 -18.525 -35.195 -18.195 ;
        RECT -35.525 -19.885 -35.195 -19.555 ;
        RECT -35.525 -26.685 -35.195 -26.355 ;
        RECT -35.525 -28.045 -35.195 -27.715 ;
        RECT -35.525 -29.405 -35.195 -29.075 ;
        RECT -35.525 -32.125 -35.195 -31.795 ;
        RECT -35.525 -34.845 -35.195 -34.515 ;
        RECT -35.525 -37.565 -35.195 -37.235 ;
        RECT -35.525 -38.925 -35.195 -38.595 ;
        RECT -35.525 -40.285 -35.195 -39.955 ;
        RECT -35.525 -41.645 -35.195 -41.315 ;
        RECT -35.525 -43.005 -35.195 -42.675 ;
        RECT -35.525 -44.365 -35.195 -44.035 ;
        RECT -35.525 -45.725 -35.195 -45.395 ;
        RECT -35.525 -47.085 -35.195 -46.755 ;
        RECT -35.525 -48.445 -35.195 -48.115 ;
        RECT -35.525 -49.805 -35.195 -49.475 ;
        RECT -35.525 -51.165 -35.195 -50.835 ;
        RECT -35.525 -52.525 -35.195 -52.195 ;
        RECT -35.525 -53.885 -35.195 -53.555 ;
        RECT -35.525 -55.245 -35.195 -54.915 ;
        RECT -35.525 -56.605 -35.195 -56.275 ;
        RECT -35.525 -57.965 -35.195 -57.635 ;
        RECT -35.525 -59.325 -35.195 -58.995 ;
        RECT -35.525 -60.685 -35.195 -60.355 ;
        RECT -35.525 -62.045 -35.195 -61.715 ;
        RECT -35.525 -63.405 -35.195 -63.075 ;
        RECT -35.525 -64.765 -35.195 -64.435 ;
        RECT -35.525 -66.125 -35.195 -65.795 ;
        RECT -35.525 -67.485 -35.195 -67.155 ;
        RECT -35.525 -68.845 -35.195 -68.515 ;
        RECT -35.525 -70.205 -35.195 -69.875 ;
        RECT -35.525 -71.565 -35.195 -71.235 ;
        RECT -35.525 -72.925 -35.195 -72.595 ;
        RECT -35.525 -74.285 -35.195 -73.955 ;
        RECT -35.525 -75.645 -35.195 -75.315 ;
        RECT -35.525 -77.005 -35.195 -76.675 ;
        RECT -35.525 -78.365 -35.195 -78.035 ;
        RECT -35.525 -79.725 -35.195 -79.395 ;
        RECT -35.525 -81.085 -35.195 -80.755 ;
        RECT -35.525 -82.445 -35.195 -82.115 ;
        RECT -35.525 -83.805 -35.195 -83.475 ;
        RECT -35.525 -85.165 -35.195 -84.835 ;
        RECT -35.525 -86.525 -35.195 -86.195 ;
        RECT -35.525 -87.885 -35.195 -87.555 ;
        RECT -35.525 -89.245 -35.195 -88.915 ;
        RECT -35.525 -90.605 -35.195 -90.275 ;
        RECT -35.525 -91.965 -35.195 -91.635 ;
        RECT -35.525 -93.325 -35.195 -92.995 ;
        RECT -35.525 -94.685 -35.195 -94.355 ;
        RECT -35.525 -96.045 -35.195 -95.715 ;
        RECT -35.525 -97.405 -35.195 -97.075 ;
        RECT -35.525 -98.765 -35.195 -98.435 ;
        RECT -35.525 -100.125 -35.195 -99.795 ;
        RECT -35.525 -101.485 -35.195 -101.155 ;
        RECT -35.525 -102.845 -35.195 -102.515 ;
        RECT -35.525 -104.205 -35.195 -103.875 ;
        RECT -35.525 -105.565 -35.195 -105.235 ;
        RECT -35.525 -106.925 -35.195 -106.595 ;
        RECT -35.525 -109.645 -35.195 -109.315 ;
        RECT -35.525 -111.005 -35.195 -110.675 ;
        RECT -35.525 -111.87 -35.195 -111.54 ;
        RECT -35.525 -113.725 -35.195 -113.395 ;
        RECT -35.525 -115.085 -35.195 -114.755 ;
        RECT -35.525 -116.445 -35.195 -116.115 ;
        RECT -35.525 -117.805 -35.195 -117.475 ;
        RECT -35.525 -120.525 -35.195 -120.195 ;
        RECT -35.525 -121.885 -35.195 -121.555 ;
        RECT -35.525 -123.245 -35.195 -122.915 ;
        RECT -35.525 -124.71 -35.195 -124.38 ;
        RECT -35.525 -125.965 -35.195 -125.635 ;
        RECT -35.525 -127.325 -35.195 -126.995 ;
        RECT -35.525 -130.045 -35.195 -129.715 ;
        RECT -35.52 -132.08 -35.2 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -35.525 -214.365 -35.195 -214.035 ;
        RECT -35.525 -215.725 -35.195 -215.395 ;
        RECT -35.525 -217.085 -35.195 -216.755 ;
        RECT -35.525 -218.445 -35.195 -218.115 ;
        RECT -35.525 -224.09 -35.195 -222.96 ;
        RECT -35.52 -224.205 -35.2 -210.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -34.165 132.52 -33.835 133.65 ;
        RECT -34.165 128.355 -33.835 128.685 ;
        RECT -34.165 126.995 -33.835 127.325 ;
        RECT -34.165 125.635 -33.835 125.965 ;
        RECT -34.165 124.275 -33.835 124.605 ;
        RECT -34.165 122.915 -33.835 123.245 ;
        RECT -34.165 121.555 -33.835 121.885 ;
        RECT -34.165 120.195 -33.835 120.525 ;
        RECT -34.165 118.835 -33.835 119.165 ;
        RECT -34.165 117.475 -33.835 117.805 ;
        RECT -34.165 116.115 -33.835 116.445 ;
        RECT -34.165 114.755 -33.835 115.085 ;
        RECT -34.165 113.395 -33.835 113.725 ;
        RECT -34.165 112.035 -33.835 112.365 ;
        RECT -34.165 110.675 -33.835 111.005 ;
        RECT -34.165 109.315 -33.835 109.645 ;
        RECT -34.165 107.955 -33.835 108.285 ;
        RECT -34.165 106.595 -33.835 106.925 ;
        RECT -34.165 105.235 -33.835 105.565 ;
        RECT -34.165 103.875 -33.835 104.205 ;
        RECT -34.165 102.515 -33.835 102.845 ;
        RECT -34.165 101.155 -33.835 101.485 ;
        RECT -34.165 99.795 -33.835 100.125 ;
        RECT -34.165 98.435 -33.835 98.765 ;
        RECT -34.165 97.075 -33.835 97.405 ;
        RECT -34.165 95.715 -33.835 96.045 ;
        RECT -34.165 94.355 -33.835 94.685 ;
        RECT -34.165 92.995 -33.835 93.325 ;
        RECT -34.165 91.635 -33.835 91.965 ;
        RECT -34.165 90.275 -33.835 90.605 ;
        RECT -34.165 88.915 -33.835 89.245 ;
        RECT -34.165 87.555 -33.835 87.885 ;
        RECT -34.165 86.195 -33.835 86.525 ;
        RECT -34.165 84.835 -33.835 85.165 ;
        RECT -34.165 83.475 -33.835 83.805 ;
        RECT -34.165 82.115 -33.835 82.445 ;
        RECT -34.165 80.755 -33.835 81.085 ;
        RECT -34.165 79.395 -33.835 79.725 ;
        RECT -34.165 78.035 -33.835 78.365 ;
        RECT -34.165 76.675 -33.835 77.005 ;
        RECT -34.165 75.315 -33.835 75.645 ;
        RECT -34.165 73.955 -33.835 74.285 ;
        RECT -34.165 72.595 -33.835 72.925 ;
        RECT -34.165 71.235 -33.835 71.565 ;
        RECT -34.165 69.875 -33.835 70.205 ;
        RECT -34.165 68.515 -33.835 68.845 ;
        RECT -34.165 67.155 -33.835 67.485 ;
        RECT -34.165 65.795 -33.835 66.125 ;
        RECT -34.165 64.435 -33.835 64.765 ;
        RECT -34.165 63.075 -33.835 63.405 ;
        RECT -34.165 61.715 -33.835 62.045 ;
        RECT -34.165 60.355 -33.835 60.685 ;
        RECT -34.165 58.995 -33.835 59.325 ;
        RECT -34.165 57.635 -33.835 57.965 ;
        RECT -34.165 56.275 -33.835 56.605 ;
        RECT -34.165 54.915 -33.835 55.245 ;
        RECT -34.165 53.555 -33.835 53.885 ;
        RECT -34.165 52.195 -33.835 52.525 ;
        RECT -34.165 50.835 -33.835 51.165 ;
        RECT -34.165 49.475 -33.835 49.805 ;
        RECT -34.165 48.115 -33.835 48.445 ;
        RECT -34.165 46.755 -33.835 47.085 ;
        RECT -34.165 45.395 -33.835 45.725 ;
        RECT -34.165 44.035 -33.835 44.365 ;
        RECT -34.165 42.675 -33.835 43.005 ;
        RECT -34.165 41.315 -33.835 41.645 ;
        RECT -34.165 39.955 -33.835 40.285 ;
        RECT -34.165 38.595 -33.835 38.925 ;
        RECT -34.165 37.235 -33.835 37.565 ;
        RECT -34.165 35.875 -33.835 36.205 ;
        RECT -34.165 34.515 -33.835 34.845 ;
        RECT -34.165 33.155 -33.835 33.485 ;
        RECT -34.165 31.795 -33.835 32.125 ;
        RECT -34.165 30.435 -33.835 30.765 ;
        RECT -34.165 29.075 -33.835 29.405 ;
        RECT -34.165 27.715 -33.835 28.045 ;
        RECT -34.165 26.355 -33.835 26.685 ;
        RECT -34.165 24.995 -33.835 25.325 ;
        RECT -34.165 23.635 -33.835 23.965 ;
        RECT -34.165 22.275 -33.835 22.605 ;
        RECT -34.165 20.915 -33.835 21.245 ;
        RECT -34.165 19.555 -33.835 19.885 ;
        RECT -34.165 18.195 -33.835 18.525 ;
        RECT -34.165 16.835 -33.835 17.165 ;
        RECT -34.165 15.475 -33.835 15.805 ;
        RECT -34.165 14.115 -33.835 14.445 ;
        RECT -34.165 12.755 -33.835 13.085 ;
        RECT -34.165 11.395 -33.835 11.725 ;
        RECT -34.165 10.035 -33.835 10.365 ;
        RECT -34.165 8.675 -33.835 9.005 ;
        RECT -34.165 7.315 -33.835 7.645 ;
        RECT -34.165 5.955 -33.835 6.285 ;
        RECT -34.165 4.595 -33.835 4.925 ;
        RECT -34.165 3.235 -33.835 3.565 ;
        RECT -34.165 1.875 -33.835 2.205 ;
        RECT -34.165 0.515 -33.835 0.845 ;
        RECT -34.165 -0.845 -33.835 -0.515 ;
        RECT -34.165 -6.285 -33.835 -5.955 ;
        RECT -34.165 -7.645 -33.835 -7.315 ;
        RECT -34.165 -9.005 -33.835 -8.675 ;
        RECT -34.165 -11.725 -33.835 -11.395 ;
        RECT -34.165 -13.085 -33.835 -12.755 ;
        RECT -34.165 -14.445 -33.835 -14.115 ;
        RECT -34.165 -15.805 -33.835 -15.475 ;
        RECT -34.165 -17.165 -33.835 -16.835 ;
        RECT -34.165 -18.525 -33.835 -18.195 ;
        RECT -34.165 -19.885 -33.835 -19.555 ;
        RECT -34.165 -26.685 -33.835 -26.355 ;
        RECT -34.165 -28.045 -33.835 -27.715 ;
        RECT -34.165 -29.405 -33.835 -29.075 ;
        RECT -34.165 -32.125 -33.835 -31.795 ;
        RECT -34.165 -34.845 -33.835 -34.515 ;
        RECT -34.165 -37.565 -33.835 -37.235 ;
        RECT -34.165 -38.925 -33.835 -38.595 ;
        RECT -34.165 -40.285 -33.835 -39.955 ;
        RECT -34.165 -41.645 -33.835 -41.315 ;
        RECT -34.165 -43.005 -33.835 -42.675 ;
        RECT -34.165 -44.365 -33.835 -44.035 ;
        RECT -34.165 -45.725 -33.835 -45.395 ;
        RECT -34.165 -47.085 -33.835 -46.755 ;
        RECT -34.165 -48.445 -33.835 -48.115 ;
        RECT -34.165 -49.805 -33.835 -49.475 ;
        RECT -34.165 -51.165 -33.835 -50.835 ;
        RECT -34.165 -52.525 -33.835 -52.195 ;
        RECT -34.165 -53.885 -33.835 -53.555 ;
        RECT -34.165 -55.245 -33.835 -54.915 ;
        RECT -34.165 -56.605 -33.835 -56.275 ;
        RECT -34.165 -57.965 -33.835 -57.635 ;
        RECT -34.165 -59.325 -33.835 -58.995 ;
        RECT -34.165 -60.685 -33.835 -60.355 ;
        RECT -34.165 -62.045 -33.835 -61.715 ;
        RECT -34.165 -63.405 -33.835 -63.075 ;
        RECT -34.165 -64.765 -33.835 -64.435 ;
        RECT -34.165 -66.125 -33.835 -65.795 ;
        RECT -34.165 -67.485 -33.835 -67.155 ;
        RECT -34.165 -68.845 -33.835 -68.515 ;
        RECT -34.165 -70.205 -33.835 -69.875 ;
        RECT -34.165 -71.565 -33.835 -71.235 ;
        RECT -34.165 -72.925 -33.835 -72.595 ;
        RECT -34.165 -74.285 -33.835 -73.955 ;
        RECT -34.165 -75.645 -33.835 -75.315 ;
        RECT -34.165 -77.005 -33.835 -76.675 ;
        RECT -34.165 -78.365 -33.835 -78.035 ;
        RECT -34.165 -79.725 -33.835 -79.395 ;
        RECT -34.165 -81.085 -33.835 -80.755 ;
        RECT -34.165 -82.445 -33.835 -82.115 ;
        RECT -34.165 -83.805 -33.835 -83.475 ;
        RECT -34.165 -85.165 -33.835 -84.835 ;
        RECT -34.165 -86.525 -33.835 -86.195 ;
        RECT -34.165 -87.885 -33.835 -87.555 ;
        RECT -34.165 -89.245 -33.835 -88.915 ;
        RECT -34.165 -90.605 -33.835 -90.275 ;
        RECT -34.165 -91.965 -33.835 -91.635 ;
        RECT -34.165 -93.325 -33.835 -92.995 ;
        RECT -34.165 -94.685 -33.835 -94.355 ;
        RECT -34.165 -96.045 -33.835 -95.715 ;
        RECT -34.165 -97.405 -33.835 -97.075 ;
        RECT -34.165 -98.765 -33.835 -98.435 ;
        RECT -34.165 -100.125 -33.835 -99.795 ;
        RECT -34.165 -101.485 -33.835 -101.155 ;
        RECT -34.165 -102.845 -33.835 -102.515 ;
        RECT -34.165 -104.205 -33.835 -103.875 ;
        RECT -34.165 -105.565 -33.835 -105.235 ;
        RECT -34.165 -109.645 -33.835 -109.315 ;
        RECT -34.165 -111.005 -33.835 -110.675 ;
        RECT -34.165 -111.87 -33.835 -111.54 ;
        RECT -34.165 -113.725 -33.835 -113.395 ;
        RECT -34.165 -115.085 -33.835 -114.755 ;
        RECT -34.165 -116.445 -33.835 -116.115 ;
        RECT -34.165 -117.805 -33.835 -117.475 ;
        RECT -34.165 -120.525 -33.835 -120.195 ;
        RECT -34.165 -121.885 -33.835 -121.555 ;
        RECT -34.165 -123.245 -33.835 -122.915 ;
        RECT -34.165 -124.71 -33.835 -124.38 ;
        RECT -34.165 -125.965 -33.835 -125.635 ;
        RECT -34.165 -127.325 -33.835 -126.995 ;
        RECT -34.165 -130.045 -33.835 -129.715 ;
        RECT -34.165 -132.765 -33.835 -132.435 ;
        RECT -34.165 -134.125 -33.835 -133.795 ;
        RECT -34.165 -135.485 -33.835 -135.155 ;
        RECT -34.165 -136.845 -33.835 -136.515 ;
        RECT -34.165 -138.205 -33.835 -137.875 ;
        RECT -34.165 -139.565 -33.835 -139.235 ;
        RECT -34.165 -142.285 -33.835 -141.955 ;
        RECT -34.165 -143.645 -33.835 -143.315 ;
        RECT -34.165 -145.005 -33.835 -144.675 ;
        RECT -34.165 -146.365 -33.835 -146.035 ;
        RECT -34.165 -147.725 -33.835 -147.395 ;
        RECT -34.165 -149.085 -33.835 -148.755 ;
        RECT -34.165 -150.445 -33.835 -150.115 ;
        RECT -34.165 -151.805 -33.835 -151.475 ;
        RECT -34.165 -153.165 -33.835 -152.835 ;
        RECT -34.165 -154.525 -33.835 -154.195 ;
        RECT -34.165 -155.885 -33.835 -155.555 ;
        RECT -34.165 -157.245 -33.835 -156.915 ;
        RECT -34.165 -158.605 -33.835 -158.275 ;
        RECT -34.165 -159.965 -33.835 -159.635 ;
        RECT -34.165 -161.325 -33.835 -160.995 ;
        RECT -34.165 -162.685 -33.835 -162.355 ;
        RECT -34.165 -164.045 -33.835 -163.715 ;
        RECT -34.165 -165.405 -33.835 -165.075 ;
        RECT -34.165 -166.765 -33.835 -166.435 ;
        RECT -34.165 -168.125 -33.835 -167.795 ;
        RECT -34.165 -170.845 -33.835 -170.515 ;
        RECT -34.165 -172.205 -33.835 -171.875 ;
        RECT -34.165 -173.565 -33.835 -173.235 ;
        RECT -34.165 -174.925 -33.835 -174.595 ;
        RECT -34.165 -176.285 -33.835 -175.955 ;
        RECT -34.165 -177.645 -33.835 -177.315 ;
        RECT -34.165 -179.005 -33.835 -178.675 ;
        RECT -34.165 -180.365 -33.835 -180.035 ;
        RECT -34.165 -181.725 -33.835 -181.395 ;
        RECT -34.165 -183.085 -33.835 -182.755 ;
        RECT -34.165 -184.445 -33.835 -184.115 ;
        RECT -34.165 -185.805 -33.835 -185.475 ;
        RECT -34.165 -188.525 -33.835 -188.195 ;
        RECT -34.165 -189.885 -33.835 -189.555 ;
        RECT -34.165 -192.605 -33.835 -192.275 ;
        RECT -34.165 -195.325 -33.835 -194.995 ;
        RECT -34.165 -196.685 -33.835 -196.355 ;
        RECT -34.165 -198.045 -33.835 -197.715 ;
        RECT -34.165 -199.405 -33.835 -199.075 ;
        RECT -34.165 -200.765 -33.835 -200.435 ;
        RECT -34.165 -202.125 -33.835 -201.795 ;
        RECT -34.165 -203.485 -33.835 -203.155 ;
        RECT -34.165 -204.845 -33.835 -204.515 ;
        RECT -34.165 -206.555 -33.835 -206.225 ;
        RECT -34.165 -207.565 -33.835 -207.235 ;
        RECT -34.165 -208.925 -33.835 -208.595 ;
        RECT -34.16 -209.6 -33.84 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -32.805 132.52 -32.475 133.65 ;
        RECT -32.805 128.355 -32.475 128.685 ;
        RECT -32.805 126.995 -32.475 127.325 ;
        RECT -32.805 125.635 -32.475 125.965 ;
        RECT -32.805 124.275 -32.475 124.605 ;
        RECT -32.805 122.915 -32.475 123.245 ;
        RECT -32.805 121.555 -32.475 121.885 ;
        RECT -32.805 120.195 -32.475 120.525 ;
        RECT -32.805 118.835 -32.475 119.165 ;
        RECT -32.805 117.475 -32.475 117.805 ;
        RECT -32.805 116.115 -32.475 116.445 ;
        RECT -32.805 114.755 -32.475 115.085 ;
        RECT -32.805 113.395 -32.475 113.725 ;
        RECT -32.805 112.035 -32.475 112.365 ;
        RECT -32.805 110.675 -32.475 111.005 ;
        RECT -32.805 109.315 -32.475 109.645 ;
        RECT -32.805 107.955 -32.475 108.285 ;
        RECT -32.805 106.595 -32.475 106.925 ;
        RECT -32.805 105.235 -32.475 105.565 ;
        RECT -32.805 103.875 -32.475 104.205 ;
        RECT -32.805 102.515 -32.475 102.845 ;
        RECT -32.805 101.155 -32.475 101.485 ;
        RECT -32.805 99.795 -32.475 100.125 ;
        RECT -32.805 98.435 -32.475 98.765 ;
        RECT -32.805 97.075 -32.475 97.405 ;
        RECT -32.805 95.715 -32.475 96.045 ;
        RECT -32.805 94.355 -32.475 94.685 ;
        RECT -32.805 92.995 -32.475 93.325 ;
        RECT -32.805 91.635 -32.475 91.965 ;
        RECT -32.805 90.275 -32.475 90.605 ;
        RECT -32.805 88.915 -32.475 89.245 ;
        RECT -32.805 87.555 -32.475 87.885 ;
        RECT -32.805 86.195 -32.475 86.525 ;
        RECT -32.805 84.835 -32.475 85.165 ;
        RECT -32.805 83.475 -32.475 83.805 ;
        RECT -32.805 82.115 -32.475 82.445 ;
        RECT -32.805 80.755 -32.475 81.085 ;
        RECT -32.805 79.395 -32.475 79.725 ;
        RECT -32.805 78.035 -32.475 78.365 ;
        RECT -32.805 76.675 -32.475 77.005 ;
        RECT -32.805 75.315 -32.475 75.645 ;
        RECT -32.805 73.955 -32.475 74.285 ;
        RECT -32.805 72.595 -32.475 72.925 ;
        RECT -32.805 71.235 -32.475 71.565 ;
        RECT -32.805 69.875 -32.475 70.205 ;
        RECT -32.805 68.515 -32.475 68.845 ;
        RECT -32.805 67.155 -32.475 67.485 ;
        RECT -32.805 65.795 -32.475 66.125 ;
        RECT -32.805 64.435 -32.475 64.765 ;
        RECT -32.805 63.075 -32.475 63.405 ;
        RECT -32.805 61.715 -32.475 62.045 ;
        RECT -32.805 60.355 -32.475 60.685 ;
        RECT -32.805 58.995 -32.475 59.325 ;
        RECT -32.805 57.635 -32.475 57.965 ;
        RECT -32.805 56.275 -32.475 56.605 ;
        RECT -32.805 54.915 -32.475 55.245 ;
        RECT -32.805 53.555 -32.475 53.885 ;
        RECT -32.805 52.195 -32.475 52.525 ;
        RECT -32.805 50.835 -32.475 51.165 ;
        RECT -32.805 49.475 -32.475 49.805 ;
        RECT -32.805 48.115 -32.475 48.445 ;
        RECT -32.805 46.755 -32.475 47.085 ;
        RECT -32.805 45.395 -32.475 45.725 ;
        RECT -32.805 44.035 -32.475 44.365 ;
        RECT -32.805 42.675 -32.475 43.005 ;
        RECT -32.805 41.315 -32.475 41.645 ;
        RECT -32.805 39.955 -32.475 40.285 ;
        RECT -32.805 38.595 -32.475 38.925 ;
        RECT -32.805 37.235 -32.475 37.565 ;
        RECT -32.805 35.875 -32.475 36.205 ;
        RECT -32.805 34.515 -32.475 34.845 ;
        RECT -32.805 33.155 -32.475 33.485 ;
        RECT -32.805 31.795 -32.475 32.125 ;
        RECT -32.805 30.435 -32.475 30.765 ;
        RECT -32.805 29.075 -32.475 29.405 ;
        RECT -32.805 27.715 -32.475 28.045 ;
        RECT -32.805 26.355 -32.475 26.685 ;
        RECT -32.805 24.995 -32.475 25.325 ;
        RECT -32.805 23.635 -32.475 23.965 ;
        RECT -32.805 22.275 -32.475 22.605 ;
        RECT -32.805 20.915 -32.475 21.245 ;
        RECT -32.805 19.555 -32.475 19.885 ;
        RECT -32.805 18.195 -32.475 18.525 ;
        RECT -32.805 16.835 -32.475 17.165 ;
        RECT -32.805 15.475 -32.475 15.805 ;
        RECT -32.805 14.115 -32.475 14.445 ;
        RECT -32.805 12.755 -32.475 13.085 ;
        RECT -32.805 11.395 -32.475 11.725 ;
        RECT -32.805 10.035 -32.475 10.365 ;
        RECT -32.805 8.675 -32.475 9.005 ;
        RECT -32.805 7.315 -32.475 7.645 ;
        RECT -32.805 5.955 -32.475 6.285 ;
        RECT -32.805 4.595 -32.475 4.925 ;
        RECT -32.805 3.235 -32.475 3.565 ;
        RECT -32.805 1.875 -32.475 2.205 ;
        RECT -32.805 0.515 -32.475 0.845 ;
        RECT -32.805 -6.285 -32.475 -5.955 ;
        RECT -32.805 -7.645 -32.475 -7.315 ;
        RECT -32.805 -9.005 -32.475 -8.675 ;
        RECT -32.805 -11.725 -32.475 -11.395 ;
        RECT -32.805 -13.085 -32.475 -12.755 ;
        RECT -32.805 -14.445 -32.475 -14.115 ;
        RECT -32.805 -15.805 -32.475 -15.475 ;
        RECT -32.805 -17.165 -32.475 -16.835 ;
        RECT -32.805 -18.525 -32.475 -18.195 ;
        RECT -32.805 -19.885 -32.475 -19.555 ;
        RECT -32.805 -26.685 -32.475 -26.355 ;
        RECT -32.805 -28.045 -32.475 -27.715 ;
        RECT -32.805 -29.405 -32.475 -29.075 ;
        RECT -32.805 -32.125 -32.475 -31.795 ;
        RECT -32.805 -34.845 -32.475 -34.515 ;
        RECT -32.805 -37.565 -32.475 -37.235 ;
        RECT -32.805 -38.925 -32.475 -38.595 ;
        RECT -32.805 -40.285 -32.475 -39.955 ;
        RECT -32.805 -41.645 -32.475 -41.315 ;
        RECT -32.805 -43.005 -32.475 -42.675 ;
        RECT -32.805 -44.365 -32.475 -44.035 ;
        RECT -32.805 -45.725 -32.475 -45.395 ;
        RECT -32.805 -47.085 -32.475 -46.755 ;
        RECT -32.805 -48.445 -32.475 -48.115 ;
        RECT -32.805 -49.805 -32.475 -49.475 ;
        RECT -32.805 -51.165 -32.475 -50.835 ;
        RECT -32.805 -52.525 -32.475 -52.195 ;
        RECT -32.805 -53.885 -32.475 -53.555 ;
        RECT -32.805 -55.245 -32.475 -54.915 ;
        RECT -32.805 -56.605 -32.475 -56.275 ;
        RECT -32.805 -57.965 -32.475 -57.635 ;
        RECT -32.805 -59.325 -32.475 -58.995 ;
        RECT -32.805 -60.685 -32.475 -60.355 ;
        RECT -32.805 -62.045 -32.475 -61.715 ;
        RECT -32.805 -63.405 -32.475 -63.075 ;
        RECT -32.805 -64.765 -32.475 -64.435 ;
        RECT -32.805 -66.125 -32.475 -65.795 ;
        RECT -32.805 -67.485 -32.475 -67.155 ;
        RECT -32.805 -68.845 -32.475 -68.515 ;
        RECT -32.805 -70.205 -32.475 -69.875 ;
        RECT -32.805 -71.565 -32.475 -71.235 ;
        RECT -32.805 -72.925 -32.475 -72.595 ;
        RECT -32.805 -74.285 -32.475 -73.955 ;
        RECT -32.805 -75.645 -32.475 -75.315 ;
        RECT -32.805 -77.005 -32.475 -76.675 ;
        RECT -32.805 -78.365 -32.475 -78.035 ;
        RECT -32.805 -79.725 -32.475 -79.395 ;
        RECT -32.805 -81.085 -32.475 -80.755 ;
        RECT -32.805 -82.445 -32.475 -82.115 ;
        RECT -32.805 -83.805 -32.475 -83.475 ;
        RECT -32.805 -85.165 -32.475 -84.835 ;
        RECT -32.805 -86.525 -32.475 -86.195 ;
        RECT -32.805 -87.885 -32.475 -87.555 ;
        RECT -32.805 -89.245 -32.475 -88.915 ;
        RECT -32.805 -90.605 -32.475 -90.275 ;
        RECT -32.805 -91.965 -32.475 -91.635 ;
        RECT -32.805 -93.325 -32.475 -92.995 ;
        RECT -32.805 -94.685 -32.475 -94.355 ;
        RECT -32.805 -96.045 -32.475 -95.715 ;
        RECT -32.805 -97.405 -32.475 -97.075 ;
        RECT -32.805 -98.765 -32.475 -98.435 ;
        RECT -32.805 -100.125 -32.475 -99.795 ;
        RECT -32.805 -101.485 -32.475 -101.155 ;
        RECT -32.805 -102.845 -32.475 -102.515 ;
        RECT -32.805 -104.205 -32.475 -103.875 ;
        RECT -32.805 -105.565 -32.475 -105.235 ;
        RECT -32.805 -109.645 -32.475 -109.315 ;
        RECT -32.805 -111.005 -32.475 -110.675 ;
        RECT -32.805 -111.87 -32.475 -111.54 ;
        RECT -32.805 -113.725 -32.475 -113.395 ;
        RECT -32.805 -115.085 -32.475 -114.755 ;
        RECT -32.805 -116.445 -32.475 -116.115 ;
        RECT -32.805 -117.805 -32.475 -117.475 ;
        RECT -32.805 -120.525 -32.475 -120.195 ;
        RECT -32.805 -121.885 -32.475 -121.555 ;
        RECT -32.805 -123.245 -32.475 -122.915 ;
        RECT -32.805 -124.71 -32.475 -124.38 ;
        RECT -32.805 -125.965 -32.475 -125.635 ;
        RECT -32.805 -127.325 -32.475 -126.995 ;
        RECT -32.805 -130.045 -32.475 -129.715 ;
        RECT -32.805 -132.765 -32.475 -132.435 ;
        RECT -32.805 -134.125 -32.475 -133.795 ;
        RECT -32.805 -135.485 -32.475 -135.155 ;
        RECT -32.805 -136.845 -32.475 -136.515 ;
        RECT -32.805 -138.205 -32.475 -137.875 ;
        RECT -32.805 -139.565 -32.475 -139.235 ;
        RECT -32.805 -142.285 -32.475 -141.955 ;
        RECT -32.805 -143.645 -32.475 -143.315 ;
        RECT -32.805 -145.005 -32.475 -144.675 ;
        RECT -32.805 -146.365 -32.475 -146.035 ;
        RECT -32.805 -147.725 -32.475 -147.395 ;
        RECT -32.805 -149.085 -32.475 -148.755 ;
        RECT -32.805 -150.445 -32.475 -150.115 ;
        RECT -32.805 -151.805 -32.475 -151.475 ;
        RECT -32.805 -153.165 -32.475 -152.835 ;
        RECT -32.805 -154.525 -32.475 -154.195 ;
        RECT -32.805 -155.885 -32.475 -155.555 ;
        RECT -32.805 -157.245 -32.475 -156.915 ;
        RECT -32.805 -158.605 -32.475 -158.275 ;
        RECT -32.805 -159.965 -32.475 -159.635 ;
        RECT -32.805 -161.325 -32.475 -160.995 ;
        RECT -32.805 -162.685 -32.475 -162.355 ;
        RECT -32.805 -164.045 -32.475 -163.715 ;
        RECT -32.805 -165.405 -32.475 -165.075 ;
        RECT -32.805 -166.765 -32.475 -166.435 ;
        RECT -32.805 -168.125 -32.475 -167.795 ;
        RECT -32.805 -170.845 -32.475 -170.515 ;
        RECT -32.805 -172.205 -32.475 -171.875 ;
        RECT -32.805 -173.565 -32.475 -173.235 ;
        RECT -32.805 -174.925 -32.475 -174.595 ;
        RECT -32.805 -176.285 -32.475 -175.955 ;
        RECT -32.805 -177.645 -32.475 -177.315 ;
        RECT -32.805 -179.005 -32.475 -178.675 ;
        RECT -32.805 -180.365 -32.475 -180.035 ;
        RECT -32.805 -181.725 -32.475 -181.395 ;
        RECT -32.805 -183.085 -32.475 -182.755 ;
        RECT -32.805 -184.445 -32.475 -184.115 ;
        RECT -32.805 -185.805 -32.475 -185.475 ;
        RECT -32.805 -188.525 -32.475 -188.195 ;
        RECT -32.805 -189.885 -32.475 -189.555 ;
        RECT -32.805 -192.605 -32.475 -192.275 ;
        RECT -32.805 -193.965 -32.475 -193.635 ;
        RECT -32.805 -195.325 -32.475 -194.995 ;
        RECT -32.805 -196.685 -32.475 -196.355 ;
        RECT -32.805 -198.045 -32.475 -197.715 ;
        RECT -32.805 -199.405 -32.475 -199.075 ;
        RECT -32.805 -200.765 -32.475 -200.435 ;
        RECT -32.805 -202.125 -32.475 -201.795 ;
        RECT -32.805 -203.485 -32.475 -203.155 ;
        RECT -32.805 -204.845 -32.475 -204.515 ;
        RECT -32.805 -206.555 -32.475 -206.225 ;
        RECT -32.805 -207.565 -32.475 -207.235 ;
        RECT -32.805 -208.925 -32.475 -208.595 ;
        RECT -32.805 -211.645 -32.475 -211.315 ;
        RECT -32.805 -214.365 -32.475 -214.035 ;
        RECT -32.805 -215.725 -32.475 -215.395 ;
        RECT -32.805 -217.085 -32.475 -216.755 ;
        RECT -32.805 -218.445 -32.475 -218.115 ;
        RECT -32.805 -224.09 -32.475 -222.96 ;
        RECT -32.8 -224.205 -32.48 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -31.445 37.235 -31.115 37.565 ;
        RECT -31.445 35.875 -31.115 36.205 ;
        RECT -31.445 34.515 -31.115 34.845 ;
        RECT -31.445 33.155 -31.115 33.485 ;
        RECT -31.445 31.795 -31.115 32.125 ;
        RECT -31.445 30.435 -31.115 30.765 ;
        RECT -31.445 29.075 -31.115 29.405 ;
        RECT -31.445 27.715 -31.115 28.045 ;
        RECT -31.445 26.355 -31.115 26.685 ;
        RECT -31.445 24.995 -31.115 25.325 ;
        RECT -31.445 23.635 -31.115 23.965 ;
        RECT -31.445 22.275 -31.115 22.605 ;
        RECT -31.445 20.915 -31.115 21.245 ;
        RECT -31.445 19.555 -31.115 19.885 ;
        RECT -31.445 18.195 -31.115 18.525 ;
        RECT -31.445 16.835 -31.115 17.165 ;
        RECT -31.445 15.475 -31.115 15.805 ;
        RECT -31.445 14.115 -31.115 14.445 ;
        RECT -31.445 12.755 -31.115 13.085 ;
        RECT -31.445 11.395 -31.115 11.725 ;
        RECT -31.445 10.035 -31.115 10.365 ;
        RECT -31.445 8.675 -31.115 9.005 ;
        RECT -31.445 7.315 -31.115 7.645 ;
        RECT -31.445 5.955 -31.115 6.285 ;
        RECT -31.445 4.595 -31.115 4.925 ;
        RECT -31.445 3.235 -31.115 3.565 ;
        RECT -31.445 1.875 -31.115 2.205 ;
        RECT -31.445 0.515 -31.115 0.845 ;
        RECT -31.445 -6.285 -31.115 -5.955 ;
        RECT -31.445 -7.645 -31.115 -7.315 ;
        RECT -31.445 -9.005 -31.115 -8.675 ;
        RECT -31.445 -11.725 -31.115 -11.395 ;
        RECT -31.445 -13.085 -31.115 -12.755 ;
        RECT -31.445 -14.445 -31.115 -14.115 ;
        RECT -31.445 -15.805 -31.115 -15.475 ;
        RECT -31.445 -17.165 -31.115 -16.835 ;
        RECT -31.445 -18.525 -31.115 -18.195 ;
        RECT -31.445 -19.885 -31.115 -19.555 ;
        RECT -31.445 -26.685 -31.115 -26.355 ;
        RECT -31.445 -28.045 -31.115 -27.715 ;
        RECT -31.445 -29.405 -31.115 -29.075 ;
        RECT -31.445 -32.125 -31.115 -31.795 ;
        RECT -31.445 -34.845 -31.115 -34.515 ;
        RECT -31.445 -37.565 -31.115 -37.235 ;
        RECT -31.445 -38.925 -31.115 -38.595 ;
        RECT -31.445 -40.285 -31.115 -39.955 ;
        RECT -31.445 -41.645 -31.115 -41.315 ;
        RECT -31.445 -43.005 -31.115 -42.675 ;
        RECT -31.445 -44.365 -31.115 -44.035 ;
        RECT -31.445 -45.725 -31.115 -45.395 ;
        RECT -31.445 -47.085 -31.115 -46.755 ;
        RECT -31.445 -48.445 -31.115 -48.115 ;
        RECT -31.445 -49.805 -31.115 -49.475 ;
        RECT -31.445 -51.165 -31.115 -50.835 ;
        RECT -31.445 -52.525 -31.115 -52.195 ;
        RECT -31.445 -53.885 -31.115 -53.555 ;
        RECT -31.445 -55.245 -31.115 -54.915 ;
        RECT -31.445 -56.605 -31.115 -56.275 ;
        RECT -31.445 -57.965 -31.115 -57.635 ;
        RECT -31.445 -59.325 -31.115 -58.995 ;
        RECT -31.445 -60.685 -31.115 -60.355 ;
        RECT -31.445 -62.045 -31.115 -61.715 ;
        RECT -31.445 -63.405 -31.115 -63.075 ;
        RECT -31.445 -64.765 -31.115 -64.435 ;
        RECT -31.445 -66.125 -31.115 -65.795 ;
        RECT -31.445 -67.485 -31.115 -67.155 ;
        RECT -31.445 -68.845 -31.115 -68.515 ;
        RECT -31.445 -70.205 -31.115 -69.875 ;
        RECT -31.445 -71.565 -31.115 -71.235 ;
        RECT -31.445 -72.925 -31.115 -72.595 ;
        RECT -31.445 -74.285 -31.115 -73.955 ;
        RECT -31.445 -75.645 -31.115 -75.315 ;
        RECT -31.445 -77.005 -31.115 -76.675 ;
        RECT -31.445 -78.365 -31.115 -78.035 ;
        RECT -31.445 -79.725 -31.115 -79.395 ;
        RECT -31.445 -81.085 -31.115 -80.755 ;
        RECT -31.445 -82.445 -31.115 -82.115 ;
        RECT -31.445 -83.805 -31.115 -83.475 ;
        RECT -31.445 -85.165 -31.115 -84.835 ;
        RECT -31.445 -86.525 -31.115 -86.195 ;
        RECT -31.445 -87.885 -31.115 -87.555 ;
        RECT -31.445 -89.245 -31.115 -88.915 ;
        RECT -31.445 -90.605 -31.115 -90.275 ;
        RECT -31.445 -91.965 -31.115 -91.635 ;
        RECT -31.445 -93.325 -31.115 -92.995 ;
        RECT -31.445 -94.685 -31.115 -94.355 ;
        RECT -31.445 -96.045 -31.115 -95.715 ;
        RECT -31.445 -97.405 -31.115 -97.075 ;
        RECT -31.445 -98.765 -31.115 -98.435 ;
        RECT -31.445 -100.125 -31.115 -99.795 ;
        RECT -31.445 -101.485 -31.115 -101.155 ;
        RECT -31.445 -102.845 -31.115 -102.515 ;
        RECT -31.445 -104.205 -31.115 -103.875 ;
        RECT -31.445 -105.565 -31.115 -105.235 ;
        RECT -31.445 -109.645 -31.115 -109.315 ;
        RECT -31.445 -111.005 -31.115 -110.675 ;
        RECT -31.445 -111.87 -31.115 -111.54 ;
        RECT -31.445 -113.725 -31.115 -113.395 ;
        RECT -31.445 -115.085 -31.115 -114.755 ;
        RECT -31.445 -116.445 -31.115 -116.115 ;
        RECT -31.445 -117.805 -31.115 -117.475 ;
        RECT -31.445 -120.525 -31.115 -120.195 ;
        RECT -31.445 -121.885 -31.115 -121.555 ;
        RECT -31.445 -123.245 -31.115 -122.915 ;
        RECT -31.445 -124.71 -31.115 -124.38 ;
        RECT -31.445 -125.965 -31.115 -125.635 ;
        RECT -31.445 -127.325 -31.115 -126.995 ;
        RECT -31.445 -130.045 -31.115 -129.715 ;
        RECT -31.445 -132.765 -31.115 -132.435 ;
        RECT -31.445 -134.125 -31.115 -133.795 ;
        RECT -31.445 -135.485 -31.115 -135.155 ;
        RECT -31.445 -136.845 -31.115 -136.515 ;
        RECT -31.445 -138.205 -31.115 -137.875 ;
        RECT -31.445 -139.565 -31.115 -139.235 ;
        RECT -31.445 -142.285 -31.115 -141.955 ;
        RECT -31.445 -143.645 -31.115 -143.315 ;
        RECT -31.445 -145.005 -31.115 -144.675 ;
        RECT -31.445 -146.365 -31.115 -146.035 ;
        RECT -31.445 -147.725 -31.115 -147.395 ;
        RECT -31.445 -149.085 -31.115 -148.755 ;
        RECT -31.445 -150.445 -31.115 -150.115 ;
        RECT -31.445 -151.805 -31.115 -151.475 ;
        RECT -31.445 -153.165 -31.115 -152.835 ;
        RECT -31.445 -154.525 -31.115 -154.195 ;
        RECT -31.445 -155.885 -31.115 -155.555 ;
        RECT -31.445 -157.245 -31.115 -156.915 ;
        RECT -31.445 -158.605 -31.115 -158.275 ;
        RECT -31.445 -159.965 -31.115 -159.635 ;
        RECT -31.445 -161.325 -31.115 -160.995 ;
        RECT -31.445 -162.685 -31.115 -162.355 ;
        RECT -31.445 -164.045 -31.115 -163.715 ;
        RECT -31.445 -165.405 -31.115 -165.075 ;
        RECT -31.445 -166.765 -31.115 -166.435 ;
        RECT -31.445 -170.845 -31.115 -170.515 ;
        RECT -31.445 -172.205 -31.115 -171.875 ;
        RECT -31.445 -173.565 -31.115 -173.235 ;
        RECT -31.445 -174.925 -31.115 -174.595 ;
        RECT -31.445 -176.285 -31.115 -175.955 ;
        RECT -31.445 -177.645 -31.115 -177.315 ;
        RECT -31.445 -179.005 -31.115 -178.675 ;
        RECT -31.445 -180.365 -31.115 -180.035 ;
        RECT -31.445 -181.725 -31.115 -181.395 ;
        RECT -31.445 -183.085 -31.115 -182.755 ;
        RECT -31.445 -184.445 -31.115 -184.115 ;
        RECT -31.445 -185.805 -31.115 -185.475 ;
        RECT -31.445 -188.525 -31.115 -188.195 ;
        RECT -31.445 -189.885 -31.115 -189.555 ;
        RECT -31.445 -193.965 -31.115 -193.635 ;
        RECT -31.445 -195.325 -31.115 -194.995 ;
        RECT -31.445 -196.685 -31.115 -196.355 ;
        RECT -31.445 -198.045 -31.115 -197.715 ;
        RECT -31.445 -199.405 -31.115 -199.075 ;
        RECT -31.445 -200.765 -31.115 -200.435 ;
        RECT -31.445 -202.125 -31.115 -201.795 ;
        RECT -31.445 -203.485 -31.115 -203.155 ;
        RECT -31.445 -204.845 -31.115 -204.515 ;
        RECT -31.445 -206.555 -31.115 -206.225 ;
        RECT -31.445 -207.565 -31.115 -207.235 ;
        RECT -31.445 -208.925 -31.115 -208.595 ;
        RECT -31.445 -210.285 -31.115 -209.955 ;
        RECT -31.445 -211.645 -31.115 -211.315 ;
        RECT -31.445 -214.365 -31.115 -214.035 ;
        RECT -31.445 -215.725 -31.115 -215.395 ;
        RECT -31.445 -217.085 -31.115 -216.755 ;
        RECT -31.445 -218.445 -31.115 -218.115 ;
        RECT -31.445 -224.09 -31.115 -222.96 ;
        RECT -31.44 -224.205 -31.12 133.765 ;
        RECT -31.445 132.52 -31.115 133.65 ;
        RECT -31.445 128.355 -31.115 128.685 ;
        RECT -31.445 126.995 -31.115 127.325 ;
        RECT -31.445 125.635 -31.115 125.965 ;
        RECT -31.445 124.275 -31.115 124.605 ;
        RECT -31.445 122.915 -31.115 123.245 ;
        RECT -31.445 121.555 -31.115 121.885 ;
        RECT -31.445 120.195 -31.115 120.525 ;
        RECT -31.445 118.835 -31.115 119.165 ;
        RECT -31.445 117.475 -31.115 117.805 ;
        RECT -31.445 116.115 -31.115 116.445 ;
        RECT -31.445 114.755 -31.115 115.085 ;
        RECT -31.445 113.395 -31.115 113.725 ;
        RECT -31.445 112.035 -31.115 112.365 ;
        RECT -31.445 110.675 -31.115 111.005 ;
        RECT -31.445 109.315 -31.115 109.645 ;
        RECT -31.445 107.955 -31.115 108.285 ;
        RECT -31.445 106.595 -31.115 106.925 ;
        RECT -31.445 105.235 -31.115 105.565 ;
        RECT -31.445 103.875 -31.115 104.205 ;
        RECT -31.445 102.515 -31.115 102.845 ;
        RECT -31.445 101.155 -31.115 101.485 ;
        RECT -31.445 99.795 -31.115 100.125 ;
        RECT -31.445 98.435 -31.115 98.765 ;
        RECT -31.445 97.075 -31.115 97.405 ;
        RECT -31.445 95.715 -31.115 96.045 ;
        RECT -31.445 94.355 -31.115 94.685 ;
        RECT -31.445 92.995 -31.115 93.325 ;
        RECT -31.445 91.635 -31.115 91.965 ;
        RECT -31.445 90.275 -31.115 90.605 ;
        RECT -31.445 88.915 -31.115 89.245 ;
        RECT -31.445 87.555 -31.115 87.885 ;
        RECT -31.445 86.195 -31.115 86.525 ;
        RECT -31.445 84.835 -31.115 85.165 ;
        RECT -31.445 83.475 -31.115 83.805 ;
        RECT -31.445 82.115 -31.115 82.445 ;
        RECT -31.445 80.755 -31.115 81.085 ;
        RECT -31.445 79.395 -31.115 79.725 ;
        RECT -31.445 78.035 -31.115 78.365 ;
        RECT -31.445 76.675 -31.115 77.005 ;
        RECT -31.445 75.315 -31.115 75.645 ;
        RECT -31.445 73.955 -31.115 74.285 ;
        RECT -31.445 72.595 -31.115 72.925 ;
        RECT -31.445 71.235 -31.115 71.565 ;
        RECT -31.445 69.875 -31.115 70.205 ;
        RECT -31.445 68.515 -31.115 68.845 ;
        RECT -31.445 67.155 -31.115 67.485 ;
        RECT -31.445 65.795 -31.115 66.125 ;
        RECT -31.445 64.435 -31.115 64.765 ;
        RECT -31.445 63.075 -31.115 63.405 ;
        RECT -31.445 61.715 -31.115 62.045 ;
        RECT -31.445 60.355 -31.115 60.685 ;
        RECT -31.445 58.995 -31.115 59.325 ;
        RECT -31.445 57.635 -31.115 57.965 ;
        RECT -31.445 56.275 -31.115 56.605 ;
        RECT -31.445 54.915 -31.115 55.245 ;
        RECT -31.445 53.555 -31.115 53.885 ;
        RECT -31.445 52.195 -31.115 52.525 ;
        RECT -31.445 50.835 -31.115 51.165 ;
        RECT -31.445 49.475 -31.115 49.805 ;
        RECT -31.445 48.115 -31.115 48.445 ;
        RECT -31.445 46.755 -31.115 47.085 ;
        RECT -31.445 45.395 -31.115 45.725 ;
        RECT -31.445 44.035 -31.115 44.365 ;
        RECT -31.445 42.675 -31.115 43.005 ;
        RECT -31.445 41.315 -31.115 41.645 ;
        RECT -31.445 39.955 -31.115 40.285 ;
        RECT -31.445 38.595 -31.115 38.925 ;
    END
    PORT
      LAYER met3 ;
        RECT -40.965 132.52 -40.635 133.65 ;
        RECT -40.965 128.355 -40.635 128.685 ;
        RECT -40.965 126.995 -40.635 127.325 ;
        RECT -40.965 125.635 -40.635 125.965 ;
        RECT -40.965 124.275 -40.635 124.605 ;
        RECT -40.965 122.915 -40.635 123.245 ;
        RECT -40.965 121.555 -40.635 121.885 ;
        RECT -40.965 120.195 -40.635 120.525 ;
        RECT -40.965 118.835 -40.635 119.165 ;
        RECT -40.965 117.475 -40.635 117.805 ;
        RECT -40.965 116.115 -40.635 116.445 ;
        RECT -40.965 114.755 -40.635 115.085 ;
        RECT -40.965 113.395 -40.635 113.725 ;
        RECT -40.965 112.035 -40.635 112.365 ;
        RECT -40.965 110.675 -40.635 111.005 ;
        RECT -40.965 109.315 -40.635 109.645 ;
        RECT -40.965 107.955 -40.635 108.285 ;
        RECT -40.965 106.595 -40.635 106.925 ;
        RECT -40.965 105.235 -40.635 105.565 ;
        RECT -40.965 103.875 -40.635 104.205 ;
        RECT -40.965 102.515 -40.635 102.845 ;
        RECT -40.965 101.155 -40.635 101.485 ;
        RECT -40.965 99.795 -40.635 100.125 ;
        RECT -40.965 98.435 -40.635 98.765 ;
        RECT -40.965 97.075 -40.635 97.405 ;
        RECT -40.965 95.715 -40.635 96.045 ;
        RECT -40.965 94.355 -40.635 94.685 ;
        RECT -40.965 92.995 -40.635 93.325 ;
        RECT -40.965 91.635 -40.635 91.965 ;
        RECT -40.965 90.275 -40.635 90.605 ;
        RECT -40.965 88.915 -40.635 89.245 ;
        RECT -40.965 87.555 -40.635 87.885 ;
        RECT -40.965 86.195 -40.635 86.525 ;
        RECT -40.965 84.835 -40.635 85.165 ;
        RECT -40.965 83.475 -40.635 83.805 ;
        RECT -40.965 82.115 -40.635 82.445 ;
        RECT -40.965 80.755 -40.635 81.085 ;
        RECT -40.965 79.395 -40.635 79.725 ;
        RECT -40.965 78.035 -40.635 78.365 ;
        RECT -40.965 76.675 -40.635 77.005 ;
        RECT -40.965 75.315 -40.635 75.645 ;
        RECT -40.965 73.955 -40.635 74.285 ;
        RECT -40.965 71.64 -40.635 71.97 ;
        RECT -40.965 69.465 -40.635 69.795 ;
        RECT -40.965 68.615 -40.635 68.945 ;
        RECT -40.965 66.305 -40.635 66.635 ;
        RECT -40.965 65.455 -40.635 65.785 ;
        RECT -40.965 63.145 -40.635 63.475 ;
        RECT -40.965 62.295 -40.635 62.625 ;
        RECT -40.965 59.985 -40.635 60.315 ;
        RECT -40.965 59.135 -40.635 59.465 ;
        RECT -40.965 56.825 -40.635 57.155 ;
        RECT -40.965 55.975 -40.635 56.305 ;
        RECT -40.965 53.665 -40.635 53.995 ;
        RECT -40.965 52.815 -40.635 53.145 ;
        RECT -40.965 50.64 -40.635 50.97 ;
        RECT -40.965 48.115 -40.635 48.445 ;
        RECT -40.965 46.755 -40.635 47.085 ;
        RECT -40.965 45.395 -40.635 45.725 ;
        RECT -40.965 44.035 -40.635 44.365 ;
        RECT -40.965 42.675 -40.635 43.005 ;
        RECT -40.965 41.315 -40.635 41.645 ;
        RECT -40.965 39.955 -40.635 40.285 ;
        RECT -40.965 38.595 -40.635 38.925 ;
        RECT -40.965 37.235 -40.635 37.565 ;
        RECT -40.965 35.875 -40.635 36.205 ;
        RECT -40.965 34.515 -40.635 34.845 ;
        RECT -40.965 33.155 -40.635 33.485 ;
        RECT -40.965 31.795 -40.635 32.125 ;
        RECT -40.965 30.435 -40.635 30.765 ;
        RECT -40.965 29.075 -40.635 29.405 ;
        RECT -40.965 27.715 -40.635 28.045 ;
        RECT -40.965 26.355 -40.635 26.685 ;
        RECT -40.965 24.995 -40.635 25.325 ;
        RECT -40.965 23.635 -40.635 23.965 ;
        RECT -40.965 22.275 -40.635 22.605 ;
        RECT -40.965 20.915 -40.635 21.245 ;
        RECT -40.965 19.555 -40.635 19.885 ;
        RECT -40.965 18.195 -40.635 18.525 ;
        RECT -40.965 16.835 -40.635 17.165 ;
        RECT -40.965 15.475 -40.635 15.805 ;
        RECT -40.965 14.115 -40.635 14.445 ;
        RECT -40.965 12.755 -40.635 13.085 ;
        RECT -40.965 11.395 -40.635 11.725 ;
        RECT -40.965 10.035 -40.635 10.365 ;
        RECT -40.965 8.675 -40.635 9.005 ;
        RECT -40.965 7.315 -40.635 7.645 ;
        RECT -40.965 5.955 -40.635 6.285 ;
        RECT -40.965 4.595 -40.635 4.925 ;
        RECT -40.965 3.235 -40.635 3.565 ;
        RECT -40.965 1.875 -40.635 2.205 ;
        RECT -40.965 0.515 -40.635 0.845 ;
        RECT -40.965 -0.845 -40.635 -0.515 ;
        RECT -40.965 -2.205 -40.635 -1.875 ;
        RECT -40.965 -3.565 -40.635 -3.235 ;
        RECT -40.965 -4.925 -40.635 -4.595 ;
        RECT -40.965 -6.285 -40.635 -5.955 ;
        RECT -40.965 -7.645 -40.635 -7.315 ;
        RECT -40.965 -9.005 -40.635 -8.675 ;
        RECT -40.965 -11.725 -40.635 -11.395 ;
        RECT -40.965 -13.085 -40.635 -12.755 ;
        RECT -40.965 -14.445 -40.635 -14.115 ;
        RECT -40.965 -15.805 -40.635 -15.475 ;
        RECT -40.965 -17.165 -40.635 -16.835 ;
        RECT -40.965 -18.525 -40.635 -18.195 ;
        RECT -40.965 -19.885 -40.635 -19.555 ;
        RECT -40.965 -21.245 -40.635 -20.915 ;
        RECT -40.965 -22.605 -40.635 -22.275 ;
        RECT -40.965 -26.685 -40.635 -26.355 ;
        RECT -40.965 -28.045 -40.635 -27.715 ;
        RECT -40.965 -29.405 -40.635 -29.075 ;
        RECT -40.965 -32.125 -40.635 -31.795 ;
        RECT -40.965 -34.845 -40.635 -34.515 ;
        RECT -40.965 -37.565 -40.635 -37.235 ;
        RECT -40.965 -38.925 -40.635 -38.595 ;
        RECT -40.965 -40.285 -40.635 -39.955 ;
        RECT -40.965 -41.645 -40.635 -41.315 ;
        RECT -40.965 -43.005 -40.635 -42.675 ;
        RECT -40.965 -44.365 -40.635 -44.035 ;
        RECT -40.965 -45.725 -40.635 -45.395 ;
        RECT -40.965 -47.085 -40.635 -46.755 ;
        RECT -40.965 -48.445 -40.635 -48.115 ;
        RECT -40.965 -49.805 -40.635 -49.475 ;
        RECT -40.965 -51.165 -40.635 -50.835 ;
        RECT -40.965 -52.525 -40.635 -52.195 ;
        RECT -40.965 -53.885 -40.635 -53.555 ;
        RECT -40.965 -55.245 -40.635 -54.915 ;
        RECT -40.965 -56.605 -40.635 -56.275 ;
        RECT -40.965 -57.965 -40.635 -57.635 ;
        RECT -40.965 -59.325 -40.635 -58.995 ;
        RECT -40.965 -60.685 -40.635 -60.355 ;
        RECT -40.965 -62.045 -40.635 -61.715 ;
        RECT -40.965 -63.405 -40.635 -63.075 ;
        RECT -40.965 -64.765 -40.635 -64.435 ;
        RECT -40.965 -66.125 -40.635 -65.795 ;
        RECT -40.965 -67.485 -40.635 -67.155 ;
        RECT -40.965 -68.845 -40.635 -68.515 ;
        RECT -40.965 -70.205 -40.635 -69.875 ;
        RECT -40.965 -71.565 -40.635 -71.235 ;
        RECT -40.965 -72.925 -40.635 -72.595 ;
        RECT -40.965 -74.285 -40.635 -73.955 ;
        RECT -40.965 -75.645 -40.635 -75.315 ;
        RECT -40.965 -77.005 -40.635 -76.675 ;
        RECT -40.965 -78.365 -40.635 -78.035 ;
        RECT -40.965 -79.725 -40.635 -79.395 ;
        RECT -40.965 -81.085 -40.635 -80.755 ;
        RECT -40.965 -82.445 -40.635 -82.115 ;
        RECT -40.965 -83.805 -40.635 -83.475 ;
        RECT -40.965 -85.165 -40.635 -84.835 ;
        RECT -40.965 -86.525 -40.635 -86.195 ;
        RECT -40.965 -87.885 -40.635 -87.555 ;
        RECT -40.965 -89.245 -40.635 -88.915 ;
        RECT -40.965 -90.605 -40.635 -90.275 ;
        RECT -40.965 -91.965 -40.635 -91.635 ;
        RECT -40.965 -93.325 -40.635 -92.995 ;
        RECT -40.965 -94.685 -40.635 -94.355 ;
        RECT -40.965 -96.045 -40.635 -95.715 ;
        RECT -40.965 -97.405 -40.635 -97.075 ;
        RECT -40.965 -98.765 -40.635 -98.435 ;
        RECT -40.965 -100.125 -40.635 -99.795 ;
        RECT -40.965 -101.485 -40.635 -101.155 ;
        RECT -40.965 -102.845 -40.635 -102.515 ;
        RECT -40.965 -104.205 -40.635 -103.875 ;
        RECT -40.965 -105.565 -40.635 -105.235 ;
        RECT -40.965 -106.925 -40.635 -106.595 ;
        RECT -40.965 -108.285 -40.635 -107.955 ;
        RECT -40.965 -109.645 -40.635 -109.315 ;
        RECT -40.965 -111.005 -40.635 -110.675 ;
        RECT -40.965 -111.87 -40.635 -111.54 ;
        RECT -40.965 -113.725 -40.635 -113.395 ;
        RECT -40.965 -115.085 -40.635 -114.755 ;
        RECT -40.965 -116.445 -40.635 -116.115 ;
        RECT -40.965 -117.805 -40.635 -117.475 ;
        RECT -40.965 -120.525 -40.635 -120.195 ;
        RECT -40.965 -121.885 -40.635 -121.555 ;
        RECT -40.965 -123.245 -40.635 -122.915 ;
        RECT -40.965 -124.71 -40.635 -124.38 ;
        RECT -40.965 -125.965 -40.635 -125.635 ;
        RECT -40.965 -127.325 -40.635 -126.995 ;
        RECT -40.965 -130.045 -40.635 -129.715 ;
        RECT -40.965 -134.125 -40.635 -133.795 ;
        RECT -40.965 -135.485 -40.635 -135.155 ;
        RECT -40.965 -136.845 -40.635 -136.515 ;
        RECT -40.965 -138.205 -40.635 -137.875 ;
        RECT -40.965 -139.565 -40.635 -139.235 ;
        RECT -40.965 -142.285 -40.635 -141.955 ;
        RECT -40.965 -143.645 -40.635 -143.315 ;
        RECT -40.965 -145.005 -40.635 -144.675 ;
        RECT -40.965 -146.365 -40.635 -146.035 ;
        RECT -40.965 -147.725 -40.635 -147.395 ;
        RECT -40.965 -149.085 -40.635 -148.755 ;
        RECT -40.965 -150.445 -40.635 -150.115 ;
        RECT -40.965 -151.805 -40.635 -151.475 ;
        RECT -40.965 -153.165 -40.635 -152.835 ;
        RECT -40.965 -154.525 -40.635 -154.195 ;
        RECT -40.965 -155.885 -40.635 -155.555 ;
        RECT -40.965 -157.245 -40.635 -156.915 ;
        RECT -40.965 -158.605 -40.635 -158.275 ;
        RECT -40.965 -159.965 -40.635 -159.635 ;
        RECT -40.965 -161.325 -40.635 -160.995 ;
        RECT -40.965 -162.685 -40.635 -162.355 ;
        RECT -40.965 -164.045 -40.635 -163.715 ;
        RECT -40.965 -165.405 -40.635 -165.075 ;
        RECT -40.965 -166.765 -40.635 -166.435 ;
        RECT -40.965 -168.125 -40.635 -167.795 ;
        RECT -40.965 -169.485 -40.635 -169.155 ;
        RECT -40.965 -170.845 -40.635 -170.515 ;
        RECT -40.965 -172.205 -40.635 -171.875 ;
        RECT -40.965 -173.565 -40.635 -173.235 ;
        RECT -40.965 -174.925 -40.635 -174.595 ;
        RECT -40.965 -176.285 -40.635 -175.955 ;
        RECT -40.965 -177.645 -40.635 -177.315 ;
        RECT -40.965 -179.005 -40.635 -178.675 ;
        RECT -40.965 -180.365 -40.635 -180.035 ;
        RECT -40.965 -181.725 -40.635 -181.395 ;
        RECT -40.965 -183.085 -40.635 -182.755 ;
        RECT -40.965 -184.445 -40.635 -184.115 ;
        RECT -40.965 -185.805 -40.635 -185.475 ;
        RECT -40.965 -187.165 -40.635 -186.835 ;
        RECT -40.965 -188.525 -40.635 -188.195 ;
        RECT -40.965 -189.885 -40.635 -189.555 ;
        RECT -40.965 -191.245 -40.635 -190.915 ;
        RECT -40.965 -192.605 -40.635 -192.275 ;
        RECT -40.965 -193.965 -40.635 -193.635 ;
        RECT -40.965 -195.325 -40.635 -194.995 ;
        RECT -40.965 -196.685 -40.635 -196.355 ;
        RECT -40.965 -198.045 -40.635 -197.715 ;
        RECT -40.965 -199.405 -40.635 -199.075 ;
        RECT -40.965 -200.765 -40.635 -200.435 ;
        RECT -40.965 -202.125 -40.635 -201.795 ;
        RECT -40.965 -203.485 -40.635 -203.155 ;
        RECT -40.965 -204.845 -40.635 -204.515 ;
        RECT -40.965 -207.565 -40.635 -207.235 ;
        RECT -40.965 -208.925 -40.635 -208.595 ;
        RECT -40.965 -214.365 -40.635 -214.035 ;
        RECT -40.965 -215.725 -40.635 -215.395 ;
        RECT -40.965 -217.085 -40.635 -216.755 ;
        RECT -40.965 -218.445 -40.635 -218.115 ;
        RECT -40.965 -224.09 -40.635 -222.96 ;
        RECT -40.96 -224.205 -40.64 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -39.605 132.52 -39.275 133.65 ;
        RECT -39.605 128.355 -39.275 128.685 ;
        RECT -39.605 126.995 -39.275 127.325 ;
        RECT -39.605 125.635 -39.275 125.965 ;
        RECT -39.605 124.275 -39.275 124.605 ;
        RECT -39.605 122.915 -39.275 123.245 ;
        RECT -39.605 121.555 -39.275 121.885 ;
        RECT -39.605 120.195 -39.275 120.525 ;
        RECT -39.605 118.835 -39.275 119.165 ;
        RECT -39.605 117.475 -39.275 117.805 ;
        RECT -39.605 116.115 -39.275 116.445 ;
        RECT -39.605 114.755 -39.275 115.085 ;
        RECT -39.605 113.395 -39.275 113.725 ;
        RECT -39.605 112.035 -39.275 112.365 ;
        RECT -39.605 110.675 -39.275 111.005 ;
        RECT -39.605 109.315 -39.275 109.645 ;
        RECT -39.605 107.955 -39.275 108.285 ;
        RECT -39.605 106.595 -39.275 106.925 ;
        RECT -39.605 105.235 -39.275 105.565 ;
        RECT -39.605 103.875 -39.275 104.205 ;
        RECT -39.605 102.515 -39.275 102.845 ;
        RECT -39.605 101.155 -39.275 101.485 ;
        RECT -39.605 99.795 -39.275 100.125 ;
        RECT -39.605 98.435 -39.275 98.765 ;
        RECT -39.605 97.075 -39.275 97.405 ;
        RECT -39.605 95.715 -39.275 96.045 ;
        RECT -39.605 94.355 -39.275 94.685 ;
        RECT -39.605 92.995 -39.275 93.325 ;
        RECT -39.605 91.635 -39.275 91.965 ;
        RECT -39.605 90.275 -39.275 90.605 ;
        RECT -39.605 88.915 -39.275 89.245 ;
        RECT -39.605 87.555 -39.275 87.885 ;
        RECT -39.605 86.195 -39.275 86.525 ;
        RECT -39.605 84.835 -39.275 85.165 ;
        RECT -39.605 83.475 -39.275 83.805 ;
        RECT -39.605 82.115 -39.275 82.445 ;
        RECT -39.605 80.755 -39.275 81.085 ;
        RECT -39.605 79.395 -39.275 79.725 ;
        RECT -39.605 78.035 -39.275 78.365 ;
        RECT -39.605 76.675 -39.275 77.005 ;
        RECT -39.605 75.315 -39.275 75.645 ;
        RECT -39.605 73.955 -39.275 74.285 ;
        RECT -39.605 72.595 -39.275 72.925 ;
        RECT -39.605 71.235 -39.275 71.565 ;
        RECT -39.605 69.875 -39.275 70.205 ;
        RECT -39.605 68.515 -39.275 68.845 ;
        RECT -39.605 67.155 -39.275 67.485 ;
        RECT -39.605 65.795 -39.275 66.125 ;
        RECT -39.605 64.435 -39.275 64.765 ;
        RECT -39.605 63.075 -39.275 63.405 ;
        RECT -39.605 61.715 -39.275 62.045 ;
        RECT -39.605 60.355 -39.275 60.685 ;
        RECT -39.605 58.995 -39.275 59.325 ;
        RECT -39.605 57.635 -39.275 57.965 ;
        RECT -39.605 56.275 -39.275 56.605 ;
        RECT -39.605 54.915 -39.275 55.245 ;
        RECT -39.605 53.555 -39.275 53.885 ;
        RECT -39.605 52.195 -39.275 52.525 ;
        RECT -39.605 50.835 -39.275 51.165 ;
        RECT -39.605 49.475 -39.275 49.805 ;
        RECT -39.605 48.115 -39.275 48.445 ;
        RECT -39.605 46.755 -39.275 47.085 ;
        RECT -39.605 45.395 -39.275 45.725 ;
        RECT -39.605 44.035 -39.275 44.365 ;
        RECT -39.605 42.675 -39.275 43.005 ;
        RECT -39.605 41.315 -39.275 41.645 ;
        RECT -39.605 39.955 -39.275 40.285 ;
        RECT -39.605 38.595 -39.275 38.925 ;
        RECT -39.605 37.235 -39.275 37.565 ;
        RECT -39.605 35.875 -39.275 36.205 ;
        RECT -39.605 34.515 -39.275 34.845 ;
        RECT -39.605 33.155 -39.275 33.485 ;
        RECT -39.605 31.795 -39.275 32.125 ;
        RECT -39.605 30.435 -39.275 30.765 ;
        RECT -39.605 29.075 -39.275 29.405 ;
        RECT -39.605 27.715 -39.275 28.045 ;
        RECT -39.605 26.355 -39.275 26.685 ;
        RECT -39.605 24.995 -39.275 25.325 ;
        RECT -39.605 23.635 -39.275 23.965 ;
        RECT -39.605 22.275 -39.275 22.605 ;
        RECT -39.605 20.915 -39.275 21.245 ;
        RECT -39.605 19.555 -39.275 19.885 ;
        RECT -39.605 18.195 -39.275 18.525 ;
        RECT -39.605 16.835 -39.275 17.165 ;
        RECT -39.605 15.475 -39.275 15.805 ;
        RECT -39.605 14.115 -39.275 14.445 ;
        RECT -39.605 12.755 -39.275 13.085 ;
        RECT -39.605 11.395 -39.275 11.725 ;
        RECT -39.605 10.035 -39.275 10.365 ;
        RECT -39.605 8.675 -39.275 9.005 ;
        RECT -39.605 7.315 -39.275 7.645 ;
        RECT -39.605 5.955 -39.275 6.285 ;
        RECT -39.605 4.595 -39.275 4.925 ;
        RECT -39.605 3.235 -39.275 3.565 ;
        RECT -39.605 1.875 -39.275 2.205 ;
        RECT -39.605 0.515 -39.275 0.845 ;
        RECT -39.605 -0.845 -39.275 -0.515 ;
        RECT -39.605 -2.205 -39.275 -1.875 ;
        RECT -39.605 -3.565 -39.275 -3.235 ;
        RECT -39.605 -4.925 -39.275 -4.595 ;
        RECT -39.605 -6.285 -39.275 -5.955 ;
        RECT -39.605 -7.645 -39.275 -7.315 ;
        RECT -39.605 -9.005 -39.275 -8.675 ;
        RECT -39.605 -11.725 -39.275 -11.395 ;
        RECT -39.605 -13.085 -39.275 -12.755 ;
        RECT -39.605 -14.445 -39.275 -14.115 ;
        RECT -39.605 -15.805 -39.275 -15.475 ;
        RECT -39.605 -17.165 -39.275 -16.835 ;
        RECT -39.605 -18.525 -39.275 -18.195 ;
        RECT -39.605 -19.885 -39.275 -19.555 ;
        RECT -39.605 -21.245 -39.275 -20.915 ;
        RECT -39.605 -26.685 -39.275 -26.355 ;
        RECT -39.605 -28.045 -39.275 -27.715 ;
        RECT -39.605 -29.405 -39.275 -29.075 ;
        RECT -39.605 -32.125 -39.275 -31.795 ;
        RECT -39.605 -34.845 -39.275 -34.515 ;
        RECT -39.605 -37.565 -39.275 -37.235 ;
        RECT -39.605 -38.925 -39.275 -38.595 ;
        RECT -39.605 -40.285 -39.275 -39.955 ;
        RECT -39.605 -41.645 -39.275 -41.315 ;
        RECT -39.605 -43.005 -39.275 -42.675 ;
        RECT -39.605 -44.365 -39.275 -44.035 ;
        RECT -39.605 -45.725 -39.275 -45.395 ;
        RECT -39.605 -47.085 -39.275 -46.755 ;
        RECT -39.605 -48.445 -39.275 -48.115 ;
        RECT -39.605 -49.805 -39.275 -49.475 ;
        RECT -39.605 -51.165 -39.275 -50.835 ;
        RECT -39.605 -52.525 -39.275 -52.195 ;
        RECT -39.605 -53.885 -39.275 -53.555 ;
        RECT -39.605 -55.245 -39.275 -54.915 ;
        RECT -39.605 -56.605 -39.275 -56.275 ;
        RECT -39.605 -57.965 -39.275 -57.635 ;
        RECT -39.605 -59.325 -39.275 -58.995 ;
        RECT -39.605 -60.685 -39.275 -60.355 ;
        RECT -39.605 -62.045 -39.275 -61.715 ;
        RECT -39.605 -63.405 -39.275 -63.075 ;
        RECT -39.605 -64.765 -39.275 -64.435 ;
        RECT -39.605 -66.125 -39.275 -65.795 ;
        RECT -39.605 -67.485 -39.275 -67.155 ;
        RECT -39.605 -68.845 -39.275 -68.515 ;
        RECT -39.605 -70.205 -39.275 -69.875 ;
        RECT -39.605 -71.565 -39.275 -71.235 ;
        RECT -39.605 -72.925 -39.275 -72.595 ;
        RECT -39.605 -74.285 -39.275 -73.955 ;
        RECT -39.605 -75.645 -39.275 -75.315 ;
        RECT -39.605 -77.005 -39.275 -76.675 ;
        RECT -39.605 -78.365 -39.275 -78.035 ;
        RECT -39.605 -79.725 -39.275 -79.395 ;
        RECT -39.605 -81.085 -39.275 -80.755 ;
        RECT -39.605 -82.445 -39.275 -82.115 ;
        RECT -39.605 -83.805 -39.275 -83.475 ;
        RECT -39.605 -85.165 -39.275 -84.835 ;
        RECT -39.605 -86.525 -39.275 -86.195 ;
        RECT -39.605 -87.885 -39.275 -87.555 ;
        RECT -39.605 -89.245 -39.275 -88.915 ;
        RECT -39.605 -90.605 -39.275 -90.275 ;
        RECT -39.605 -91.965 -39.275 -91.635 ;
        RECT -39.605 -93.325 -39.275 -92.995 ;
        RECT -39.605 -94.685 -39.275 -94.355 ;
        RECT -39.605 -96.045 -39.275 -95.715 ;
        RECT -39.605 -97.405 -39.275 -97.075 ;
        RECT -39.605 -98.765 -39.275 -98.435 ;
        RECT -39.605 -100.125 -39.275 -99.795 ;
        RECT -39.605 -101.485 -39.275 -101.155 ;
        RECT -39.605 -102.845 -39.275 -102.515 ;
        RECT -39.605 -104.205 -39.275 -103.875 ;
        RECT -39.605 -105.565 -39.275 -105.235 ;
        RECT -39.605 -106.925 -39.275 -106.595 ;
        RECT -39.605 -109.645 -39.275 -109.315 ;
        RECT -39.605 -111.005 -39.275 -110.675 ;
        RECT -39.605 -111.87 -39.275 -111.54 ;
        RECT -39.605 -113.725 -39.275 -113.395 ;
        RECT -39.605 -115.085 -39.275 -114.755 ;
        RECT -39.605 -116.445 -39.275 -116.115 ;
        RECT -39.605 -117.805 -39.275 -117.475 ;
        RECT -39.605 -120.525 -39.275 -120.195 ;
        RECT -39.605 -121.885 -39.275 -121.555 ;
        RECT -39.605 -123.245 -39.275 -122.915 ;
        RECT -39.605 -124.71 -39.275 -124.38 ;
        RECT -39.605 -125.965 -39.275 -125.635 ;
        RECT -39.605 -127.325 -39.275 -126.995 ;
        RECT -39.605 -130.045 -39.275 -129.715 ;
        RECT -39.605 -134.125 -39.275 -133.795 ;
        RECT -39.605 -135.485 -39.275 -135.155 ;
        RECT -39.605 -136.845 -39.275 -136.515 ;
        RECT -39.605 -138.205 -39.275 -137.875 ;
        RECT -39.605 -139.565 -39.275 -139.235 ;
        RECT -39.605 -142.285 -39.275 -141.955 ;
        RECT -39.605 -143.645 -39.275 -143.315 ;
        RECT -39.605 -145.005 -39.275 -144.675 ;
        RECT -39.605 -146.365 -39.275 -146.035 ;
        RECT -39.605 -147.725 -39.275 -147.395 ;
        RECT -39.605 -149.085 -39.275 -148.755 ;
        RECT -39.605 -150.445 -39.275 -150.115 ;
        RECT -39.605 -151.805 -39.275 -151.475 ;
        RECT -39.605 -153.165 -39.275 -152.835 ;
        RECT -39.605 -154.525 -39.275 -154.195 ;
        RECT -39.605 -155.885 -39.275 -155.555 ;
        RECT -39.605 -157.245 -39.275 -156.915 ;
        RECT -39.605 -158.605 -39.275 -158.275 ;
        RECT -39.605 -159.965 -39.275 -159.635 ;
        RECT -39.605 -161.325 -39.275 -160.995 ;
        RECT -39.605 -162.685 -39.275 -162.355 ;
        RECT -39.605 -164.045 -39.275 -163.715 ;
        RECT -39.605 -165.405 -39.275 -165.075 ;
        RECT -39.605 -166.765 -39.275 -166.435 ;
        RECT -39.605 -168.125 -39.275 -167.795 ;
        RECT -39.605 -169.485 -39.275 -169.155 ;
        RECT -39.605 -170.845 -39.275 -170.515 ;
        RECT -39.605 -172.205 -39.275 -171.875 ;
        RECT -39.605 -173.565 -39.275 -173.235 ;
        RECT -39.605 -174.925 -39.275 -174.595 ;
        RECT -39.605 -176.285 -39.275 -175.955 ;
        RECT -39.605 -177.645 -39.275 -177.315 ;
        RECT -39.605 -179.005 -39.275 -178.675 ;
        RECT -39.605 -180.365 -39.275 -180.035 ;
        RECT -39.605 -181.725 -39.275 -181.395 ;
        RECT -39.605 -183.085 -39.275 -182.755 ;
        RECT -39.605 -184.445 -39.275 -184.115 ;
        RECT -39.605 -185.805 -39.275 -185.475 ;
        RECT -39.605 -187.165 -39.275 -186.835 ;
        RECT -39.605 -188.525 -39.275 -188.195 ;
        RECT -39.605 -189.885 -39.275 -189.555 ;
        RECT -39.605 -191.245 -39.275 -190.915 ;
        RECT -39.605 -192.605 -39.275 -192.275 ;
        RECT -39.605 -193.965 -39.275 -193.635 ;
        RECT -39.605 -195.325 -39.275 -194.995 ;
        RECT -39.605 -196.685 -39.275 -196.355 ;
        RECT -39.605 -198.045 -39.275 -197.715 ;
        RECT -39.605 -199.405 -39.275 -199.075 ;
        RECT -39.605 -200.765 -39.275 -200.435 ;
        RECT -39.605 -202.125 -39.275 -201.795 ;
        RECT -39.605 -203.485 -39.275 -203.155 ;
        RECT -39.605 -204.845 -39.275 -204.515 ;
        RECT -39.605 -206.555 -39.275 -206.225 ;
        RECT -39.605 -207.565 -39.275 -207.235 ;
        RECT -39.605 -208.925 -39.275 -208.595 ;
        RECT -39.605 -214.365 -39.275 -214.035 ;
        RECT -39.605 -215.725 -39.275 -215.395 ;
        RECT -39.605 -217.085 -39.275 -216.755 ;
        RECT -39.605 -218.445 -39.275 -218.115 ;
        RECT -39.605 -224.09 -39.275 -222.96 ;
        RECT -39.6 -224.205 -39.28 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.245 132.52 -37.915 133.65 ;
        RECT -38.245 128.355 -37.915 128.685 ;
        RECT -38.245 126.995 -37.915 127.325 ;
        RECT -38.245 125.635 -37.915 125.965 ;
        RECT -38.245 124.275 -37.915 124.605 ;
        RECT -38.245 122.915 -37.915 123.245 ;
        RECT -38.245 121.555 -37.915 121.885 ;
        RECT -38.245 120.195 -37.915 120.525 ;
        RECT -38.245 118.835 -37.915 119.165 ;
        RECT -38.245 117.475 -37.915 117.805 ;
        RECT -38.245 116.115 -37.915 116.445 ;
        RECT -38.245 114.755 -37.915 115.085 ;
        RECT -38.245 113.395 -37.915 113.725 ;
        RECT -38.245 112.035 -37.915 112.365 ;
        RECT -38.245 110.675 -37.915 111.005 ;
        RECT -38.245 109.315 -37.915 109.645 ;
        RECT -38.245 107.955 -37.915 108.285 ;
        RECT -38.245 106.595 -37.915 106.925 ;
        RECT -38.245 105.235 -37.915 105.565 ;
        RECT -38.245 103.875 -37.915 104.205 ;
        RECT -38.245 102.515 -37.915 102.845 ;
        RECT -38.245 101.155 -37.915 101.485 ;
        RECT -38.245 99.795 -37.915 100.125 ;
        RECT -38.245 98.435 -37.915 98.765 ;
        RECT -38.245 97.075 -37.915 97.405 ;
        RECT -38.245 95.715 -37.915 96.045 ;
        RECT -38.245 94.355 -37.915 94.685 ;
        RECT -38.245 92.995 -37.915 93.325 ;
        RECT -38.245 91.635 -37.915 91.965 ;
        RECT -38.245 90.275 -37.915 90.605 ;
        RECT -38.245 88.915 -37.915 89.245 ;
        RECT -38.245 87.555 -37.915 87.885 ;
        RECT -38.245 86.195 -37.915 86.525 ;
        RECT -38.245 84.835 -37.915 85.165 ;
        RECT -38.245 83.475 -37.915 83.805 ;
        RECT -38.245 82.115 -37.915 82.445 ;
        RECT -38.245 80.755 -37.915 81.085 ;
        RECT -38.245 79.395 -37.915 79.725 ;
        RECT -38.245 78.035 -37.915 78.365 ;
        RECT -38.245 76.675 -37.915 77.005 ;
        RECT -38.245 75.315 -37.915 75.645 ;
        RECT -38.245 73.955 -37.915 74.285 ;
        RECT -38.245 72.595 -37.915 72.925 ;
        RECT -38.245 71.235 -37.915 71.565 ;
        RECT -38.245 69.875 -37.915 70.205 ;
        RECT -38.245 68.515 -37.915 68.845 ;
        RECT -38.245 67.155 -37.915 67.485 ;
        RECT -38.245 65.795 -37.915 66.125 ;
        RECT -38.245 64.435 -37.915 64.765 ;
        RECT -38.245 63.075 -37.915 63.405 ;
        RECT -38.245 61.715 -37.915 62.045 ;
        RECT -38.245 60.355 -37.915 60.685 ;
        RECT -38.245 58.995 -37.915 59.325 ;
        RECT -38.245 57.635 -37.915 57.965 ;
        RECT -38.245 56.275 -37.915 56.605 ;
        RECT -38.245 54.915 -37.915 55.245 ;
        RECT -38.245 53.555 -37.915 53.885 ;
        RECT -38.245 52.195 -37.915 52.525 ;
        RECT -38.245 50.835 -37.915 51.165 ;
        RECT -38.245 49.475 -37.915 49.805 ;
        RECT -38.245 48.115 -37.915 48.445 ;
        RECT -38.245 46.755 -37.915 47.085 ;
        RECT -38.245 45.395 -37.915 45.725 ;
        RECT -38.245 44.035 -37.915 44.365 ;
        RECT -38.245 42.675 -37.915 43.005 ;
        RECT -38.245 41.315 -37.915 41.645 ;
        RECT -38.245 39.955 -37.915 40.285 ;
        RECT -38.245 38.595 -37.915 38.925 ;
        RECT -38.245 37.235 -37.915 37.565 ;
        RECT -38.245 35.875 -37.915 36.205 ;
        RECT -38.245 34.515 -37.915 34.845 ;
        RECT -38.245 33.155 -37.915 33.485 ;
        RECT -38.245 31.795 -37.915 32.125 ;
        RECT -38.245 30.435 -37.915 30.765 ;
        RECT -38.245 29.075 -37.915 29.405 ;
        RECT -38.245 27.715 -37.915 28.045 ;
        RECT -38.245 26.355 -37.915 26.685 ;
        RECT -38.245 24.995 -37.915 25.325 ;
        RECT -38.245 23.635 -37.915 23.965 ;
        RECT -38.245 22.275 -37.915 22.605 ;
        RECT -38.245 20.915 -37.915 21.245 ;
        RECT -38.245 19.555 -37.915 19.885 ;
        RECT -38.245 18.195 -37.915 18.525 ;
        RECT -38.245 16.835 -37.915 17.165 ;
        RECT -38.245 15.475 -37.915 15.805 ;
        RECT -38.245 14.115 -37.915 14.445 ;
        RECT -38.245 12.755 -37.915 13.085 ;
        RECT -38.245 11.395 -37.915 11.725 ;
        RECT -38.245 10.035 -37.915 10.365 ;
        RECT -38.245 8.675 -37.915 9.005 ;
        RECT -38.245 7.315 -37.915 7.645 ;
        RECT -38.245 5.955 -37.915 6.285 ;
        RECT -38.245 4.595 -37.915 4.925 ;
        RECT -38.245 3.235 -37.915 3.565 ;
        RECT -38.245 1.875 -37.915 2.205 ;
        RECT -38.245 0.515 -37.915 0.845 ;
        RECT -38.245 -0.845 -37.915 -0.515 ;
        RECT -38.245 -2.205 -37.915 -1.875 ;
        RECT -38.245 -3.565 -37.915 -3.235 ;
        RECT -38.245 -4.925 -37.915 -4.595 ;
        RECT -38.245 -6.285 -37.915 -5.955 ;
        RECT -38.245 -7.645 -37.915 -7.315 ;
        RECT -38.245 -9.005 -37.915 -8.675 ;
        RECT -38.245 -11.725 -37.915 -11.395 ;
        RECT -38.245 -13.085 -37.915 -12.755 ;
        RECT -38.245 -14.445 -37.915 -14.115 ;
        RECT -38.245 -15.805 -37.915 -15.475 ;
        RECT -38.245 -17.165 -37.915 -16.835 ;
        RECT -38.245 -18.525 -37.915 -18.195 ;
        RECT -38.245 -19.885 -37.915 -19.555 ;
        RECT -38.245 -26.685 -37.915 -26.355 ;
        RECT -38.245 -28.045 -37.915 -27.715 ;
        RECT -38.245 -29.405 -37.915 -29.075 ;
        RECT -38.245 -32.125 -37.915 -31.795 ;
        RECT -38.245 -34.845 -37.915 -34.515 ;
        RECT -38.245 -37.565 -37.915 -37.235 ;
        RECT -38.245 -38.925 -37.915 -38.595 ;
        RECT -38.245 -40.285 -37.915 -39.955 ;
        RECT -38.245 -41.645 -37.915 -41.315 ;
        RECT -38.245 -43.005 -37.915 -42.675 ;
        RECT -38.245 -44.365 -37.915 -44.035 ;
        RECT -38.245 -45.725 -37.915 -45.395 ;
        RECT -38.245 -47.085 -37.915 -46.755 ;
        RECT -38.245 -48.445 -37.915 -48.115 ;
        RECT -38.245 -49.805 -37.915 -49.475 ;
        RECT -38.245 -51.165 -37.915 -50.835 ;
        RECT -38.245 -52.525 -37.915 -52.195 ;
        RECT -38.245 -53.885 -37.915 -53.555 ;
        RECT -38.245 -55.245 -37.915 -54.915 ;
        RECT -38.245 -56.605 -37.915 -56.275 ;
        RECT -38.245 -57.965 -37.915 -57.635 ;
        RECT -38.245 -59.325 -37.915 -58.995 ;
        RECT -38.245 -60.685 -37.915 -60.355 ;
        RECT -38.245 -62.045 -37.915 -61.715 ;
        RECT -38.245 -63.405 -37.915 -63.075 ;
        RECT -38.245 -64.765 -37.915 -64.435 ;
        RECT -38.245 -66.125 -37.915 -65.795 ;
        RECT -38.245 -67.485 -37.915 -67.155 ;
        RECT -38.245 -68.845 -37.915 -68.515 ;
        RECT -38.245 -70.205 -37.915 -69.875 ;
        RECT -38.245 -71.565 -37.915 -71.235 ;
        RECT -38.245 -72.925 -37.915 -72.595 ;
        RECT -38.245 -74.285 -37.915 -73.955 ;
        RECT -38.245 -75.645 -37.915 -75.315 ;
        RECT -38.245 -77.005 -37.915 -76.675 ;
        RECT -38.245 -78.365 -37.915 -78.035 ;
        RECT -38.245 -79.725 -37.915 -79.395 ;
        RECT -38.245 -81.085 -37.915 -80.755 ;
        RECT -38.245 -82.445 -37.915 -82.115 ;
        RECT -38.245 -83.805 -37.915 -83.475 ;
        RECT -38.245 -85.165 -37.915 -84.835 ;
        RECT -38.245 -86.525 -37.915 -86.195 ;
        RECT -38.245 -87.885 -37.915 -87.555 ;
        RECT -38.245 -89.245 -37.915 -88.915 ;
        RECT -38.245 -90.605 -37.915 -90.275 ;
        RECT -38.245 -91.965 -37.915 -91.635 ;
        RECT -38.245 -93.325 -37.915 -92.995 ;
        RECT -38.245 -94.685 -37.915 -94.355 ;
        RECT -38.245 -96.045 -37.915 -95.715 ;
        RECT -38.245 -97.405 -37.915 -97.075 ;
        RECT -38.245 -98.765 -37.915 -98.435 ;
        RECT -38.245 -100.125 -37.915 -99.795 ;
        RECT -38.245 -101.485 -37.915 -101.155 ;
        RECT -38.245 -102.845 -37.915 -102.515 ;
        RECT -38.245 -104.205 -37.915 -103.875 ;
        RECT -38.245 -105.565 -37.915 -105.235 ;
        RECT -38.245 -106.925 -37.915 -106.595 ;
        RECT -38.245 -109.645 -37.915 -109.315 ;
        RECT -38.245 -111.005 -37.915 -110.675 ;
        RECT -38.245 -111.87 -37.915 -111.54 ;
        RECT -38.245 -113.725 -37.915 -113.395 ;
        RECT -38.245 -115.085 -37.915 -114.755 ;
        RECT -38.245 -116.445 -37.915 -116.115 ;
        RECT -38.245 -117.805 -37.915 -117.475 ;
        RECT -38.245 -120.525 -37.915 -120.195 ;
        RECT -38.245 -121.885 -37.915 -121.555 ;
        RECT -38.245 -123.245 -37.915 -122.915 ;
        RECT -38.245 -124.71 -37.915 -124.38 ;
        RECT -38.245 -125.965 -37.915 -125.635 ;
        RECT -38.245 -127.325 -37.915 -126.995 ;
        RECT -38.245 -130.045 -37.915 -129.715 ;
        RECT -38.245 -132.765 -37.915 -132.435 ;
        RECT -38.245 -134.125 -37.915 -133.795 ;
        RECT -38.245 -135.485 -37.915 -135.155 ;
        RECT -38.245 -136.845 -37.915 -136.515 ;
        RECT -38.245 -138.205 -37.915 -137.875 ;
        RECT -38.245 -139.565 -37.915 -139.235 ;
        RECT -38.245 -142.285 -37.915 -141.955 ;
        RECT -38.245 -143.645 -37.915 -143.315 ;
        RECT -38.245 -145.005 -37.915 -144.675 ;
        RECT -38.245 -146.365 -37.915 -146.035 ;
        RECT -38.245 -147.725 -37.915 -147.395 ;
        RECT -38.245 -149.085 -37.915 -148.755 ;
        RECT -38.245 -150.445 -37.915 -150.115 ;
        RECT -38.245 -151.805 -37.915 -151.475 ;
        RECT -38.245 -153.165 -37.915 -152.835 ;
        RECT -38.245 -154.525 -37.915 -154.195 ;
        RECT -38.245 -155.885 -37.915 -155.555 ;
        RECT -38.245 -157.245 -37.915 -156.915 ;
        RECT -38.245 -158.605 -37.915 -158.275 ;
        RECT -38.245 -159.965 -37.915 -159.635 ;
        RECT -38.245 -161.325 -37.915 -160.995 ;
        RECT -38.245 -162.685 -37.915 -162.355 ;
        RECT -38.245 -164.045 -37.915 -163.715 ;
        RECT -38.245 -165.405 -37.915 -165.075 ;
        RECT -38.245 -166.765 -37.915 -166.435 ;
        RECT -38.245 -168.125 -37.915 -167.795 ;
        RECT -38.245 -169.485 -37.915 -169.155 ;
        RECT -38.245 -170.845 -37.915 -170.515 ;
        RECT -38.245 -172.205 -37.915 -171.875 ;
        RECT -38.245 -173.565 -37.915 -173.235 ;
        RECT -38.245 -174.925 -37.915 -174.595 ;
        RECT -38.245 -176.285 -37.915 -175.955 ;
        RECT -38.245 -177.645 -37.915 -177.315 ;
        RECT -38.245 -179.005 -37.915 -178.675 ;
        RECT -38.245 -180.365 -37.915 -180.035 ;
        RECT -38.245 -181.725 -37.915 -181.395 ;
        RECT -38.245 -183.085 -37.915 -182.755 ;
        RECT -38.245 -184.445 -37.915 -184.115 ;
        RECT -38.245 -185.805 -37.915 -185.475 ;
        RECT -38.245 -187.165 -37.915 -186.835 ;
        RECT -38.245 -188.525 -37.915 -188.195 ;
        RECT -38.245 -189.885 -37.915 -189.555 ;
        RECT -38.245 -191.245 -37.915 -190.915 ;
        RECT -38.245 -192.605 -37.915 -192.275 ;
        RECT -38.245 -193.965 -37.915 -193.635 ;
        RECT -38.245 -195.325 -37.915 -194.995 ;
        RECT -38.245 -196.685 -37.915 -196.355 ;
        RECT -38.245 -198.045 -37.915 -197.715 ;
        RECT -38.245 -199.405 -37.915 -199.075 ;
        RECT -38.245 -200.765 -37.915 -200.435 ;
        RECT -38.245 -202.125 -37.915 -201.795 ;
        RECT -38.245 -203.485 -37.915 -203.155 ;
        RECT -38.245 -204.845 -37.915 -204.515 ;
        RECT -38.245 -206.555 -37.915 -206.225 ;
        RECT -38.245 -207.565 -37.915 -207.235 ;
        RECT -38.245 -208.925 -37.915 -208.595 ;
        RECT -38.245 -210.285 -37.915 -209.955 ;
        RECT -38.245 -211.645 -37.915 -211.315 ;
        RECT -38.245 -214.365 -37.915 -214.035 ;
        RECT -38.245 -215.725 -37.915 -215.395 ;
        RECT -38.245 -217.085 -37.915 -216.755 ;
        RECT -38.245 -218.445 -37.915 -218.115 ;
        RECT -38.245 -224.09 -37.915 -222.96 ;
        RECT -38.24 -224.205 -37.92 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.885 -134.125 -36.555 -133.795 ;
        RECT -36.885 -135.485 -36.555 -135.155 ;
        RECT -36.885 -136.845 -36.555 -136.515 ;
        RECT -36.885 -138.205 -36.555 -137.875 ;
        RECT -36.885 -139.565 -36.555 -139.235 ;
        RECT -36.885 -142.285 -36.555 -141.955 ;
        RECT -36.885 -143.645 -36.555 -143.315 ;
        RECT -36.885 -145.005 -36.555 -144.675 ;
        RECT -36.885 -146.365 -36.555 -146.035 ;
        RECT -36.885 -147.725 -36.555 -147.395 ;
        RECT -36.885 -149.085 -36.555 -148.755 ;
        RECT -36.885 -150.445 -36.555 -150.115 ;
        RECT -36.885 -151.805 -36.555 -151.475 ;
        RECT -36.885 -153.165 -36.555 -152.835 ;
        RECT -36.885 -154.525 -36.555 -154.195 ;
        RECT -36.885 -155.885 -36.555 -155.555 ;
        RECT -36.885 -157.245 -36.555 -156.915 ;
        RECT -36.885 -158.605 -36.555 -158.275 ;
        RECT -36.885 -159.965 -36.555 -159.635 ;
        RECT -36.885 -161.325 -36.555 -160.995 ;
        RECT -36.885 -162.685 -36.555 -162.355 ;
        RECT -36.885 -164.045 -36.555 -163.715 ;
        RECT -36.885 -165.405 -36.555 -165.075 ;
        RECT -36.885 -166.765 -36.555 -166.435 ;
        RECT -36.885 -168.125 -36.555 -167.795 ;
        RECT -36.885 -169.485 -36.555 -169.155 ;
        RECT -36.885 -170.845 -36.555 -170.515 ;
        RECT -36.885 -172.205 -36.555 -171.875 ;
        RECT -36.885 -173.565 -36.555 -173.235 ;
        RECT -36.885 -174.925 -36.555 -174.595 ;
        RECT -36.885 -176.285 -36.555 -175.955 ;
        RECT -36.885 -177.645 -36.555 -177.315 ;
        RECT -36.885 -179.005 -36.555 -178.675 ;
        RECT -36.885 -180.365 -36.555 -180.035 ;
        RECT -36.885 -181.725 -36.555 -181.395 ;
        RECT -36.885 -183.085 -36.555 -182.755 ;
        RECT -36.885 -184.445 -36.555 -184.115 ;
        RECT -36.885 -185.805 -36.555 -185.475 ;
        RECT -36.885 -187.165 -36.555 -186.835 ;
        RECT -36.885 -188.525 -36.555 -188.195 ;
        RECT -36.885 -189.885 -36.555 -189.555 ;
        RECT -36.885 -191.245 -36.555 -190.915 ;
        RECT -36.885 -192.605 -36.555 -192.275 ;
        RECT -36.885 -193.965 -36.555 -193.635 ;
        RECT -36.885 -195.325 -36.555 -194.995 ;
        RECT -36.885 -196.685 -36.555 -196.355 ;
        RECT -36.885 -198.045 -36.555 -197.715 ;
        RECT -36.885 -199.405 -36.555 -199.075 ;
        RECT -36.885 -200.765 -36.555 -200.435 ;
        RECT -36.885 -202.125 -36.555 -201.795 ;
        RECT -36.885 -203.485 -36.555 -203.155 ;
        RECT -36.885 -204.845 -36.555 -204.515 ;
        RECT -36.885 -206.555 -36.555 -206.225 ;
        RECT -36.885 -207.565 -36.555 -207.235 ;
        RECT -36.885 -208.925 -36.555 -208.595 ;
        RECT -36.885 -210.285 -36.555 -209.955 ;
        RECT -36.885 -211.645 -36.555 -211.315 ;
        RECT -36.885 -214.365 -36.555 -214.035 ;
        RECT -36.885 -215.725 -36.555 -215.395 ;
        RECT -36.885 -217.085 -36.555 -216.755 ;
        RECT -36.885 -218.445 -36.555 -218.115 ;
        RECT -36.885 -224.09 -36.555 -222.96 ;
        RECT -36.88 -224.205 -36.56 133.765 ;
        RECT -36.885 132.52 -36.555 133.65 ;
        RECT -36.885 128.355 -36.555 128.685 ;
        RECT -36.885 126.995 -36.555 127.325 ;
        RECT -36.885 125.635 -36.555 125.965 ;
        RECT -36.885 124.275 -36.555 124.605 ;
        RECT -36.885 122.915 -36.555 123.245 ;
        RECT -36.885 121.555 -36.555 121.885 ;
        RECT -36.885 120.195 -36.555 120.525 ;
        RECT -36.885 118.835 -36.555 119.165 ;
        RECT -36.885 117.475 -36.555 117.805 ;
        RECT -36.885 116.115 -36.555 116.445 ;
        RECT -36.885 114.755 -36.555 115.085 ;
        RECT -36.885 113.395 -36.555 113.725 ;
        RECT -36.885 112.035 -36.555 112.365 ;
        RECT -36.885 110.675 -36.555 111.005 ;
        RECT -36.885 109.315 -36.555 109.645 ;
        RECT -36.885 107.955 -36.555 108.285 ;
        RECT -36.885 106.595 -36.555 106.925 ;
        RECT -36.885 105.235 -36.555 105.565 ;
        RECT -36.885 103.875 -36.555 104.205 ;
        RECT -36.885 102.515 -36.555 102.845 ;
        RECT -36.885 101.155 -36.555 101.485 ;
        RECT -36.885 99.795 -36.555 100.125 ;
        RECT -36.885 98.435 -36.555 98.765 ;
        RECT -36.885 97.075 -36.555 97.405 ;
        RECT -36.885 95.715 -36.555 96.045 ;
        RECT -36.885 94.355 -36.555 94.685 ;
        RECT -36.885 92.995 -36.555 93.325 ;
        RECT -36.885 91.635 -36.555 91.965 ;
        RECT -36.885 90.275 -36.555 90.605 ;
        RECT -36.885 88.915 -36.555 89.245 ;
        RECT -36.885 87.555 -36.555 87.885 ;
        RECT -36.885 86.195 -36.555 86.525 ;
        RECT -36.885 84.835 -36.555 85.165 ;
        RECT -36.885 83.475 -36.555 83.805 ;
        RECT -36.885 82.115 -36.555 82.445 ;
        RECT -36.885 80.755 -36.555 81.085 ;
        RECT -36.885 79.395 -36.555 79.725 ;
        RECT -36.885 78.035 -36.555 78.365 ;
        RECT -36.885 76.675 -36.555 77.005 ;
        RECT -36.885 75.315 -36.555 75.645 ;
        RECT -36.885 73.955 -36.555 74.285 ;
        RECT -36.885 72.595 -36.555 72.925 ;
        RECT -36.885 71.235 -36.555 71.565 ;
        RECT -36.885 69.875 -36.555 70.205 ;
        RECT -36.885 68.515 -36.555 68.845 ;
        RECT -36.885 67.155 -36.555 67.485 ;
        RECT -36.885 65.795 -36.555 66.125 ;
        RECT -36.885 64.435 -36.555 64.765 ;
        RECT -36.885 63.075 -36.555 63.405 ;
        RECT -36.885 61.715 -36.555 62.045 ;
        RECT -36.885 60.355 -36.555 60.685 ;
        RECT -36.885 58.995 -36.555 59.325 ;
        RECT -36.885 57.635 -36.555 57.965 ;
        RECT -36.885 56.275 -36.555 56.605 ;
        RECT -36.885 54.915 -36.555 55.245 ;
        RECT -36.885 53.555 -36.555 53.885 ;
        RECT -36.885 52.195 -36.555 52.525 ;
        RECT -36.885 50.835 -36.555 51.165 ;
        RECT -36.885 49.475 -36.555 49.805 ;
        RECT -36.885 48.115 -36.555 48.445 ;
        RECT -36.885 46.755 -36.555 47.085 ;
        RECT -36.885 45.395 -36.555 45.725 ;
        RECT -36.885 44.035 -36.555 44.365 ;
        RECT -36.885 42.675 -36.555 43.005 ;
        RECT -36.885 41.315 -36.555 41.645 ;
        RECT -36.885 39.955 -36.555 40.285 ;
        RECT -36.885 38.595 -36.555 38.925 ;
        RECT -36.885 37.235 -36.555 37.565 ;
        RECT -36.885 35.875 -36.555 36.205 ;
        RECT -36.885 34.515 -36.555 34.845 ;
        RECT -36.885 33.155 -36.555 33.485 ;
        RECT -36.885 31.795 -36.555 32.125 ;
        RECT -36.885 30.435 -36.555 30.765 ;
        RECT -36.885 29.075 -36.555 29.405 ;
        RECT -36.885 27.715 -36.555 28.045 ;
        RECT -36.885 26.355 -36.555 26.685 ;
        RECT -36.885 24.995 -36.555 25.325 ;
        RECT -36.885 23.635 -36.555 23.965 ;
        RECT -36.885 22.275 -36.555 22.605 ;
        RECT -36.885 20.915 -36.555 21.245 ;
        RECT -36.885 19.555 -36.555 19.885 ;
        RECT -36.885 18.195 -36.555 18.525 ;
        RECT -36.885 16.835 -36.555 17.165 ;
        RECT -36.885 15.475 -36.555 15.805 ;
        RECT -36.885 14.115 -36.555 14.445 ;
        RECT -36.885 12.755 -36.555 13.085 ;
        RECT -36.885 11.395 -36.555 11.725 ;
        RECT -36.885 10.035 -36.555 10.365 ;
        RECT -36.885 8.675 -36.555 9.005 ;
        RECT -36.885 7.315 -36.555 7.645 ;
        RECT -36.885 5.955 -36.555 6.285 ;
        RECT -36.885 4.595 -36.555 4.925 ;
        RECT -36.885 3.235 -36.555 3.565 ;
        RECT -36.885 1.875 -36.555 2.205 ;
        RECT -36.885 0.515 -36.555 0.845 ;
        RECT -36.885 -0.845 -36.555 -0.515 ;
        RECT -36.885 -2.205 -36.555 -1.875 ;
        RECT -36.885 -3.565 -36.555 -3.235 ;
        RECT -36.885 -6.285 -36.555 -5.955 ;
        RECT -36.885 -7.645 -36.555 -7.315 ;
        RECT -36.885 -9.005 -36.555 -8.675 ;
        RECT -36.885 -11.725 -36.555 -11.395 ;
        RECT -36.885 -13.085 -36.555 -12.755 ;
        RECT -36.885 -14.445 -36.555 -14.115 ;
        RECT -36.885 -15.805 -36.555 -15.475 ;
        RECT -36.885 -17.165 -36.555 -16.835 ;
        RECT -36.885 -18.525 -36.555 -18.195 ;
        RECT -36.885 -19.885 -36.555 -19.555 ;
        RECT -36.885 -26.685 -36.555 -26.355 ;
        RECT -36.885 -28.045 -36.555 -27.715 ;
        RECT -36.885 -29.405 -36.555 -29.075 ;
        RECT -36.885 -32.125 -36.555 -31.795 ;
        RECT -36.885 -34.845 -36.555 -34.515 ;
        RECT -36.885 -37.565 -36.555 -37.235 ;
        RECT -36.885 -38.925 -36.555 -38.595 ;
        RECT -36.885 -40.285 -36.555 -39.955 ;
        RECT -36.885 -41.645 -36.555 -41.315 ;
        RECT -36.885 -43.005 -36.555 -42.675 ;
        RECT -36.885 -44.365 -36.555 -44.035 ;
        RECT -36.885 -45.725 -36.555 -45.395 ;
        RECT -36.885 -47.085 -36.555 -46.755 ;
        RECT -36.885 -48.445 -36.555 -48.115 ;
        RECT -36.885 -49.805 -36.555 -49.475 ;
        RECT -36.885 -51.165 -36.555 -50.835 ;
        RECT -36.885 -52.525 -36.555 -52.195 ;
        RECT -36.885 -53.885 -36.555 -53.555 ;
        RECT -36.885 -55.245 -36.555 -54.915 ;
        RECT -36.885 -56.605 -36.555 -56.275 ;
        RECT -36.885 -57.965 -36.555 -57.635 ;
        RECT -36.885 -59.325 -36.555 -58.995 ;
        RECT -36.885 -60.685 -36.555 -60.355 ;
        RECT -36.885 -62.045 -36.555 -61.715 ;
        RECT -36.885 -63.405 -36.555 -63.075 ;
        RECT -36.885 -64.765 -36.555 -64.435 ;
        RECT -36.885 -66.125 -36.555 -65.795 ;
        RECT -36.885 -67.485 -36.555 -67.155 ;
        RECT -36.885 -68.845 -36.555 -68.515 ;
        RECT -36.885 -70.205 -36.555 -69.875 ;
        RECT -36.885 -71.565 -36.555 -71.235 ;
        RECT -36.885 -72.925 -36.555 -72.595 ;
        RECT -36.885 -74.285 -36.555 -73.955 ;
        RECT -36.885 -75.645 -36.555 -75.315 ;
        RECT -36.885 -77.005 -36.555 -76.675 ;
        RECT -36.885 -78.365 -36.555 -78.035 ;
        RECT -36.885 -79.725 -36.555 -79.395 ;
        RECT -36.885 -81.085 -36.555 -80.755 ;
        RECT -36.885 -82.445 -36.555 -82.115 ;
        RECT -36.885 -83.805 -36.555 -83.475 ;
        RECT -36.885 -85.165 -36.555 -84.835 ;
        RECT -36.885 -86.525 -36.555 -86.195 ;
        RECT -36.885 -87.885 -36.555 -87.555 ;
        RECT -36.885 -89.245 -36.555 -88.915 ;
        RECT -36.885 -90.605 -36.555 -90.275 ;
        RECT -36.885 -91.965 -36.555 -91.635 ;
        RECT -36.885 -93.325 -36.555 -92.995 ;
        RECT -36.885 -94.685 -36.555 -94.355 ;
        RECT -36.885 -96.045 -36.555 -95.715 ;
        RECT -36.885 -97.405 -36.555 -97.075 ;
        RECT -36.885 -98.765 -36.555 -98.435 ;
        RECT -36.885 -100.125 -36.555 -99.795 ;
        RECT -36.885 -101.485 -36.555 -101.155 ;
        RECT -36.885 -102.845 -36.555 -102.515 ;
        RECT -36.885 -104.205 -36.555 -103.875 ;
        RECT -36.885 -105.565 -36.555 -105.235 ;
        RECT -36.885 -106.925 -36.555 -106.595 ;
        RECT -36.885 -109.645 -36.555 -109.315 ;
        RECT -36.885 -111.005 -36.555 -110.675 ;
        RECT -36.885 -111.87 -36.555 -111.54 ;
        RECT -36.885 -113.725 -36.555 -113.395 ;
        RECT -36.885 -115.085 -36.555 -114.755 ;
        RECT -36.885 -116.445 -36.555 -116.115 ;
        RECT -36.885 -117.805 -36.555 -117.475 ;
        RECT -36.885 -120.525 -36.555 -120.195 ;
        RECT -36.885 -121.885 -36.555 -121.555 ;
        RECT -36.885 -123.245 -36.555 -122.915 ;
        RECT -36.885 -124.71 -36.555 -124.38 ;
        RECT -36.885 -125.965 -36.555 -125.635 ;
        RECT -36.885 -127.325 -36.555 -126.995 ;
        RECT -36.885 -130.045 -36.555 -129.715 ;
        RECT -36.885 -132.765 -36.555 -132.435 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.765 132.52 -47.435 133.65 ;
        RECT -47.765 128.355 -47.435 128.685 ;
        RECT -47.765 126.995 -47.435 127.325 ;
        RECT -47.765 125.635 -47.435 125.965 ;
        RECT -47.765 124.275 -47.435 124.605 ;
        RECT -47.765 122.915 -47.435 123.245 ;
        RECT -47.765 121.555 -47.435 121.885 ;
        RECT -47.765 120.195 -47.435 120.525 ;
        RECT -47.765 118.835 -47.435 119.165 ;
        RECT -47.765 117.475 -47.435 117.805 ;
        RECT -47.765 116.115 -47.435 116.445 ;
        RECT -47.765 114.755 -47.435 115.085 ;
        RECT -47.765 113.395 -47.435 113.725 ;
        RECT -47.765 112.035 -47.435 112.365 ;
        RECT -47.765 110.675 -47.435 111.005 ;
        RECT -47.765 109.315 -47.435 109.645 ;
        RECT -47.765 107.955 -47.435 108.285 ;
        RECT -47.765 106.595 -47.435 106.925 ;
        RECT -47.765 105.235 -47.435 105.565 ;
        RECT -47.765 103.875 -47.435 104.205 ;
        RECT -47.765 102.515 -47.435 102.845 ;
        RECT -47.765 101.155 -47.435 101.485 ;
        RECT -47.765 99.795 -47.435 100.125 ;
        RECT -47.765 98.435 -47.435 98.765 ;
        RECT -47.765 97.075 -47.435 97.405 ;
        RECT -47.765 95.715 -47.435 96.045 ;
        RECT -47.765 94.355 -47.435 94.685 ;
        RECT -47.765 92.995 -47.435 93.325 ;
        RECT -47.765 91.635 -47.435 91.965 ;
        RECT -47.765 90.275 -47.435 90.605 ;
        RECT -47.765 88.915 -47.435 89.245 ;
        RECT -47.765 87.555 -47.435 87.885 ;
        RECT -47.765 86.195 -47.435 86.525 ;
        RECT -47.765 84.835 -47.435 85.165 ;
        RECT -47.765 83.475 -47.435 83.805 ;
        RECT -47.765 82.115 -47.435 82.445 ;
        RECT -47.765 80.755 -47.435 81.085 ;
        RECT -47.765 79.395 -47.435 79.725 ;
        RECT -47.765 78.035 -47.435 78.365 ;
        RECT -47.765 76.675 -47.435 77.005 ;
        RECT -47.765 75.315 -47.435 75.645 ;
        RECT -47.765 73.955 -47.435 74.285 ;
        RECT -47.76 73.28 -47.44 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.765 48.115 -47.435 48.445 ;
        RECT -47.765 46.755 -47.435 47.085 ;
        RECT -47.765 45.395 -47.435 45.725 ;
        RECT -47.765 44.035 -47.435 44.365 ;
        RECT -47.765 39.955 -47.435 40.285 ;
        RECT -47.765 38.595 -47.435 38.925 ;
        RECT -47.765 35.875 -47.435 36.205 ;
        RECT -47.765 34.515 -47.435 34.845 ;
        RECT -47.765 33.155 -47.435 33.485 ;
        RECT -47.765 31.795 -47.435 32.125 ;
        RECT -47.765 30.435 -47.435 30.765 ;
        RECT -47.765 29.075 -47.435 29.405 ;
        RECT -47.765 27.715 -47.435 28.045 ;
        RECT -47.765 26.355 -47.435 26.685 ;
        RECT -47.765 24.995 -47.435 25.325 ;
        RECT -47.765 23.635 -47.435 23.965 ;
        RECT -47.765 22.275 -47.435 22.605 ;
        RECT -47.765 20.915 -47.435 21.245 ;
        RECT -47.765 19.555 -47.435 19.885 ;
        RECT -47.765 18.195 -47.435 18.525 ;
        RECT -47.765 16.835 -47.435 17.165 ;
        RECT -47.765 15.475 -47.435 15.805 ;
        RECT -47.765 14.115 -47.435 14.445 ;
        RECT -47.765 12.755 -47.435 13.085 ;
        RECT -47.765 11.395 -47.435 11.725 ;
        RECT -47.765 10.035 -47.435 10.365 ;
        RECT -47.765 8.675 -47.435 9.005 ;
        RECT -47.765 7.315 -47.435 7.645 ;
        RECT -47.765 5.955 -47.435 6.285 ;
        RECT -47.765 4.595 -47.435 4.925 ;
        RECT -47.765 3.235 -47.435 3.565 ;
        RECT -47.765 1.875 -47.435 2.205 ;
        RECT -47.765 0.515 -47.435 0.845 ;
        RECT -47.765 -0.845 -47.435 -0.515 ;
        RECT -47.765 -2.205 -47.435 -1.875 ;
        RECT -47.765 -3.565 -47.435 -3.235 ;
        RECT -47.765 -4.925 -47.435 -4.595 ;
        RECT -47.765 -6.285 -47.435 -5.955 ;
        RECT -47.765 -7.645 -47.435 -7.315 ;
        RECT -47.765 -9.005 -47.435 -8.675 ;
        RECT -47.765 -11.725 -47.435 -11.395 ;
        RECT -47.765 -13.085 -47.435 -12.755 ;
        RECT -47.765 -14.445 -47.435 -14.115 ;
        RECT -47.765 -15.805 -47.435 -15.475 ;
        RECT -47.765 -17.165 -47.435 -16.835 ;
        RECT -47.765 -18.525 -47.435 -18.195 ;
        RECT -47.765 -19.885 -47.435 -19.555 ;
        RECT -47.765 -21.245 -47.435 -20.915 ;
        RECT -47.765 -22.605 -47.435 -22.275 ;
        RECT -47.765 -23.965 -47.435 -23.635 ;
        RECT -47.765 -25.325 -47.435 -24.995 ;
        RECT -47.765 -26.685 -47.435 -26.355 ;
        RECT -47.765 -28.045 -47.435 -27.715 ;
        RECT -47.765 -29.405 -47.435 -29.075 ;
        RECT -47.765 -30.765 -47.435 -30.435 ;
        RECT -47.765 -32.125 -47.435 -31.795 ;
        RECT -47.765 -34.845 -47.435 -34.515 ;
        RECT -47.765 -37.565 -47.435 -37.235 ;
        RECT -47.765 -38.925 -47.435 -38.595 ;
        RECT -47.765 -40.285 -47.435 -39.955 ;
        RECT -47.765 -41.645 -47.435 -41.315 ;
        RECT -47.765 -43.005 -47.435 -42.675 ;
        RECT -47.765 -44.365 -47.435 -44.035 ;
        RECT -47.765 -45.725 -47.435 -45.395 ;
        RECT -47.765 -47.085 -47.435 -46.755 ;
        RECT -47.765 -48.445 -47.435 -48.115 ;
        RECT -47.765 -49.805 -47.435 -49.475 ;
        RECT -47.765 -51.165 -47.435 -50.835 ;
        RECT -47.765 -52.525 -47.435 -52.195 ;
        RECT -47.765 -53.885 -47.435 -53.555 ;
        RECT -47.765 -55.245 -47.435 -54.915 ;
        RECT -47.765 -56.605 -47.435 -56.275 ;
        RECT -47.765 -57.965 -47.435 -57.635 ;
        RECT -47.765 -59.325 -47.435 -58.995 ;
        RECT -47.765 -60.685 -47.435 -60.355 ;
        RECT -47.765 -62.045 -47.435 -61.715 ;
        RECT -47.765 -63.405 -47.435 -63.075 ;
        RECT -47.765 -64.765 -47.435 -64.435 ;
        RECT -47.765 -66.125 -47.435 -65.795 ;
        RECT -47.765 -67.485 -47.435 -67.155 ;
        RECT -47.765 -68.845 -47.435 -68.515 ;
        RECT -47.765 -70.205 -47.435 -69.875 ;
        RECT -47.765 -71.565 -47.435 -71.235 ;
        RECT -47.765 -72.925 -47.435 -72.595 ;
        RECT -47.765 -74.285 -47.435 -73.955 ;
        RECT -47.765 -75.645 -47.435 -75.315 ;
        RECT -47.765 -77.005 -47.435 -76.675 ;
        RECT -47.765 -78.365 -47.435 -78.035 ;
        RECT -47.765 -79.725 -47.435 -79.395 ;
        RECT -47.765 -81.085 -47.435 -80.755 ;
        RECT -47.765 -82.445 -47.435 -82.115 ;
        RECT -47.765 -83.805 -47.435 -83.475 ;
        RECT -47.765 -85.165 -47.435 -84.835 ;
        RECT -47.765 -86.525 -47.435 -86.195 ;
        RECT -47.765 -87.885 -47.435 -87.555 ;
        RECT -47.765 -89.245 -47.435 -88.915 ;
        RECT -47.765 -90.605 -47.435 -90.275 ;
        RECT -47.765 -91.965 -47.435 -91.635 ;
        RECT -47.765 -93.325 -47.435 -92.995 ;
        RECT -47.765 -94.685 -47.435 -94.355 ;
        RECT -47.765 -96.045 -47.435 -95.715 ;
        RECT -47.765 -97.405 -47.435 -97.075 ;
        RECT -47.765 -98.765 -47.435 -98.435 ;
        RECT -47.765 -100.125 -47.435 -99.795 ;
        RECT -47.765 -101.485 -47.435 -101.155 ;
        RECT -47.765 -102.845 -47.435 -102.515 ;
        RECT -47.765 -104.205 -47.435 -103.875 ;
        RECT -47.765 -105.565 -47.435 -105.235 ;
        RECT -47.765 -106.925 -47.435 -106.595 ;
        RECT -47.765 -108.285 -47.435 -107.955 ;
        RECT -47.765 -109.645 -47.435 -109.315 ;
        RECT -47.765 -111.005 -47.435 -110.675 ;
        RECT -47.765 -111.87 -47.435 -111.54 ;
        RECT -47.765 -113.725 -47.435 -113.395 ;
        RECT -47.765 -115.085 -47.435 -114.755 ;
        RECT -47.765 -116.445 -47.435 -116.115 ;
        RECT -47.765 -117.805 -47.435 -117.475 ;
        RECT -47.765 -120.525 -47.435 -120.195 ;
        RECT -47.765 -121.885 -47.435 -121.555 ;
        RECT -47.765 -123.245 -47.435 -122.915 ;
        RECT -47.765 -124.71 -47.435 -124.38 ;
        RECT -47.765 -125.965 -47.435 -125.635 ;
        RECT -47.765 -127.325 -47.435 -126.995 ;
        RECT -47.765 -130.045 -47.435 -129.715 ;
        RECT -47.765 -132.765 -47.435 -132.435 ;
        RECT -47.765 -134.125 -47.435 -133.795 ;
        RECT -47.765 -135.485 -47.435 -135.155 ;
        RECT -47.765 -136.845 -47.435 -136.515 ;
        RECT -47.765 -138.205 -47.435 -137.875 ;
        RECT -47.765 -139.565 -47.435 -139.235 ;
        RECT -47.765 -142.285 -47.435 -141.955 ;
        RECT -47.765 -143.645 -47.435 -143.315 ;
        RECT -47.765 -145.005 -47.435 -144.675 ;
        RECT -47.765 -146.365 -47.435 -146.035 ;
        RECT -47.765 -147.725 -47.435 -147.395 ;
        RECT -47.765 -149.085 -47.435 -148.755 ;
        RECT -47.765 -150.445 -47.435 -150.115 ;
        RECT -47.765 -151.805 -47.435 -151.475 ;
        RECT -47.765 -153.165 -47.435 -152.835 ;
        RECT -47.765 -154.525 -47.435 -154.195 ;
        RECT -47.765 -155.885 -47.435 -155.555 ;
        RECT -47.765 -157.245 -47.435 -156.915 ;
        RECT -47.765 -158.605 -47.435 -158.275 ;
        RECT -47.765 -159.965 -47.435 -159.635 ;
        RECT -47.765 -161.325 -47.435 -160.995 ;
        RECT -47.765 -162.685 -47.435 -162.355 ;
        RECT -47.765 -164.045 -47.435 -163.715 ;
        RECT -47.765 -165.405 -47.435 -165.075 ;
        RECT -47.765 -166.765 -47.435 -166.435 ;
        RECT -47.765 -168.125 -47.435 -167.795 ;
        RECT -47.765 -169.485 -47.435 -169.155 ;
        RECT -47.765 -170.845 -47.435 -170.515 ;
        RECT -47.765 -172.205 -47.435 -171.875 ;
        RECT -47.765 -173.565 -47.435 -173.235 ;
        RECT -47.765 -174.925 -47.435 -174.595 ;
        RECT -47.765 -176.285 -47.435 -175.955 ;
        RECT -47.765 -177.645 -47.435 -177.315 ;
        RECT -47.765 -179.005 -47.435 -178.675 ;
        RECT -47.765 -180.365 -47.435 -180.035 ;
        RECT -47.765 -181.725 -47.435 -181.395 ;
        RECT -47.765 -183.085 -47.435 -182.755 ;
        RECT -47.765 -184.445 -47.435 -184.115 ;
        RECT -47.765 -185.805 -47.435 -185.475 ;
        RECT -47.765 -187.165 -47.435 -186.835 ;
        RECT -47.765 -188.525 -47.435 -188.195 ;
        RECT -47.765 -189.885 -47.435 -189.555 ;
        RECT -47.765 -191.245 -47.435 -190.915 ;
        RECT -47.765 -192.605 -47.435 -192.275 ;
        RECT -47.765 -193.965 -47.435 -193.635 ;
        RECT -47.765 -195.325 -47.435 -194.995 ;
        RECT -47.765 -196.685 -47.435 -196.355 ;
        RECT -47.765 -198.045 -47.435 -197.715 ;
        RECT -47.765 -199.405 -47.435 -199.075 ;
        RECT -47.765 -200.765 -47.435 -200.435 ;
        RECT -47.765 -202.125 -47.435 -201.795 ;
        RECT -47.765 -203.485 -47.435 -203.155 ;
        RECT -47.765 -204.845 -47.435 -204.515 ;
        RECT -47.765 -206.555 -47.435 -206.225 ;
        RECT -47.765 -207.565 -47.435 -207.235 ;
        RECT -47.765 -208.925 -47.435 -208.595 ;
        RECT -47.765 -214.365 -47.435 -214.035 ;
        RECT -47.765 -215.725 -47.435 -215.395 ;
        RECT -47.765 -217.085 -47.435 -216.755 ;
        RECT -47.765 -218.445 -47.435 -218.115 ;
        RECT -47.765 -224.09 -47.435 -222.96 ;
        RECT -47.76 -224.205 -47.44 49.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -46.405 132.52 -46.075 133.65 ;
        RECT -46.405 128.355 -46.075 128.685 ;
        RECT -46.405 126.995 -46.075 127.325 ;
        RECT -46.405 125.635 -46.075 125.965 ;
        RECT -46.405 124.275 -46.075 124.605 ;
        RECT -46.405 122.915 -46.075 123.245 ;
        RECT -46.405 121.555 -46.075 121.885 ;
        RECT -46.405 120.195 -46.075 120.525 ;
        RECT -46.405 118.835 -46.075 119.165 ;
        RECT -46.405 117.475 -46.075 117.805 ;
        RECT -46.405 116.115 -46.075 116.445 ;
        RECT -46.405 114.755 -46.075 115.085 ;
        RECT -46.405 113.395 -46.075 113.725 ;
        RECT -46.405 112.035 -46.075 112.365 ;
        RECT -46.405 110.675 -46.075 111.005 ;
        RECT -46.405 109.315 -46.075 109.645 ;
        RECT -46.405 107.955 -46.075 108.285 ;
        RECT -46.405 106.595 -46.075 106.925 ;
        RECT -46.405 105.235 -46.075 105.565 ;
        RECT -46.405 103.875 -46.075 104.205 ;
        RECT -46.405 102.515 -46.075 102.845 ;
        RECT -46.405 101.155 -46.075 101.485 ;
        RECT -46.405 99.795 -46.075 100.125 ;
        RECT -46.405 98.435 -46.075 98.765 ;
        RECT -46.405 97.075 -46.075 97.405 ;
        RECT -46.405 95.715 -46.075 96.045 ;
        RECT -46.405 94.355 -46.075 94.685 ;
        RECT -46.405 92.995 -46.075 93.325 ;
        RECT -46.405 91.635 -46.075 91.965 ;
        RECT -46.405 90.275 -46.075 90.605 ;
        RECT -46.405 88.915 -46.075 89.245 ;
        RECT -46.405 87.555 -46.075 87.885 ;
        RECT -46.405 86.195 -46.075 86.525 ;
        RECT -46.405 84.835 -46.075 85.165 ;
        RECT -46.405 83.475 -46.075 83.805 ;
        RECT -46.405 82.115 -46.075 82.445 ;
        RECT -46.405 80.755 -46.075 81.085 ;
        RECT -46.405 79.395 -46.075 79.725 ;
        RECT -46.405 78.035 -46.075 78.365 ;
        RECT -46.405 76.675 -46.075 77.005 ;
        RECT -46.405 75.315 -46.075 75.645 ;
        RECT -46.405 73.955 -46.075 74.285 ;
        RECT -46.4 73.28 -46.08 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -46.405 48.115 -46.075 48.445 ;
        RECT -46.405 46.755 -46.075 47.085 ;
        RECT -46.405 45.395 -46.075 45.725 ;
        RECT -46.405 44.035 -46.075 44.365 ;
        RECT -46.405 39.955 -46.075 40.285 ;
        RECT -46.405 38.595 -46.075 38.925 ;
        RECT -46.405 35.875 -46.075 36.205 ;
        RECT -46.405 34.515 -46.075 34.845 ;
        RECT -46.405 33.155 -46.075 33.485 ;
        RECT -46.405 31.795 -46.075 32.125 ;
        RECT -46.405 30.435 -46.075 30.765 ;
        RECT -46.405 29.075 -46.075 29.405 ;
        RECT -46.405 27.715 -46.075 28.045 ;
        RECT -46.405 26.355 -46.075 26.685 ;
        RECT -46.405 24.995 -46.075 25.325 ;
        RECT -46.405 23.635 -46.075 23.965 ;
        RECT -46.405 22.275 -46.075 22.605 ;
        RECT -46.405 20.915 -46.075 21.245 ;
        RECT -46.405 19.555 -46.075 19.885 ;
        RECT -46.405 18.195 -46.075 18.525 ;
        RECT -46.405 16.835 -46.075 17.165 ;
        RECT -46.405 15.475 -46.075 15.805 ;
        RECT -46.405 14.115 -46.075 14.445 ;
        RECT -46.405 12.755 -46.075 13.085 ;
        RECT -46.405 11.395 -46.075 11.725 ;
        RECT -46.405 10.035 -46.075 10.365 ;
        RECT -46.405 8.675 -46.075 9.005 ;
        RECT -46.405 7.315 -46.075 7.645 ;
        RECT -46.405 5.955 -46.075 6.285 ;
        RECT -46.405 4.595 -46.075 4.925 ;
        RECT -46.405 3.235 -46.075 3.565 ;
        RECT -46.405 1.875 -46.075 2.205 ;
        RECT -46.405 0.515 -46.075 0.845 ;
        RECT -46.405 -0.845 -46.075 -0.515 ;
        RECT -46.405 -2.205 -46.075 -1.875 ;
        RECT -46.405 -3.565 -46.075 -3.235 ;
        RECT -46.405 -4.925 -46.075 -4.595 ;
        RECT -46.405 -6.285 -46.075 -5.955 ;
        RECT -46.405 -7.645 -46.075 -7.315 ;
        RECT -46.405 -9.005 -46.075 -8.675 ;
        RECT -46.405 -11.725 -46.075 -11.395 ;
        RECT -46.405 -13.085 -46.075 -12.755 ;
        RECT -46.405 -14.445 -46.075 -14.115 ;
        RECT -46.405 -15.805 -46.075 -15.475 ;
        RECT -46.405 -17.165 -46.075 -16.835 ;
        RECT -46.405 -18.525 -46.075 -18.195 ;
        RECT -46.405 -19.885 -46.075 -19.555 ;
        RECT -46.405 -21.245 -46.075 -20.915 ;
        RECT -46.405 -22.605 -46.075 -22.275 ;
        RECT -46.405 -23.965 -46.075 -23.635 ;
        RECT -46.405 -25.325 -46.075 -24.995 ;
        RECT -46.405 -26.685 -46.075 -26.355 ;
        RECT -46.405 -28.045 -46.075 -27.715 ;
        RECT -46.405 -29.405 -46.075 -29.075 ;
        RECT -46.405 -30.765 -46.075 -30.435 ;
        RECT -46.405 -32.125 -46.075 -31.795 ;
        RECT -46.405 -34.845 -46.075 -34.515 ;
        RECT -46.405 -37.565 -46.075 -37.235 ;
        RECT -46.405 -38.925 -46.075 -38.595 ;
        RECT -46.405 -40.285 -46.075 -39.955 ;
        RECT -46.405 -41.645 -46.075 -41.315 ;
        RECT -46.405 -43.005 -46.075 -42.675 ;
        RECT -46.405 -44.365 -46.075 -44.035 ;
        RECT -46.405 -45.725 -46.075 -45.395 ;
        RECT -46.405 -47.085 -46.075 -46.755 ;
        RECT -46.405 -48.445 -46.075 -48.115 ;
        RECT -46.405 -49.805 -46.075 -49.475 ;
        RECT -46.405 -51.165 -46.075 -50.835 ;
        RECT -46.405 -52.525 -46.075 -52.195 ;
        RECT -46.405 -53.885 -46.075 -53.555 ;
        RECT -46.405 -55.245 -46.075 -54.915 ;
        RECT -46.405 -56.605 -46.075 -56.275 ;
        RECT -46.405 -57.965 -46.075 -57.635 ;
        RECT -46.405 -59.325 -46.075 -58.995 ;
        RECT -46.405 -60.685 -46.075 -60.355 ;
        RECT -46.405 -62.045 -46.075 -61.715 ;
        RECT -46.405 -63.405 -46.075 -63.075 ;
        RECT -46.405 -64.765 -46.075 -64.435 ;
        RECT -46.405 -66.125 -46.075 -65.795 ;
        RECT -46.405 -67.485 -46.075 -67.155 ;
        RECT -46.405 -68.845 -46.075 -68.515 ;
        RECT -46.405 -70.205 -46.075 -69.875 ;
        RECT -46.405 -71.565 -46.075 -71.235 ;
        RECT -46.405 -72.925 -46.075 -72.595 ;
        RECT -46.405 -74.285 -46.075 -73.955 ;
        RECT -46.405 -75.645 -46.075 -75.315 ;
        RECT -46.405 -77.005 -46.075 -76.675 ;
        RECT -46.405 -78.365 -46.075 -78.035 ;
        RECT -46.405 -79.725 -46.075 -79.395 ;
        RECT -46.405 -81.085 -46.075 -80.755 ;
        RECT -46.405 -82.445 -46.075 -82.115 ;
        RECT -46.405 -83.805 -46.075 -83.475 ;
        RECT -46.405 -85.165 -46.075 -84.835 ;
        RECT -46.405 -86.525 -46.075 -86.195 ;
        RECT -46.405 -87.885 -46.075 -87.555 ;
        RECT -46.405 -89.245 -46.075 -88.915 ;
        RECT -46.405 -90.605 -46.075 -90.275 ;
        RECT -46.405 -91.965 -46.075 -91.635 ;
        RECT -46.405 -93.325 -46.075 -92.995 ;
        RECT -46.405 -94.685 -46.075 -94.355 ;
        RECT -46.405 -96.045 -46.075 -95.715 ;
        RECT -46.405 -97.405 -46.075 -97.075 ;
        RECT -46.405 -98.765 -46.075 -98.435 ;
        RECT -46.405 -100.125 -46.075 -99.795 ;
        RECT -46.405 -101.485 -46.075 -101.155 ;
        RECT -46.405 -102.845 -46.075 -102.515 ;
        RECT -46.405 -104.205 -46.075 -103.875 ;
        RECT -46.405 -105.565 -46.075 -105.235 ;
        RECT -46.405 -106.925 -46.075 -106.595 ;
        RECT -46.405 -108.285 -46.075 -107.955 ;
        RECT -46.405 -109.645 -46.075 -109.315 ;
        RECT -46.405 -111.005 -46.075 -110.675 ;
        RECT -46.405 -111.87 -46.075 -111.54 ;
        RECT -46.405 -113.725 -46.075 -113.395 ;
        RECT -46.405 -115.085 -46.075 -114.755 ;
        RECT -46.405 -116.445 -46.075 -116.115 ;
        RECT -46.405 -117.805 -46.075 -117.475 ;
        RECT -46.405 -120.525 -46.075 -120.195 ;
        RECT -46.405 -121.885 -46.075 -121.555 ;
        RECT -46.405 -123.245 -46.075 -122.915 ;
        RECT -46.405 -124.71 -46.075 -124.38 ;
        RECT -46.405 -125.965 -46.075 -125.635 ;
        RECT -46.405 -127.325 -46.075 -126.995 ;
        RECT -46.405 -130.045 -46.075 -129.715 ;
        RECT -46.405 -134.125 -46.075 -133.795 ;
        RECT -46.405 -135.485 -46.075 -135.155 ;
        RECT -46.405 -136.845 -46.075 -136.515 ;
        RECT -46.405 -138.205 -46.075 -137.875 ;
        RECT -46.405 -139.565 -46.075 -139.235 ;
        RECT -46.405 -142.285 -46.075 -141.955 ;
        RECT -46.405 -143.645 -46.075 -143.315 ;
        RECT -46.405 -145.005 -46.075 -144.675 ;
        RECT -46.405 -146.365 -46.075 -146.035 ;
        RECT -46.405 -147.725 -46.075 -147.395 ;
        RECT -46.405 -149.085 -46.075 -148.755 ;
        RECT -46.405 -150.445 -46.075 -150.115 ;
        RECT -46.405 -151.805 -46.075 -151.475 ;
        RECT -46.405 -153.165 -46.075 -152.835 ;
        RECT -46.405 -154.525 -46.075 -154.195 ;
        RECT -46.405 -155.885 -46.075 -155.555 ;
        RECT -46.405 -157.245 -46.075 -156.915 ;
        RECT -46.405 -158.605 -46.075 -158.275 ;
        RECT -46.405 -159.965 -46.075 -159.635 ;
        RECT -46.405 -161.325 -46.075 -160.995 ;
        RECT -46.405 -162.685 -46.075 -162.355 ;
        RECT -46.405 -164.045 -46.075 -163.715 ;
        RECT -46.405 -165.405 -46.075 -165.075 ;
        RECT -46.405 -166.765 -46.075 -166.435 ;
        RECT -46.405 -168.125 -46.075 -167.795 ;
        RECT -46.405 -169.485 -46.075 -169.155 ;
        RECT -46.405 -170.845 -46.075 -170.515 ;
        RECT -46.405 -172.205 -46.075 -171.875 ;
        RECT -46.405 -173.565 -46.075 -173.235 ;
        RECT -46.405 -174.925 -46.075 -174.595 ;
        RECT -46.405 -176.285 -46.075 -175.955 ;
        RECT -46.405 -177.645 -46.075 -177.315 ;
        RECT -46.405 -179.005 -46.075 -178.675 ;
        RECT -46.405 -180.365 -46.075 -180.035 ;
        RECT -46.405 -181.725 -46.075 -181.395 ;
        RECT -46.405 -183.085 -46.075 -182.755 ;
        RECT -46.405 -184.445 -46.075 -184.115 ;
        RECT -46.405 -185.805 -46.075 -185.475 ;
        RECT -46.405 -187.165 -46.075 -186.835 ;
        RECT -46.405 -188.525 -46.075 -188.195 ;
        RECT -46.405 -189.885 -46.075 -189.555 ;
        RECT -46.405 -191.245 -46.075 -190.915 ;
        RECT -46.405 -192.605 -46.075 -192.275 ;
        RECT -46.405 -193.965 -46.075 -193.635 ;
        RECT -46.405 -195.325 -46.075 -194.995 ;
        RECT -46.405 -196.685 -46.075 -196.355 ;
        RECT -46.405 -198.045 -46.075 -197.715 ;
        RECT -46.405 -199.405 -46.075 -199.075 ;
        RECT -46.405 -200.765 -46.075 -200.435 ;
        RECT -46.405 -202.125 -46.075 -201.795 ;
        RECT -46.405 -203.485 -46.075 -203.155 ;
        RECT -46.405 -204.845 -46.075 -204.515 ;
        RECT -46.405 -206.555 -46.075 -206.225 ;
        RECT -46.405 -207.565 -46.075 -207.235 ;
        RECT -46.405 -208.925 -46.075 -208.595 ;
        RECT -46.4 -209.6 -46.08 49.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.045 132.52 -44.715 133.65 ;
        RECT -45.045 128.355 -44.715 128.685 ;
        RECT -45.045 126.995 -44.715 127.325 ;
        RECT -45.045 125.635 -44.715 125.965 ;
        RECT -45.045 124.275 -44.715 124.605 ;
        RECT -45.045 122.915 -44.715 123.245 ;
        RECT -45.045 121.555 -44.715 121.885 ;
        RECT -45.045 120.195 -44.715 120.525 ;
        RECT -45.045 118.835 -44.715 119.165 ;
        RECT -45.045 117.475 -44.715 117.805 ;
        RECT -45.045 116.115 -44.715 116.445 ;
        RECT -45.045 114.755 -44.715 115.085 ;
        RECT -45.045 113.395 -44.715 113.725 ;
        RECT -45.045 112.035 -44.715 112.365 ;
        RECT -45.045 110.675 -44.715 111.005 ;
        RECT -45.045 109.315 -44.715 109.645 ;
        RECT -45.045 107.955 -44.715 108.285 ;
        RECT -45.045 106.595 -44.715 106.925 ;
        RECT -45.045 105.235 -44.715 105.565 ;
        RECT -45.045 103.875 -44.715 104.205 ;
        RECT -45.045 102.515 -44.715 102.845 ;
        RECT -45.045 101.155 -44.715 101.485 ;
        RECT -45.045 99.795 -44.715 100.125 ;
        RECT -45.045 98.435 -44.715 98.765 ;
        RECT -45.045 97.075 -44.715 97.405 ;
        RECT -45.045 95.715 -44.715 96.045 ;
        RECT -45.045 94.355 -44.715 94.685 ;
        RECT -45.045 92.995 -44.715 93.325 ;
        RECT -45.045 91.635 -44.715 91.965 ;
        RECT -45.045 90.275 -44.715 90.605 ;
        RECT -45.045 88.915 -44.715 89.245 ;
        RECT -45.045 87.555 -44.715 87.885 ;
        RECT -45.045 86.195 -44.715 86.525 ;
        RECT -45.045 84.835 -44.715 85.165 ;
        RECT -45.045 83.475 -44.715 83.805 ;
        RECT -45.045 82.115 -44.715 82.445 ;
        RECT -45.045 80.755 -44.715 81.085 ;
        RECT -45.045 79.395 -44.715 79.725 ;
        RECT -45.045 78.035 -44.715 78.365 ;
        RECT -45.045 76.675 -44.715 77.005 ;
        RECT -45.045 75.315 -44.715 75.645 ;
        RECT -45.045 73.955 -44.715 74.285 ;
        RECT -45.045 71.64 -44.715 71.97 ;
        RECT -45.045 69.465 -44.715 69.795 ;
        RECT -45.045 68.615 -44.715 68.945 ;
        RECT -45.045 66.305 -44.715 66.635 ;
        RECT -45.045 65.455 -44.715 65.785 ;
        RECT -45.045 63.145 -44.715 63.475 ;
        RECT -45.04 62.4 -44.72 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.045 -139.565 -44.715 -139.235 ;
        RECT -45.045 -142.285 -44.715 -141.955 ;
        RECT -45.045 -143.645 -44.715 -143.315 ;
        RECT -45.045 -145.005 -44.715 -144.675 ;
        RECT -45.045 -146.365 -44.715 -146.035 ;
        RECT -45.045 -147.725 -44.715 -147.395 ;
        RECT -45.045 -149.085 -44.715 -148.755 ;
        RECT -45.045 -150.445 -44.715 -150.115 ;
        RECT -45.045 -151.805 -44.715 -151.475 ;
        RECT -45.045 -153.165 -44.715 -152.835 ;
        RECT -45.045 -154.525 -44.715 -154.195 ;
        RECT -45.045 -155.885 -44.715 -155.555 ;
        RECT -45.045 -157.245 -44.715 -156.915 ;
        RECT -45.045 -158.605 -44.715 -158.275 ;
        RECT -45.045 -159.965 -44.715 -159.635 ;
        RECT -45.045 -161.325 -44.715 -160.995 ;
        RECT -45.045 -162.685 -44.715 -162.355 ;
        RECT -45.045 -164.045 -44.715 -163.715 ;
        RECT -45.045 -165.405 -44.715 -165.075 ;
        RECT -45.045 -166.765 -44.715 -166.435 ;
        RECT -45.045 -168.125 -44.715 -167.795 ;
        RECT -45.045 -169.485 -44.715 -169.155 ;
        RECT -45.045 -170.845 -44.715 -170.515 ;
        RECT -45.045 -172.205 -44.715 -171.875 ;
        RECT -45.045 -173.565 -44.715 -173.235 ;
        RECT -45.045 -174.925 -44.715 -174.595 ;
        RECT -45.045 -176.285 -44.715 -175.955 ;
        RECT -45.045 -177.645 -44.715 -177.315 ;
        RECT -45.045 -179.005 -44.715 -178.675 ;
        RECT -45.045 -180.365 -44.715 -180.035 ;
        RECT -45.045 -181.725 -44.715 -181.395 ;
        RECT -45.045 -183.085 -44.715 -182.755 ;
        RECT -45.045 -184.445 -44.715 -184.115 ;
        RECT -45.045 -185.805 -44.715 -185.475 ;
        RECT -45.045 -187.165 -44.715 -186.835 ;
        RECT -45.045 -188.525 -44.715 -188.195 ;
        RECT -45.045 -189.885 -44.715 -189.555 ;
        RECT -45.045 -191.245 -44.715 -190.915 ;
        RECT -45.045 -192.605 -44.715 -192.275 ;
        RECT -45.045 -193.965 -44.715 -193.635 ;
        RECT -45.045 -195.325 -44.715 -194.995 ;
        RECT -45.045 -196.685 -44.715 -196.355 ;
        RECT -45.045 -198.045 -44.715 -197.715 ;
        RECT -45.045 -199.405 -44.715 -199.075 ;
        RECT -45.045 -200.765 -44.715 -200.435 ;
        RECT -45.045 -202.125 -44.715 -201.795 ;
        RECT -45.045 -203.485 -44.715 -203.155 ;
        RECT -45.045 -204.845 -44.715 -204.515 ;
        RECT -45.045 -206.555 -44.715 -206.225 ;
        RECT -45.045 -207.565 -44.715 -207.235 ;
        RECT -45.045 -208.925 -44.715 -208.595 ;
        RECT -45.045 -211.645 -44.715 -211.315 ;
        RECT -45.045 -214.365 -44.715 -214.035 ;
        RECT -45.045 -215.725 -44.715 -215.395 ;
        RECT -45.045 -217.085 -44.715 -216.755 ;
        RECT -45.045 -218.445 -44.715 -218.115 ;
        RECT -45.045 -224.09 -44.715 -222.96 ;
        RECT -45.04 -224.205 -44.72 -139.235 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.685 132.52 -43.355 133.65 ;
        RECT -43.685 128.355 -43.355 128.685 ;
        RECT -43.685 126.995 -43.355 127.325 ;
        RECT -43.685 125.635 -43.355 125.965 ;
        RECT -43.685 124.275 -43.355 124.605 ;
        RECT -43.685 122.915 -43.355 123.245 ;
        RECT -43.685 121.555 -43.355 121.885 ;
        RECT -43.685 120.195 -43.355 120.525 ;
        RECT -43.685 118.835 -43.355 119.165 ;
        RECT -43.685 117.475 -43.355 117.805 ;
        RECT -43.685 116.115 -43.355 116.445 ;
        RECT -43.685 114.755 -43.355 115.085 ;
        RECT -43.685 113.395 -43.355 113.725 ;
        RECT -43.685 112.035 -43.355 112.365 ;
        RECT -43.685 110.675 -43.355 111.005 ;
        RECT -43.685 109.315 -43.355 109.645 ;
        RECT -43.685 107.955 -43.355 108.285 ;
        RECT -43.685 106.595 -43.355 106.925 ;
        RECT -43.685 105.235 -43.355 105.565 ;
        RECT -43.685 103.875 -43.355 104.205 ;
        RECT -43.685 102.515 -43.355 102.845 ;
        RECT -43.685 101.155 -43.355 101.485 ;
        RECT -43.685 99.795 -43.355 100.125 ;
        RECT -43.685 98.435 -43.355 98.765 ;
        RECT -43.685 97.075 -43.355 97.405 ;
        RECT -43.685 95.715 -43.355 96.045 ;
        RECT -43.685 94.355 -43.355 94.685 ;
        RECT -43.685 92.995 -43.355 93.325 ;
        RECT -43.685 91.635 -43.355 91.965 ;
        RECT -43.685 90.275 -43.355 90.605 ;
        RECT -43.685 88.915 -43.355 89.245 ;
        RECT -43.685 87.555 -43.355 87.885 ;
        RECT -43.685 86.195 -43.355 86.525 ;
        RECT -43.685 84.835 -43.355 85.165 ;
        RECT -43.685 83.475 -43.355 83.805 ;
        RECT -43.685 82.115 -43.355 82.445 ;
        RECT -43.685 80.755 -43.355 81.085 ;
        RECT -43.685 79.395 -43.355 79.725 ;
        RECT -43.685 78.035 -43.355 78.365 ;
        RECT -43.685 76.675 -43.355 77.005 ;
        RECT -43.685 75.315 -43.355 75.645 ;
        RECT -43.685 73.955 -43.355 74.285 ;
        RECT -43.685 71.64 -43.355 71.97 ;
        RECT -43.685 69.465 -43.355 69.795 ;
        RECT -43.685 68.615 -43.355 68.945 ;
        RECT -43.685 66.305 -43.355 66.635 ;
        RECT -43.685 65.455 -43.355 65.785 ;
        RECT -43.685 63.145 -43.355 63.475 ;
        RECT -43.685 62.295 -43.355 62.625 ;
        RECT -43.685 59.985 -43.355 60.315 ;
        RECT -43.685 59.135 -43.355 59.465 ;
        RECT -43.685 56.825 -43.355 57.155 ;
        RECT -43.685 55.975 -43.355 56.305 ;
        RECT -43.685 53.665 -43.355 53.995 ;
        RECT -43.685 52.815 -43.355 53.145 ;
        RECT -43.685 50.64 -43.355 50.97 ;
        RECT -43.685 48.115 -43.355 48.445 ;
        RECT -43.685 46.755 -43.355 47.085 ;
        RECT -43.685 45.395 -43.355 45.725 ;
        RECT -43.685 44.035 -43.355 44.365 ;
        RECT -43.685 42.675 -43.355 43.005 ;
        RECT -43.685 41.315 -43.355 41.645 ;
        RECT -43.685 39.955 -43.355 40.285 ;
        RECT -43.685 38.595 -43.355 38.925 ;
        RECT -43.685 37.235 -43.355 37.565 ;
        RECT -43.685 35.875 -43.355 36.205 ;
        RECT -43.685 34.515 -43.355 34.845 ;
        RECT -43.685 33.155 -43.355 33.485 ;
        RECT -43.685 31.795 -43.355 32.125 ;
        RECT -43.685 30.435 -43.355 30.765 ;
        RECT -43.685 29.075 -43.355 29.405 ;
        RECT -43.685 27.715 -43.355 28.045 ;
        RECT -43.685 26.355 -43.355 26.685 ;
        RECT -43.685 24.995 -43.355 25.325 ;
        RECT -43.685 23.635 -43.355 23.965 ;
        RECT -43.685 22.275 -43.355 22.605 ;
        RECT -43.685 20.915 -43.355 21.245 ;
        RECT -43.685 19.555 -43.355 19.885 ;
        RECT -43.685 18.195 -43.355 18.525 ;
        RECT -43.685 16.835 -43.355 17.165 ;
        RECT -43.685 15.475 -43.355 15.805 ;
        RECT -43.685 14.115 -43.355 14.445 ;
        RECT -43.685 12.755 -43.355 13.085 ;
        RECT -43.685 11.395 -43.355 11.725 ;
        RECT -43.685 10.035 -43.355 10.365 ;
        RECT -43.685 8.675 -43.355 9.005 ;
        RECT -43.685 7.315 -43.355 7.645 ;
        RECT -43.685 5.955 -43.355 6.285 ;
        RECT -43.685 4.595 -43.355 4.925 ;
        RECT -43.685 3.235 -43.355 3.565 ;
        RECT -43.685 1.875 -43.355 2.205 ;
        RECT -43.685 0.515 -43.355 0.845 ;
        RECT -43.685 -0.845 -43.355 -0.515 ;
        RECT -43.685 -2.205 -43.355 -1.875 ;
        RECT -43.685 -3.565 -43.355 -3.235 ;
        RECT -43.685 -4.925 -43.355 -4.595 ;
        RECT -43.685 -6.285 -43.355 -5.955 ;
        RECT -43.685 -7.645 -43.355 -7.315 ;
        RECT -43.685 -9.005 -43.355 -8.675 ;
        RECT -43.685 -11.725 -43.355 -11.395 ;
        RECT -43.685 -13.085 -43.355 -12.755 ;
        RECT -43.685 -14.445 -43.355 -14.115 ;
        RECT -43.685 -15.805 -43.355 -15.475 ;
        RECT -43.685 -17.165 -43.355 -16.835 ;
        RECT -43.685 -18.525 -43.355 -18.195 ;
        RECT -43.685 -19.885 -43.355 -19.555 ;
        RECT -43.685 -21.245 -43.355 -20.915 ;
        RECT -43.685 -22.605 -43.355 -22.275 ;
        RECT -43.685 -23.965 -43.355 -23.635 ;
        RECT -43.685 -25.325 -43.355 -24.995 ;
        RECT -43.685 -26.685 -43.355 -26.355 ;
        RECT -43.685 -28.045 -43.355 -27.715 ;
        RECT -43.685 -29.405 -43.355 -29.075 ;
        RECT -43.685 -32.125 -43.355 -31.795 ;
        RECT -43.685 -34.845 -43.355 -34.515 ;
        RECT -43.685 -37.565 -43.355 -37.235 ;
        RECT -43.685 -38.925 -43.355 -38.595 ;
        RECT -43.685 -40.285 -43.355 -39.955 ;
        RECT -43.685 -41.645 -43.355 -41.315 ;
        RECT -43.685 -43.005 -43.355 -42.675 ;
        RECT -43.685 -44.365 -43.355 -44.035 ;
        RECT -43.685 -45.725 -43.355 -45.395 ;
        RECT -43.685 -47.085 -43.355 -46.755 ;
        RECT -43.685 -48.445 -43.355 -48.115 ;
        RECT -43.685 -49.805 -43.355 -49.475 ;
        RECT -43.685 -51.165 -43.355 -50.835 ;
        RECT -43.685 -52.525 -43.355 -52.195 ;
        RECT -43.685 -53.885 -43.355 -53.555 ;
        RECT -43.685 -55.245 -43.355 -54.915 ;
        RECT -43.685 -56.605 -43.355 -56.275 ;
        RECT -43.685 -57.965 -43.355 -57.635 ;
        RECT -43.685 -59.325 -43.355 -58.995 ;
        RECT -43.685 -60.685 -43.355 -60.355 ;
        RECT -43.685 -62.045 -43.355 -61.715 ;
        RECT -43.685 -63.405 -43.355 -63.075 ;
        RECT -43.685 -64.765 -43.355 -64.435 ;
        RECT -43.685 -66.125 -43.355 -65.795 ;
        RECT -43.685 -67.485 -43.355 -67.155 ;
        RECT -43.685 -68.845 -43.355 -68.515 ;
        RECT -43.685 -70.205 -43.355 -69.875 ;
        RECT -43.685 -71.565 -43.355 -71.235 ;
        RECT -43.685 -72.925 -43.355 -72.595 ;
        RECT -43.685 -74.285 -43.355 -73.955 ;
        RECT -43.685 -75.645 -43.355 -75.315 ;
        RECT -43.685 -77.005 -43.355 -76.675 ;
        RECT -43.685 -78.365 -43.355 -78.035 ;
        RECT -43.685 -79.725 -43.355 -79.395 ;
        RECT -43.685 -81.085 -43.355 -80.755 ;
        RECT -43.685 -82.445 -43.355 -82.115 ;
        RECT -43.685 -83.805 -43.355 -83.475 ;
        RECT -43.685 -85.165 -43.355 -84.835 ;
        RECT -43.685 -86.525 -43.355 -86.195 ;
        RECT -43.685 -87.885 -43.355 -87.555 ;
        RECT -43.685 -89.245 -43.355 -88.915 ;
        RECT -43.685 -90.605 -43.355 -90.275 ;
        RECT -43.685 -91.965 -43.355 -91.635 ;
        RECT -43.685 -93.325 -43.355 -92.995 ;
        RECT -43.685 -94.685 -43.355 -94.355 ;
        RECT -43.685 -96.045 -43.355 -95.715 ;
        RECT -43.685 -97.405 -43.355 -97.075 ;
        RECT -43.685 -98.765 -43.355 -98.435 ;
        RECT -43.685 -100.125 -43.355 -99.795 ;
        RECT -43.685 -101.485 -43.355 -101.155 ;
        RECT -43.685 -102.845 -43.355 -102.515 ;
        RECT -43.685 -104.205 -43.355 -103.875 ;
        RECT -43.685 -105.565 -43.355 -105.235 ;
        RECT -43.685 -106.925 -43.355 -106.595 ;
        RECT -43.685 -108.285 -43.355 -107.955 ;
        RECT -43.685 -109.645 -43.355 -109.315 ;
        RECT -43.685 -111.005 -43.355 -110.675 ;
        RECT -43.685 -111.87 -43.355 -111.54 ;
        RECT -43.685 -113.725 -43.355 -113.395 ;
        RECT -43.685 -115.085 -43.355 -114.755 ;
        RECT -43.685 -116.445 -43.355 -116.115 ;
        RECT -43.685 -117.805 -43.355 -117.475 ;
        RECT -43.685 -120.525 -43.355 -120.195 ;
        RECT -43.685 -121.885 -43.355 -121.555 ;
        RECT -43.685 -123.245 -43.355 -122.915 ;
        RECT -43.685 -124.71 -43.355 -124.38 ;
        RECT -43.685 -125.965 -43.355 -125.635 ;
        RECT -43.685 -127.325 -43.355 -126.995 ;
        RECT -43.685 -130.045 -43.355 -129.715 ;
        RECT -43.685 -132.765 -43.355 -132.435 ;
        RECT -43.685 -134.125 -43.355 -133.795 ;
        RECT -43.685 -135.485 -43.355 -135.155 ;
        RECT -43.685 -136.845 -43.355 -136.515 ;
        RECT -43.685 -138.205 -43.355 -137.875 ;
        RECT -43.685 -139.565 -43.355 -139.235 ;
        RECT -43.685 -142.285 -43.355 -141.955 ;
        RECT -43.685 -143.645 -43.355 -143.315 ;
        RECT -43.685 -145.005 -43.355 -144.675 ;
        RECT -43.685 -146.365 -43.355 -146.035 ;
        RECT -43.685 -147.725 -43.355 -147.395 ;
        RECT -43.685 -149.085 -43.355 -148.755 ;
        RECT -43.685 -150.445 -43.355 -150.115 ;
        RECT -43.685 -151.805 -43.355 -151.475 ;
        RECT -43.685 -153.165 -43.355 -152.835 ;
        RECT -43.685 -154.525 -43.355 -154.195 ;
        RECT -43.685 -155.885 -43.355 -155.555 ;
        RECT -43.685 -157.245 -43.355 -156.915 ;
        RECT -43.685 -158.605 -43.355 -158.275 ;
        RECT -43.685 -159.965 -43.355 -159.635 ;
        RECT -43.685 -161.325 -43.355 -160.995 ;
        RECT -43.685 -162.685 -43.355 -162.355 ;
        RECT -43.685 -164.045 -43.355 -163.715 ;
        RECT -43.685 -165.405 -43.355 -165.075 ;
        RECT -43.685 -166.765 -43.355 -166.435 ;
        RECT -43.685 -168.125 -43.355 -167.795 ;
        RECT -43.685 -169.485 -43.355 -169.155 ;
        RECT -43.685 -170.845 -43.355 -170.515 ;
        RECT -43.685 -172.205 -43.355 -171.875 ;
        RECT -43.685 -173.565 -43.355 -173.235 ;
        RECT -43.685 -174.925 -43.355 -174.595 ;
        RECT -43.685 -176.285 -43.355 -175.955 ;
        RECT -43.685 -177.645 -43.355 -177.315 ;
        RECT -43.685 -179.005 -43.355 -178.675 ;
        RECT -43.685 -180.365 -43.355 -180.035 ;
        RECT -43.685 -181.725 -43.355 -181.395 ;
        RECT -43.685 -183.085 -43.355 -182.755 ;
        RECT -43.685 -184.445 -43.355 -184.115 ;
        RECT -43.685 -185.805 -43.355 -185.475 ;
        RECT -43.685 -187.165 -43.355 -186.835 ;
        RECT -43.685 -188.525 -43.355 -188.195 ;
        RECT -43.685 -189.885 -43.355 -189.555 ;
        RECT -43.685 -191.245 -43.355 -190.915 ;
        RECT -43.685 -192.605 -43.355 -192.275 ;
        RECT -43.685 -193.965 -43.355 -193.635 ;
        RECT -43.685 -195.325 -43.355 -194.995 ;
        RECT -43.685 -196.685 -43.355 -196.355 ;
        RECT -43.685 -198.045 -43.355 -197.715 ;
        RECT -43.685 -199.405 -43.355 -199.075 ;
        RECT -43.685 -200.765 -43.355 -200.435 ;
        RECT -43.685 -202.125 -43.355 -201.795 ;
        RECT -43.685 -203.485 -43.355 -203.155 ;
        RECT -43.685 -204.845 -43.355 -204.515 ;
        RECT -43.685 -206.555 -43.355 -206.225 ;
        RECT -43.685 -207.565 -43.355 -207.235 ;
        RECT -43.685 -208.925 -43.355 -208.595 ;
        RECT -43.685 -210.285 -43.355 -209.955 ;
        RECT -43.685 -211.645 -43.355 -211.315 ;
        RECT -43.685 -214.365 -43.355 -214.035 ;
        RECT -43.685 -215.725 -43.355 -215.395 ;
        RECT -43.685 -217.085 -43.355 -216.755 ;
        RECT -43.685 -218.445 -43.355 -218.115 ;
        RECT -43.685 -224.09 -43.355 -222.96 ;
        RECT -43.68 -224.205 -43.36 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -42.325 -172.205 -41.995 -171.875 ;
        RECT -42.325 -173.565 -41.995 -173.235 ;
        RECT -42.325 -174.925 -41.995 -174.595 ;
        RECT -42.325 -176.285 -41.995 -175.955 ;
        RECT -42.325 -177.645 -41.995 -177.315 ;
        RECT -42.325 -179.005 -41.995 -178.675 ;
        RECT -42.325 -180.365 -41.995 -180.035 ;
        RECT -42.325 -181.725 -41.995 -181.395 ;
        RECT -42.325 -183.085 -41.995 -182.755 ;
        RECT -42.325 -184.445 -41.995 -184.115 ;
        RECT -42.325 -185.805 -41.995 -185.475 ;
        RECT -42.325 -187.165 -41.995 -186.835 ;
        RECT -42.325 -188.525 -41.995 -188.195 ;
        RECT -42.325 -189.885 -41.995 -189.555 ;
        RECT -42.325 -191.245 -41.995 -190.915 ;
        RECT -42.325 -192.605 -41.995 -192.275 ;
        RECT -42.325 -193.965 -41.995 -193.635 ;
        RECT -42.325 -195.325 -41.995 -194.995 ;
        RECT -42.325 -196.685 -41.995 -196.355 ;
        RECT -42.325 -198.045 -41.995 -197.715 ;
        RECT -42.325 -199.405 -41.995 -199.075 ;
        RECT -42.325 -200.765 -41.995 -200.435 ;
        RECT -42.325 -202.125 -41.995 -201.795 ;
        RECT -42.325 -203.485 -41.995 -203.155 ;
        RECT -42.325 -204.845 -41.995 -204.515 ;
        RECT -42.325 -206.555 -41.995 -206.225 ;
        RECT -42.325 -207.565 -41.995 -207.235 ;
        RECT -42.325 -208.925 -41.995 -208.595 ;
        RECT -42.325 -210.285 -41.995 -209.955 ;
        RECT -42.325 -214.365 -41.995 -214.035 ;
        RECT -42.325 -215.725 -41.995 -215.395 ;
        RECT -42.325 -217.085 -41.995 -216.755 ;
        RECT -42.325 -218.445 -41.995 -218.115 ;
        RECT -42.325 -224.09 -41.995 -222.96 ;
        RECT -42.32 -224.205 -42 133.765 ;
        RECT -42.325 132.52 -41.995 133.65 ;
        RECT -42.325 128.355 -41.995 128.685 ;
        RECT -42.325 126.995 -41.995 127.325 ;
        RECT -42.325 125.635 -41.995 125.965 ;
        RECT -42.325 124.275 -41.995 124.605 ;
        RECT -42.325 122.915 -41.995 123.245 ;
        RECT -42.325 121.555 -41.995 121.885 ;
        RECT -42.325 120.195 -41.995 120.525 ;
        RECT -42.325 118.835 -41.995 119.165 ;
        RECT -42.325 117.475 -41.995 117.805 ;
        RECT -42.325 116.115 -41.995 116.445 ;
        RECT -42.325 114.755 -41.995 115.085 ;
        RECT -42.325 113.395 -41.995 113.725 ;
        RECT -42.325 112.035 -41.995 112.365 ;
        RECT -42.325 110.675 -41.995 111.005 ;
        RECT -42.325 109.315 -41.995 109.645 ;
        RECT -42.325 107.955 -41.995 108.285 ;
        RECT -42.325 106.595 -41.995 106.925 ;
        RECT -42.325 105.235 -41.995 105.565 ;
        RECT -42.325 103.875 -41.995 104.205 ;
        RECT -42.325 102.515 -41.995 102.845 ;
        RECT -42.325 101.155 -41.995 101.485 ;
        RECT -42.325 99.795 -41.995 100.125 ;
        RECT -42.325 98.435 -41.995 98.765 ;
        RECT -42.325 97.075 -41.995 97.405 ;
        RECT -42.325 95.715 -41.995 96.045 ;
        RECT -42.325 94.355 -41.995 94.685 ;
        RECT -42.325 92.995 -41.995 93.325 ;
        RECT -42.325 91.635 -41.995 91.965 ;
        RECT -42.325 90.275 -41.995 90.605 ;
        RECT -42.325 88.915 -41.995 89.245 ;
        RECT -42.325 87.555 -41.995 87.885 ;
        RECT -42.325 86.195 -41.995 86.525 ;
        RECT -42.325 84.835 -41.995 85.165 ;
        RECT -42.325 83.475 -41.995 83.805 ;
        RECT -42.325 82.115 -41.995 82.445 ;
        RECT -42.325 80.755 -41.995 81.085 ;
        RECT -42.325 79.395 -41.995 79.725 ;
        RECT -42.325 78.035 -41.995 78.365 ;
        RECT -42.325 76.675 -41.995 77.005 ;
        RECT -42.325 75.315 -41.995 75.645 ;
        RECT -42.325 73.955 -41.995 74.285 ;
        RECT -42.325 71.64 -41.995 71.97 ;
        RECT -42.325 69.465 -41.995 69.795 ;
        RECT -42.325 68.615 -41.995 68.945 ;
        RECT -42.325 66.305 -41.995 66.635 ;
        RECT -42.325 65.455 -41.995 65.785 ;
        RECT -42.325 63.145 -41.995 63.475 ;
        RECT -42.325 62.295 -41.995 62.625 ;
        RECT -42.325 59.985 -41.995 60.315 ;
        RECT -42.325 59.135 -41.995 59.465 ;
        RECT -42.325 56.825 -41.995 57.155 ;
        RECT -42.325 55.975 -41.995 56.305 ;
        RECT -42.325 53.665 -41.995 53.995 ;
        RECT -42.325 52.815 -41.995 53.145 ;
        RECT -42.325 50.64 -41.995 50.97 ;
        RECT -42.325 48.115 -41.995 48.445 ;
        RECT -42.325 46.755 -41.995 47.085 ;
        RECT -42.325 45.395 -41.995 45.725 ;
        RECT -42.325 44.035 -41.995 44.365 ;
        RECT -42.325 42.675 -41.995 43.005 ;
        RECT -42.325 41.315 -41.995 41.645 ;
        RECT -42.325 39.955 -41.995 40.285 ;
        RECT -42.325 38.595 -41.995 38.925 ;
        RECT -42.325 37.235 -41.995 37.565 ;
        RECT -42.325 35.875 -41.995 36.205 ;
        RECT -42.325 34.515 -41.995 34.845 ;
        RECT -42.325 33.155 -41.995 33.485 ;
        RECT -42.325 31.795 -41.995 32.125 ;
        RECT -42.325 30.435 -41.995 30.765 ;
        RECT -42.325 29.075 -41.995 29.405 ;
        RECT -42.325 27.715 -41.995 28.045 ;
        RECT -42.325 26.355 -41.995 26.685 ;
        RECT -42.325 24.995 -41.995 25.325 ;
        RECT -42.325 23.635 -41.995 23.965 ;
        RECT -42.325 22.275 -41.995 22.605 ;
        RECT -42.325 20.915 -41.995 21.245 ;
        RECT -42.325 19.555 -41.995 19.885 ;
        RECT -42.325 18.195 -41.995 18.525 ;
        RECT -42.325 16.835 -41.995 17.165 ;
        RECT -42.325 15.475 -41.995 15.805 ;
        RECT -42.325 14.115 -41.995 14.445 ;
        RECT -42.325 12.755 -41.995 13.085 ;
        RECT -42.325 11.395 -41.995 11.725 ;
        RECT -42.325 10.035 -41.995 10.365 ;
        RECT -42.325 8.675 -41.995 9.005 ;
        RECT -42.325 7.315 -41.995 7.645 ;
        RECT -42.325 5.955 -41.995 6.285 ;
        RECT -42.325 4.595 -41.995 4.925 ;
        RECT -42.325 3.235 -41.995 3.565 ;
        RECT -42.325 1.875 -41.995 2.205 ;
        RECT -42.325 0.515 -41.995 0.845 ;
        RECT -42.325 -0.845 -41.995 -0.515 ;
        RECT -42.325 -2.205 -41.995 -1.875 ;
        RECT -42.325 -3.565 -41.995 -3.235 ;
        RECT -42.325 -4.925 -41.995 -4.595 ;
        RECT -42.325 -6.285 -41.995 -5.955 ;
        RECT -42.325 -7.645 -41.995 -7.315 ;
        RECT -42.325 -9.005 -41.995 -8.675 ;
        RECT -42.325 -11.725 -41.995 -11.395 ;
        RECT -42.325 -13.085 -41.995 -12.755 ;
        RECT -42.325 -14.445 -41.995 -14.115 ;
        RECT -42.325 -15.805 -41.995 -15.475 ;
        RECT -42.325 -17.165 -41.995 -16.835 ;
        RECT -42.325 -18.525 -41.995 -18.195 ;
        RECT -42.325 -19.885 -41.995 -19.555 ;
        RECT -42.325 -21.245 -41.995 -20.915 ;
        RECT -42.325 -22.605 -41.995 -22.275 ;
        RECT -42.325 -23.965 -41.995 -23.635 ;
        RECT -42.325 -26.685 -41.995 -26.355 ;
        RECT -42.325 -28.045 -41.995 -27.715 ;
        RECT -42.325 -29.405 -41.995 -29.075 ;
        RECT -42.325 -32.125 -41.995 -31.795 ;
        RECT -42.325 -34.845 -41.995 -34.515 ;
        RECT -42.325 -37.565 -41.995 -37.235 ;
        RECT -42.325 -38.925 -41.995 -38.595 ;
        RECT -42.325 -40.285 -41.995 -39.955 ;
        RECT -42.325 -41.645 -41.995 -41.315 ;
        RECT -42.325 -43.005 -41.995 -42.675 ;
        RECT -42.325 -44.365 -41.995 -44.035 ;
        RECT -42.325 -45.725 -41.995 -45.395 ;
        RECT -42.325 -47.085 -41.995 -46.755 ;
        RECT -42.325 -48.445 -41.995 -48.115 ;
        RECT -42.325 -49.805 -41.995 -49.475 ;
        RECT -42.325 -51.165 -41.995 -50.835 ;
        RECT -42.325 -52.525 -41.995 -52.195 ;
        RECT -42.325 -53.885 -41.995 -53.555 ;
        RECT -42.325 -55.245 -41.995 -54.915 ;
        RECT -42.325 -56.605 -41.995 -56.275 ;
        RECT -42.325 -57.965 -41.995 -57.635 ;
        RECT -42.325 -59.325 -41.995 -58.995 ;
        RECT -42.325 -60.685 -41.995 -60.355 ;
        RECT -42.325 -62.045 -41.995 -61.715 ;
        RECT -42.325 -63.405 -41.995 -63.075 ;
        RECT -42.325 -64.765 -41.995 -64.435 ;
        RECT -42.325 -66.125 -41.995 -65.795 ;
        RECT -42.325 -67.485 -41.995 -67.155 ;
        RECT -42.325 -68.845 -41.995 -68.515 ;
        RECT -42.325 -70.205 -41.995 -69.875 ;
        RECT -42.325 -71.565 -41.995 -71.235 ;
        RECT -42.325 -72.925 -41.995 -72.595 ;
        RECT -42.325 -74.285 -41.995 -73.955 ;
        RECT -42.325 -75.645 -41.995 -75.315 ;
        RECT -42.325 -77.005 -41.995 -76.675 ;
        RECT -42.325 -78.365 -41.995 -78.035 ;
        RECT -42.325 -79.725 -41.995 -79.395 ;
        RECT -42.325 -81.085 -41.995 -80.755 ;
        RECT -42.325 -82.445 -41.995 -82.115 ;
        RECT -42.325 -83.805 -41.995 -83.475 ;
        RECT -42.325 -85.165 -41.995 -84.835 ;
        RECT -42.325 -86.525 -41.995 -86.195 ;
        RECT -42.325 -87.885 -41.995 -87.555 ;
        RECT -42.325 -89.245 -41.995 -88.915 ;
        RECT -42.325 -90.605 -41.995 -90.275 ;
        RECT -42.325 -91.965 -41.995 -91.635 ;
        RECT -42.325 -93.325 -41.995 -92.995 ;
        RECT -42.325 -94.685 -41.995 -94.355 ;
        RECT -42.325 -96.045 -41.995 -95.715 ;
        RECT -42.325 -97.405 -41.995 -97.075 ;
        RECT -42.325 -98.765 -41.995 -98.435 ;
        RECT -42.325 -100.125 -41.995 -99.795 ;
        RECT -42.325 -101.485 -41.995 -101.155 ;
        RECT -42.325 -102.845 -41.995 -102.515 ;
        RECT -42.325 -104.205 -41.995 -103.875 ;
        RECT -42.325 -105.565 -41.995 -105.235 ;
        RECT -42.325 -106.925 -41.995 -106.595 ;
        RECT -42.325 -108.285 -41.995 -107.955 ;
        RECT -42.325 -109.645 -41.995 -109.315 ;
        RECT -42.325 -111.005 -41.995 -110.675 ;
        RECT -42.325 -111.87 -41.995 -111.54 ;
        RECT -42.325 -113.725 -41.995 -113.395 ;
        RECT -42.325 -115.085 -41.995 -114.755 ;
        RECT -42.325 -116.445 -41.995 -116.115 ;
        RECT -42.325 -117.805 -41.995 -117.475 ;
        RECT -42.325 -120.525 -41.995 -120.195 ;
        RECT -42.325 -121.885 -41.995 -121.555 ;
        RECT -42.325 -123.245 -41.995 -122.915 ;
        RECT -42.325 -124.71 -41.995 -124.38 ;
        RECT -42.325 -125.965 -41.995 -125.635 ;
        RECT -42.325 -127.325 -41.995 -126.995 ;
        RECT -42.325 -130.045 -41.995 -129.715 ;
        RECT -42.325 -132.765 -41.995 -132.435 ;
        RECT -42.325 -134.125 -41.995 -133.795 ;
        RECT -42.325 -135.485 -41.995 -135.155 ;
        RECT -42.325 -136.845 -41.995 -136.515 ;
        RECT -42.325 -138.205 -41.995 -137.875 ;
        RECT -42.325 -139.565 -41.995 -139.235 ;
        RECT -42.325 -142.285 -41.995 -141.955 ;
        RECT -42.325 -143.645 -41.995 -143.315 ;
        RECT -42.325 -145.005 -41.995 -144.675 ;
        RECT -42.325 -146.365 -41.995 -146.035 ;
        RECT -42.325 -147.725 -41.995 -147.395 ;
        RECT -42.325 -149.085 -41.995 -148.755 ;
        RECT -42.325 -150.445 -41.995 -150.115 ;
        RECT -42.325 -151.805 -41.995 -151.475 ;
        RECT -42.325 -153.165 -41.995 -152.835 ;
        RECT -42.325 -154.525 -41.995 -154.195 ;
        RECT -42.325 -155.885 -41.995 -155.555 ;
        RECT -42.325 -157.245 -41.995 -156.915 ;
        RECT -42.325 -158.605 -41.995 -158.275 ;
        RECT -42.325 -159.965 -41.995 -159.635 ;
        RECT -42.325 -161.325 -41.995 -160.995 ;
        RECT -42.325 -162.685 -41.995 -162.355 ;
        RECT -42.325 -164.045 -41.995 -163.715 ;
        RECT -42.325 -165.405 -41.995 -165.075 ;
        RECT -42.325 -166.765 -41.995 -166.435 ;
        RECT -42.325 -168.125 -41.995 -167.795 ;
        RECT -42.325 -169.485 -41.995 -169.155 ;
        RECT -42.325 -170.845 -41.995 -170.515 ;
    END
    PORT
      LAYER met3 ;
        RECT -54.565 132.52 -54.235 133.65 ;
        RECT -54.565 128.355 -54.235 128.685 ;
        RECT -54.565 126.995 -54.235 127.325 ;
        RECT -54.565 125.635 -54.235 125.965 ;
        RECT -54.565 124.275 -54.235 124.605 ;
        RECT -54.565 122.915 -54.235 123.245 ;
        RECT -54.565 121.555 -54.235 121.885 ;
        RECT -54.565 120.195 -54.235 120.525 ;
        RECT -54.565 118.835 -54.235 119.165 ;
        RECT -54.565 117.475 -54.235 117.805 ;
        RECT -54.565 116.115 -54.235 116.445 ;
        RECT -54.565 114.755 -54.235 115.085 ;
        RECT -54.565 113.395 -54.235 113.725 ;
        RECT -54.565 112.035 -54.235 112.365 ;
        RECT -54.565 110.675 -54.235 111.005 ;
        RECT -54.565 109.315 -54.235 109.645 ;
        RECT -54.565 107.955 -54.235 108.285 ;
        RECT -54.565 106.595 -54.235 106.925 ;
        RECT -54.565 105.235 -54.235 105.565 ;
        RECT -54.565 103.875 -54.235 104.205 ;
        RECT -54.565 102.515 -54.235 102.845 ;
        RECT -54.565 101.155 -54.235 101.485 ;
        RECT -54.565 99.795 -54.235 100.125 ;
        RECT -54.565 98.435 -54.235 98.765 ;
        RECT -54.565 97.075 -54.235 97.405 ;
        RECT -54.565 95.715 -54.235 96.045 ;
        RECT -54.565 94.355 -54.235 94.685 ;
        RECT -54.565 92.995 -54.235 93.325 ;
        RECT -54.565 91.635 -54.235 91.965 ;
        RECT -54.565 90.275 -54.235 90.605 ;
        RECT -54.565 88.915 -54.235 89.245 ;
        RECT -54.565 87.555 -54.235 87.885 ;
        RECT -54.565 86.195 -54.235 86.525 ;
        RECT -54.565 84.835 -54.235 85.165 ;
        RECT -54.565 83.475 -54.235 83.805 ;
        RECT -54.565 82.115 -54.235 82.445 ;
        RECT -54.565 80.755 -54.235 81.085 ;
        RECT -54.565 79.395 -54.235 79.725 ;
        RECT -54.565 78.035 -54.235 78.365 ;
        RECT -54.565 76.675 -54.235 77.005 ;
        RECT -54.565 75.315 -54.235 75.645 ;
        RECT -54.565 73.955 -54.235 74.285 ;
        RECT -54.565 71.64 -54.235 71.97 ;
        RECT -54.565 69.465 -54.235 69.795 ;
        RECT -54.565 68.615 -54.235 68.945 ;
        RECT -54.565 66.305 -54.235 66.635 ;
        RECT -54.565 65.455 -54.235 65.785 ;
        RECT -54.565 63.145 -54.235 63.475 ;
        RECT -54.565 62.295 -54.235 62.625 ;
        RECT -54.565 59.985 -54.235 60.315 ;
        RECT -54.565 59.135 -54.235 59.465 ;
        RECT -54.565 56.825 -54.235 57.155 ;
        RECT -54.565 55.975 -54.235 56.305 ;
        RECT -54.565 53.665 -54.235 53.995 ;
        RECT -54.565 52.815 -54.235 53.145 ;
        RECT -54.565 50.64 -54.235 50.97 ;
        RECT -54.565 48.115 -54.235 48.445 ;
        RECT -54.565 46.755 -54.235 47.085 ;
        RECT -54.565 45.395 -54.235 45.725 ;
        RECT -54.565 44.035 -54.235 44.365 ;
        RECT -54.565 42.675 -54.235 43.005 ;
        RECT -54.565 41.315 -54.235 41.645 ;
        RECT -54.565 39.955 -54.235 40.285 ;
        RECT -54.565 38.595 -54.235 38.925 ;
        RECT -54.565 37.235 -54.235 37.565 ;
        RECT -54.565 35.875 -54.235 36.205 ;
        RECT -54.565 34.515 -54.235 34.845 ;
        RECT -54.565 33.155 -54.235 33.485 ;
        RECT -54.565 31.795 -54.235 32.125 ;
        RECT -54.565 30.435 -54.235 30.765 ;
        RECT -54.565 29.075 -54.235 29.405 ;
        RECT -54.565 27.715 -54.235 28.045 ;
        RECT -54.565 26.355 -54.235 26.685 ;
        RECT -54.565 24.995 -54.235 25.325 ;
        RECT -54.565 23.635 -54.235 23.965 ;
        RECT -54.565 22.275 -54.235 22.605 ;
        RECT -54.565 20.915 -54.235 21.245 ;
        RECT -54.565 19.555 -54.235 19.885 ;
        RECT -54.565 18.195 -54.235 18.525 ;
        RECT -54.565 16.835 -54.235 17.165 ;
        RECT -54.565 15.475 -54.235 15.805 ;
        RECT -54.565 14.115 -54.235 14.445 ;
        RECT -54.565 12.755 -54.235 13.085 ;
        RECT -54.565 11.395 -54.235 11.725 ;
        RECT -54.565 10.035 -54.235 10.365 ;
        RECT -54.565 8.675 -54.235 9.005 ;
        RECT -54.565 7.315 -54.235 7.645 ;
        RECT -54.565 5.955 -54.235 6.285 ;
        RECT -54.565 4.595 -54.235 4.925 ;
        RECT -54.565 3.235 -54.235 3.565 ;
        RECT -54.565 1.875 -54.235 2.205 ;
        RECT -54.565 0.515 -54.235 0.845 ;
        RECT -54.565 -0.845 -54.235 -0.515 ;
        RECT -54.565 -2.205 -54.235 -1.875 ;
        RECT -54.565 -3.565 -54.235 -3.235 ;
        RECT -54.565 -4.925 -54.235 -4.595 ;
        RECT -54.565 -6.285 -54.235 -5.955 ;
        RECT -54.565 -7.645 -54.235 -7.315 ;
        RECT -54.565 -9.005 -54.235 -8.675 ;
        RECT -54.565 -10.365 -54.235 -10.035 ;
        RECT -54.565 -11.725 -54.235 -11.395 ;
        RECT -54.565 -13.085 -54.235 -12.755 ;
        RECT -54.565 -14.445 -54.235 -14.115 ;
        RECT -54.565 -15.805 -54.235 -15.475 ;
        RECT -54.565 -17.165 -54.235 -16.835 ;
        RECT -54.565 -18.525 -54.235 -18.195 ;
        RECT -54.565 -19.885 -54.235 -19.555 ;
        RECT -54.565 -21.245 -54.235 -20.915 ;
        RECT -54.565 -22.605 -54.235 -22.275 ;
        RECT -54.565 -23.965 -54.235 -23.635 ;
        RECT -54.565 -25.325 -54.235 -24.995 ;
        RECT -54.565 -26.685 -54.235 -26.355 ;
        RECT -54.565 -28.045 -54.235 -27.715 ;
        RECT -54.565 -29.405 -54.235 -29.075 ;
        RECT -54.565 -30.765 -54.235 -30.435 ;
        RECT -54.565 -32.125 -54.235 -31.795 ;
        RECT -54.565 -33.485 -54.235 -33.155 ;
        RECT -54.565 -34.845 -54.235 -34.515 ;
        RECT -54.565 -36.205 -54.235 -35.875 ;
        RECT -54.565 -37.565 -54.235 -37.235 ;
        RECT -54.565 -38.925 -54.235 -38.595 ;
        RECT -54.565 -40.285 -54.235 -39.955 ;
        RECT -54.565 -41.645 -54.235 -41.315 ;
        RECT -54.565 -43.005 -54.235 -42.675 ;
        RECT -54.565 -44.365 -54.235 -44.035 ;
        RECT -54.565 -45.725 -54.235 -45.395 ;
        RECT -54.565 -47.085 -54.235 -46.755 ;
        RECT -54.565 -48.445 -54.235 -48.115 ;
        RECT -54.565 -49.805 -54.235 -49.475 ;
        RECT -54.565 -51.165 -54.235 -50.835 ;
        RECT -54.565 -52.525 -54.235 -52.195 ;
        RECT -54.565 -53.885 -54.235 -53.555 ;
        RECT -54.565 -55.245 -54.235 -54.915 ;
        RECT -54.565 -56.605 -54.235 -56.275 ;
        RECT -54.565 -57.965 -54.235 -57.635 ;
        RECT -54.565 -59.325 -54.235 -58.995 ;
        RECT -54.565 -60.685 -54.235 -60.355 ;
        RECT -54.565 -62.045 -54.235 -61.715 ;
        RECT -54.565 -63.405 -54.235 -63.075 ;
        RECT -54.565 -64.765 -54.235 -64.435 ;
        RECT -54.565 -66.125 -54.235 -65.795 ;
        RECT -54.565 -67.485 -54.235 -67.155 ;
        RECT -54.565 -68.845 -54.235 -68.515 ;
        RECT -54.565 -70.205 -54.235 -69.875 ;
        RECT -54.565 -71.565 -54.235 -71.235 ;
        RECT -54.565 -72.925 -54.235 -72.595 ;
        RECT -54.565 -74.285 -54.235 -73.955 ;
        RECT -54.565 -75.645 -54.235 -75.315 ;
        RECT -54.565 -77.005 -54.235 -76.675 ;
        RECT -54.565 -78.365 -54.235 -78.035 ;
        RECT -54.565 -79.725 -54.235 -79.395 ;
        RECT -54.565 -81.085 -54.235 -80.755 ;
        RECT -54.565 -82.445 -54.235 -82.115 ;
        RECT -54.565 -83.805 -54.235 -83.475 ;
        RECT -54.565 -85.165 -54.235 -84.835 ;
        RECT -54.565 -86.525 -54.235 -86.195 ;
        RECT -54.565 -87.885 -54.235 -87.555 ;
        RECT -54.565 -89.245 -54.235 -88.915 ;
        RECT -54.565 -90.605 -54.235 -90.275 ;
        RECT -54.565 -91.965 -54.235 -91.635 ;
        RECT -54.565 -93.325 -54.235 -92.995 ;
        RECT -54.565 -94.685 -54.235 -94.355 ;
        RECT -54.565 -96.045 -54.235 -95.715 ;
        RECT -54.565 -97.405 -54.235 -97.075 ;
        RECT -54.565 -98.765 -54.235 -98.435 ;
        RECT -54.565 -100.125 -54.235 -99.795 ;
        RECT -54.565 -101.485 -54.235 -101.155 ;
        RECT -54.565 -102.845 -54.235 -102.515 ;
        RECT -54.565 -104.205 -54.235 -103.875 ;
        RECT -54.565 -105.565 -54.235 -105.235 ;
        RECT -54.565 -106.925 -54.235 -106.595 ;
        RECT -54.565 -108.285 -54.235 -107.955 ;
        RECT -54.565 -109.645 -54.235 -109.315 ;
        RECT -54.565 -111.005 -54.235 -110.675 ;
        RECT -54.565 -111.87 -54.235 -111.54 ;
        RECT -54.565 -113.725 -54.235 -113.395 ;
        RECT -54.565 -115.085 -54.235 -114.755 ;
        RECT -54.565 -116.445 -54.235 -116.115 ;
        RECT -54.565 -117.805 -54.235 -117.475 ;
        RECT -54.565 -120.525 -54.235 -120.195 ;
        RECT -54.565 -121.885 -54.235 -121.555 ;
        RECT -54.565 -123.245 -54.235 -122.915 ;
        RECT -54.565 -124.71 -54.235 -124.38 ;
        RECT -54.565 -125.965 -54.235 -125.635 ;
        RECT -54.565 -127.325 -54.235 -126.995 ;
        RECT -54.565 -130.045 -54.235 -129.715 ;
        RECT -54.56 -133.44 -54.24 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -54.565 -214.365 -54.235 -214.035 ;
        RECT -54.565 -215.725 -54.235 -215.395 ;
        RECT -54.565 -217.085 -54.235 -216.755 ;
        RECT -54.565 -218.445 -54.235 -218.115 ;
        RECT -54.565 -224.09 -54.235 -222.96 ;
        RECT -54.56 -224.205 -54.24 -212 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.205 132.52 -52.875 133.65 ;
        RECT -53.205 128.355 -52.875 128.685 ;
        RECT -53.205 126.995 -52.875 127.325 ;
        RECT -53.205 125.635 -52.875 125.965 ;
        RECT -53.205 124.275 -52.875 124.605 ;
        RECT -53.205 122.915 -52.875 123.245 ;
        RECT -53.205 121.555 -52.875 121.885 ;
        RECT -53.205 120.195 -52.875 120.525 ;
        RECT -53.205 118.835 -52.875 119.165 ;
        RECT -53.205 117.475 -52.875 117.805 ;
        RECT -53.205 116.115 -52.875 116.445 ;
        RECT -53.205 114.755 -52.875 115.085 ;
        RECT -53.205 113.395 -52.875 113.725 ;
        RECT -53.205 112.035 -52.875 112.365 ;
        RECT -53.205 110.675 -52.875 111.005 ;
        RECT -53.205 109.315 -52.875 109.645 ;
        RECT -53.205 107.955 -52.875 108.285 ;
        RECT -53.205 106.595 -52.875 106.925 ;
        RECT -53.205 105.235 -52.875 105.565 ;
        RECT -53.205 103.875 -52.875 104.205 ;
        RECT -53.205 102.515 -52.875 102.845 ;
        RECT -53.205 101.155 -52.875 101.485 ;
        RECT -53.205 99.795 -52.875 100.125 ;
        RECT -53.205 98.435 -52.875 98.765 ;
        RECT -53.205 97.075 -52.875 97.405 ;
        RECT -53.205 95.715 -52.875 96.045 ;
        RECT -53.205 94.355 -52.875 94.685 ;
        RECT -53.205 92.995 -52.875 93.325 ;
        RECT -53.205 91.635 -52.875 91.965 ;
        RECT -53.205 90.275 -52.875 90.605 ;
        RECT -53.205 88.915 -52.875 89.245 ;
        RECT -53.205 87.555 -52.875 87.885 ;
        RECT -53.205 86.195 -52.875 86.525 ;
        RECT -53.205 84.835 -52.875 85.165 ;
        RECT -53.205 83.475 -52.875 83.805 ;
        RECT -53.205 82.115 -52.875 82.445 ;
        RECT -53.205 80.755 -52.875 81.085 ;
        RECT -53.205 79.395 -52.875 79.725 ;
        RECT -53.205 78.035 -52.875 78.365 ;
        RECT -53.205 76.675 -52.875 77.005 ;
        RECT -53.205 75.315 -52.875 75.645 ;
        RECT -53.205 73.955 -52.875 74.285 ;
        RECT -53.205 71.64 -52.875 71.97 ;
        RECT -53.205 69.465 -52.875 69.795 ;
        RECT -53.205 68.615 -52.875 68.945 ;
        RECT -53.205 66.305 -52.875 66.635 ;
        RECT -53.205 65.455 -52.875 65.785 ;
        RECT -53.205 63.145 -52.875 63.475 ;
        RECT -53.205 62.295 -52.875 62.625 ;
        RECT -53.205 59.985 -52.875 60.315 ;
        RECT -53.205 59.135 -52.875 59.465 ;
        RECT -53.205 56.825 -52.875 57.155 ;
        RECT -53.205 55.975 -52.875 56.305 ;
        RECT -53.205 53.665 -52.875 53.995 ;
        RECT -53.205 52.815 -52.875 53.145 ;
        RECT -53.205 50.64 -52.875 50.97 ;
        RECT -53.205 48.115 -52.875 48.445 ;
        RECT -53.205 46.755 -52.875 47.085 ;
        RECT -53.205 45.395 -52.875 45.725 ;
        RECT -53.205 44.035 -52.875 44.365 ;
        RECT -53.205 42.675 -52.875 43.005 ;
        RECT -53.205 41.315 -52.875 41.645 ;
        RECT -53.205 39.955 -52.875 40.285 ;
        RECT -53.205 38.595 -52.875 38.925 ;
        RECT -53.205 37.235 -52.875 37.565 ;
        RECT -53.205 35.875 -52.875 36.205 ;
        RECT -53.205 34.515 -52.875 34.845 ;
        RECT -53.205 33.155 -52.875 33.485 ;
        RECT -53.205 31.795 -52.875 32.125 ;
        RECT -53.205 30.435 -52.875 30.765 ;
        RECT -53.205 29.075 -52.875 29.405 ;
        RECT -53.205 27.715 -52.875 28.045 ;
        RECT -53.205 26.355 -52.875 26.685 ;
        RECT -53.205 24.995 -52.875 25.325 ;
        RECT -53.205 23.635 -52.875 23.965 ;
        RECT -53.205 22.275 -52.875 22.605 ;
        RECT -53.205 20.915 -52.875 21.245 ;
        RECT -53.205 19.555 -52.875 19.885 ;
        RECT -53.205 18.195 -52.875 18.525 ;
        RECT -53.205 16.835 -52.875 17.165 ;
        RECT -53.205 15.475 -52.875 15.805 ;
        RECT -53.205 14.115 -52.875 14.445 ;
        RECT -53.205 12.755 -52.875 13.085 ;
        RECT -53.205 11.395 -52.875 11.725 ;
        RECT -53.205 10.035 -52.875 10.365 ;
        RECT -53.205 8.675 -52.875 9.005 ;
        RECT -53.205 7.315 -52.875 7.645 ;
        RECT -53.205 5.955 -52.875 6.285 ;
        RECT -53.205 4.595 -52.875 4.925 ;
        RECT -53.205 3.235 -52.875 3.565 ;
        RECT -53.205 1.875 -52.875 2.205 ;
        RECT -53.205 0.515 -52.875 0.845 ;
        RECT -53.205 -0.845 -52.875 -0.515 ;
        RECT -53.205 -2.205 -52.875 -1.875 ;
        RECT -53.205 -3.565 -52.875 -3.235 ;
        RECT -53.205 -4.925 -52.875 -4.595 ;
        RECT -53.205 -6.285 -52.875 -5.955 ;
        RECT -53.205 -7.645 -52.875 -7.315 ;
        RECT -53.205 -9.005 -52.875 -8.675 ;
        RECT -53.205 -10.365 -52.875 -10.035 ;
        RECT -53.205 -11.725 -52.875 -11.395 ;
        RECT -53.205 -13.085 -52.875 -12.755 ;
        RECT -53.205 -14.445 -52.875 -14.115 ;
        RECT -53.205 -15.805 -52.875 -15.475 ;
        RECT -53.205 -17.165 -52.875 -16.835 ;
        RECT -53.205 -18.525 -52.875 -18.195 ;
        RECT -53.205 -19.885 -52.875 -19.555 ;
        RECT -53.205 -21.245 -52.875 -20.915 ;
        RECT -53.205 -22.605 -52.875 -22.275 ;
        RECT -53.205 -23.965 -52.875 -23.635 ;
        RECT -53.205 -25.325 -52.875 -24.995 ;
        RECT -53.205 -26.685 -52.875 -26.355 ;
        RECT -53.205 -28.045 -52.875 -27.715 ;
        RECT -53.205 -29.405 -52.875 -29.075 ;
        RECT -53.205 -30.765 -52.875 -30.435 ;
        RECT -53.205 -32.125 -52.875 -31.795 ;
        RECT -53.205 -33.485 -52.875 -33.155 ;
        RECT -53.205 -34.845 -52.875 -34.515 ;
        RECT -53.205 -37.565 -52.875 -37.235 ;
        RECT -53.205 -38.925 -52.875 -38.595 ;
        RECT -53.205 -40.285 -52.875 -39.955 ;
        RECT -53.205 -41.645 -52.875 -41.315 ;
        RECT -53.205 -43.005 -52.875 -42.675 ;
        RECT -53.205 -44.365 -52.875 -44.035 ;
        RECT -53.205 -45.725 -52.875 -45.395 ;
        RECT -53.205 -47.085 -52.875 -46.755 ;
        RECT -53.205 -48.445 -52.875 -48.115 ;
        RECT -53.205 -49.805 -52.875 -49.475 ;
        RECT -53.205 -51.165 -52.875 -50.835 ;
        RECT -53.205 -52.525 -52.875 -52.195 ;
        RECT -53.205 -53.885 -52.875 -53.555 ;
        RECT -53.205 -55.245 -52.875 -54.915 ;
        RECT -53.205 -56.605 -52.875 -56.275 ;
        RECT -53.205 -57.965 -52.875 -57.635 ;
        RECT -53.205 -59.325 -52.875 -58.995 ;
        RECT -53.205 -60.685 -52.875 -60.355 ;
        RECT -53.205 -62.045 -52.875 -61.715 ;
        RECT -53.205 -63.405 -52.875 -63.075 ;
        RECT -53.205 -64.765 -52.875 -64.435 ;
        RECT -53.205 -66.125 -52.875 -65.795 ;
        RECT -53.205 -67.485 -52.875 -67.155 ;
        RECT -53.205 -68.845 -52.875 -68.515 ;
        RECT -53.205 -70.205 -52.875 -69.875 ;
        RECT -53.205 -71.565 -52.875 -71.235 ;
        RECT -53.205 -72.925 -52.875 -72.595 ;
        RECT -53.205 -74.285 -52.875 -73.955 ;
        RECT -53.205 -75.645 -52.875 -75.315 ;
        RECT -53.205 -77.005 -52.875 -76.675 ;
        RECT -53.205 -78.365 -52.875 -78.035 ;
        RECT -53.205 -79.725 -52.875 -79.395 ;
        RECT -53.205 -81.085 -52.875 -80.755 ;
        RECT -53.205 -82.445 -52.875 -82.115 ;
        RECT -53.205 -83.805 -52.875 -83.475 ;
        RECT -53.205 -85.165 -52.875 -84.835 ;
        RECT -53.205 -86.525 -52.875 -86.195 ;
        RECT -53.205 -87.885 -52.875 -87.555 ;
        RECT -53.205 -89.245 -52.875 -88.915 ;
        RECT -53.205 -90.605 -52.875 -90.275 ;
        RECT -53.205 -91.965 -52.875 -91.635 ;
        RECT -53.205 -93.325 -52.875 -92.995 ;
        RECT -53.205 -94.685 -52.875 -94.355 ;
        RECT -53.205 -96.045 -52.875 -95.715 ;
        RECT -53.205 -97.405 -52.875 -97.075 ;
        RECT -53.205 -98.765 -52.875 -98.435 ;
        RECT -53.205 -100.125 -52.875 -99.795 ;
        RECT -53.205 -101.485 -52.875 -101.155 ;
        RECT -53.205 -102.845 -52.875 -102.515 ;
        RECT -53.205 -104.205 -52.875 -103.875 ;
        RECT -53.205 -105.565 -52.875 -105.235 ;
        RECT -53.205 -106.925 -52.875 -106.595 ;
        RECT -53.205 -108.285 -52.875 -107.955 ;
        RECT -53.205 -109.645 -52.875 -109.315 ;
        RECT -53.205 -111.005 -52.875 -110.675 ;
        RECT -53.205 -111.87 -52.875 -111.54 ;
        RECT -53.205 -113.725 -52.875 -113.395 ;
        RECT -53.205 -115.085 -52.875 -114.755 ;
        RECT -53.205 -116.445 -52.875 -116.115 ;
        RECT -53.205 -117.805 -52.875 -117.475 ;
        RECT -53.205 -120.525 -52.875 -120.195 ;
        RECT -53.205 -121.885 -52.875 -121.555 ;
        RECT -53.205 -123.245 -52.875 -122.915 ;
        RECT -53.205 -124.71 -52.875 -124.38 ;
        RECT -53.205 -125.965 -52.875 -125.635 ;
        RECT -53.205 -127.325 -52.875 -126.995 ;
        RECT -53.205 -130.045 -52.875 -129.715 ;
        RECT -53.2 -132.08 -52.88 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.205 -211.645 -52.875 -211.315 ;
        RECT -53.205 -214.365 -52.875 -214.035 ;
        RECT -53.205 -215.725 -52.875 -215.395 ;
        RECT -53.205 -217.085 -52.875 -216.755 ;
        RECT -53.205 -218.445 -52.875 -218.115 ;
        RECT -53.205 -224.09 -52.875 -222.96 ;
        RECT -53.2 -224.205 -52.88 -210.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -51.845 132.52 -51.515 133.65 ;
        RECT -51.845 128.355 -51.515 128.685 ;
        RECT -51.845 126.995 -51.515 127.325 ;
        RECT -51.845 125.635 -51.515 125.965 ;
        RECT -51.845 124.275 -51.515 124.605 ;
        RECT -51.845 122.915 -51.515 123.245 ;
        RECT -51.845 121.555 -51.515 121.885 ;
        RECT -51.845 120.195 -51.515 120.525 ;
        RECT -51.845 118.835 -51.515 119.165 ;
        RECT -51.845 117.475 -51.515 117.805 ;
        RECT -51.845 116.115 -51.515 116.445 ;
        RECT -51.845 114.755 -51.515 115.085 ;
        RECT -51.845 113.395 -51.515 113.725 ;
        RECT -51.845 112.035 -51.515 112.365 ;
        RECT -51.845 110.675 -51.515 111.005 ;
        RECT -51.845 109.315 -51.515 109.645 ;
        RECT -51.845 107.955 -51.515 108.285 ;
        RECT -51.845 106.595 -51.515 106.925 ;
        RECT -51.845 105.235 -51.515 105.565 ;
        RECT -51.845 103.875 -51.515 104.205 ;
        RECT -51.845 102.515 -51.515 102.845 ;
        RECT -51.845 101.155 -51.515 101.485 ;
        RECT -51.845 99.795 -51.515 100.125 ;
        RECT -51.845 98.435 -51.515 98.765 ;
        RECT -51.845 97.075 -51.515 97.405 ;
        RECT -51.845 95.715 -51.515 96.045 ;
        RECT -51.845 94.355 -51.515 94.685 ;
        RECT -51.845 92.995 -51.515 93.325 ;
        RECT -51.845 91.635 -51.515 91.965 ;
        RECT -51.845 90.275 -51.515 90.605 ;
        RECT -51.845 88.915 -51.515 89.245 ;
        RECT -51.845 87.555 -51.515 87.885 ;
        RECT -51.845 86.195 -51.515 86.525 ;
        RECT -51.845 84.835 -51.515 85.165 ;
        RECT -51.845 83.475 -51.515 83.805 ;
        RECT -51.845 82.115 -51.515 82.445 ;
        RECT -51.845 80.755 -51.515 81.085 ;
        RECT -51.845 79.395 -51.515 79.725 ;
        RECT -51.845 78.035 -51.515 78.365 ;
        RECT -51.845 76.675 -51.515 77.005 ;
        RECT -51.845 75.315 -51.515 75.645 ;
        RECT -51.845 73.955 -51.515 74.285 ;
        RECT -51.845 71.64 -51.515 71.97 ;
        RECT -51.845 69.465 -51.515 69.795 ;
        RECT -51.845 68.615 -51.515 68.945 ;
        RECT -51.845 66.305 -51.515 66.635 ;
        RECT -51.845 65.455 -51.515 65.785 ;
        RECT -51.845 63.145 -51.515 63.475 ;
        RECT -51.845 62.295 -51.515 62.625 ;
        RECT -51.845 59.985 -51.515 60.315 ;
        RECT -51.845 59.135 -51.515 59.465 ;
        RECT -51.845 56.825 -51.515 57.155 ;
        RECT -51.845 55.975 -51.515 56.305 ;
        RECT -51.845 53.665 -51.515 53.995 ;
        RECT -51.845 52.815 -51.515 53.145 ;
        RECT -51.845 50.64 -51.515 50.97 ;
        RECT -51.845 48.115 -51.515 48.445 ;
        RECT -51.845 46.755 -51.515 47.085 ;
        RECT -51.845 45.395 -51.515 45.725 ;
        RECT -51.845 44.035 -51.515 44.365 ;
        RECT -51.845 42.675 -51.515 43.005 ;
        RECT -51.845 41.315 -51.515 41.645 ;
        RECT -51.845 39.955 -51.515 40.285 ;
        RECT -51.845 38.595 -51.515 38.925 ;
        RECT -51.84 38.595 -51.52 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -51.845 -11.725 -51.515 -11.395 ;
        RECT -51.845 -13.085 -51.515 -12.755 ;
        RECT -51.845 -14.445 -51.515 -14.115 ;
        RECT -51.845 -15.805 -51.515 -15.475 ;
        RECT -51.845 -17.165 -51.515 -16.835 ;
        RECT -51.845 -18.525 -51.515 -18.195 ;
        RECT -51.845 -19.885 -51.515 -19.555 ;
        RECT -51.845 -21.245 -51.515 -20.915 ;
        RECT -51.845 -22.605 -51.515 -22.275 ;
        RECT -51.845 -23.965 -51.515 -23.635 ;
        RECT -51.845 -25.325 -51.515 -24.995 ;
        RECT -51.845 -26.685 -51.515 -26.355 ;
        RECT -51.845 -28.045 -51.515 -27.715 ;
        RECT -51.845 -29.405 -51.515 -29.075 ;
        RECT -51.845 -30.765 -51.515 -30.435 ;
        RECT -51.845 -32.125 -51.515 -31.795 ;
        RECT -51.845 -33.485 -51.515 -33.155 ;
        RECT -51.845 -34.845 -51.515 -34.515 ;
        RECT -51.845 -37.565 -51.515 -37.235 ;
        RECT -51.845 -38.925 -51.515 -38.595 ;
        RECT -51.845 -40.285 -51.515 -39.955 ;
        RECT -51.845 -41.645 -51.515 -41.315 ;
        RECT -51.845 -43.005 -51.515 -42.675 ;
        RECT -51.845 -44.365 -51.515 -44.035 ;
        RECT -51.845 -45.725 -51.515 -45.395 ;
        RECT -51.845 -47.085 -51.515 -46.755 ;
        RECT -51.845 -48.445 -51.515 -48.115 ;
        RECT -51.845 -49.805 -51.515 -49.475 ;
        RECT -51.845 -51.165 -51.515 -50.835 ;
        RECT -51.845 -52.525 -51.515 -52.195 ;
        RECT -51.845 -53.885 -51.515 -53.555 ;
        RECT -51.845 -55.245 -51.515 -54.915 ;
        RECT -51.845 -56.605 -51.515 -56.275 ;
        RECT -51.845 -57.965 -51.515 -57.635 ;
        RECT -51.845 -59.325 -51.515 -58.995 ;
        RECT -51.845 -60.685 -51.515 -60.355 ;
        RECT -51.845 -62.045 -51.515 -61.715 ;
        RECT -51.845 -63.405 -51.515 -63.075 ;
        RECT -51.845 -64.765 -51.515 -64.435 ;
        RECT -51.845 -66.125 -51.515 -65.795 ;
        RECT -51.845 -67.485 -51.515 -67.155 ;
        RECT -51.845 -68.845 -51.515 -68.515 ;
        RECT -51.845 -70.205 -51.515 -69.875 ;
        RECT -51.845 -71.565 -51.515 -71.235 ;
        RECT -51.845 -72.925 -51.515 -72.595 ;
        RECT -51.845 -74.285 -51.515 -73.955 ;
        RECT -51.845 -75.645 -51.515 -75.315 ;
        RECT -51.845 -77.005 -51.515 -76.675 ;
        RECT -51.845 -78.365 -51.515 -78.035 ;
        RECT -51.845 -79.725 -51.515 -79.395 ;
        RECT -51.845 -81.085 -51.515 -80.755 ;
        RECT -51.845 -82.445 -51.515 -82.115 ;
        RECT -51.845 -83.805 -51.515 -83.475 ;
        RECT -51.845 -85.165 -51.515 -84.835 ;
        RECT -51.845 -86.525 -51.515 -86.195 ;
        RECT -51.845 -87.885 -51.515 -87.555 ;
        RECT -51.845 -89.245 -51.515 -88.915 ;
        RECT -51.845 -90.605 -51.515 -90.275 ;
        RECT -51.845 -91.965 -51.515 -91.635 ;
        RECT -51.845 -93.325 -51.515 -92.995 ;
        RECT -51.845 -94.685 -51.515 -94.355 ;
        RECT -51.845 -96.045 -51.515 -95.715 ;
        RECT -51.845 -97.405 -51.515 -97.075 ;
        RECT -51.845 -98.765 -51.515 -98.435 ;
        RECT -51.845 -100.125 -51.515 -99.795 ;
        RECT -51.845 -101.485 -51.515 -101.155 ;
        RECT -51.845 -102.845 -51.515 -102.515 ;
        RECT -51.845 -104.205 -51.515 -103.875 ;
        RECT -51.845 -105.565 -51.515 -105.235 ;
        RECT -51.845 -106.925 -51.515 -106.595 ;
        RECT -51.845 -108.285 -51.515 -107.955 ;
        RECT -51.845 -109.645 -51.515 -109.315 ;
        RECT -51.845 -111.005 -51.515 -110.675 ;
        RECT -51.845 -111.87 -51.515 -111.54 ;
        RECT -51.845 -113.725 -51.515 -113.395 ;
        RECT -51.845 -115.085 -51.515 -114.755 ;
        RECT -51.845 -116.445 -51.515 -116.115 ;
        RECT -51.845 -117.805 -51.515 -117.475 ;
        RECT -51.845 -120.525 -51.515 -120.195 ;
        RECT -51.845 -121.885 -51.515 -121.555 ;
        RECT -51.845 -123.245 -51.515 -122.915 ;
        RECT -51.845 -124.71 -51.515 -124.38 ;
        RECT -51.845 -125.965 -51.515 -125.635 ;
        RECT -51.845 -127.325 -51.515 -126.995 ;
        RECT -51.845 -130.045 -51.515 -129.715 ;
        RECT -51.845 -135.485 -51.515 -135.155 ;
        RECT -51.845 -136.845 -51.515 -136.515 ;
        RECT -51.845 -138.205 -51.515 -137.875 ;
        RECT -51.845 -139.565 -51.515 -139.235 ;
        RECT -51.845 -142.285 -51.515 -141.955 ;
        RECT -51.845 -143.645 -51.515 -143.315 ;
        RECT -51.845 -145.005 -51.515 -144.675 ;
        RECT -51.845 -146.365 -51.515 -146.035 ;
        RECT -51.845 -147.725 -51.515 -147.395 ;
        RECT -51.845 -149.085 -51.515 -148.755 ;
        RECT -51.845 -150.445 -51.515 -150.115 ;
        RECT -51.845 -151.805 -51.515 -151.475 ;
        RECT -51.845 -153.165 -51.515 -152.835 ;
        RECT -51.845 -154.525 -51.515 -154.195 ;
        RECT -51.845 -155.885 -51.515 -155.555 ;
        RECT -51.845 -157.245 -51.515 -156.915 ;
        RECT -51.845 -158.605 -51.515 -158.275 ;
        RECT -51.845 -159.965 -51.515 -159.635 ;
        RECT -51.845 -161.325 -51.515 -160.995 ;
        RECT -51.845 -162.685 -51.515 -162.355 ;
        RECT -51.845 -164.045 -51.515 -163.715 ;
        RECT -51.845 -165.405 -51.515 -165.075 ;
        RECT -51.845 -166.765 -51.515 -166.435 ;
        RECT -51.845 -168.125 -51.515 -167.795 ;
        RECT -51.845 -169.485 -51.515 -169.155 ;
        RECT -51.845 -170.845 -51.515 -170.515 ;
        RECT -51.845 -172.205 -51.515 -171.875 ;
        RECT -51.845 -173.565 -51.515 -173.235 ;
        RECT -51.845 -174.925 -51.515 -174.595 ;
        RECT -51.845 -176.285 -51.515 -175.955 ;
        RECT -51.845 -177.645 -51.515 -177.315 ;
        RECT -51.845 -179.005 -51.515 -178.675 ;
        RECT -51.845 -180.365 -51.515 -180.035 ;
        RECT -51.845 -181.725 -51.515 -181.395 ;
        RECT -51.845 -183.085 -51.515 -182.755 ;
        RECT -51.845 -184.445 -51.515 -184.115 ;
        RECT -51.845 -185.805 -51.515 -185.475 ;
        RECT -51.845 -187.165 -51.515 -186.835 ;
        RECT -51.845 -188.525 -51.515 -188.195 ;
        RECT -51.845 -189.885 -51.515 -189.555 ;
        RECT -51.845 -191.245 -51.515 -190.915 ;
        RECT -51.845 -192.605 -51.515 -192.275 ;
        RECT -51.845 -193.965 -51.515 -193.635 ;
        RECT -51.845 -195.325 -51.515 -194.995 ;
        RECT -51.845 -196.685 -51.515 -196.355 ;
        RECT -51.845 -198.045 -51.515 -197.715 ;
        RECT -51.845 -199.405 -51.515 -199.075 ;
        RECT -51.845 -200.765 -51.515 -200.435 ;
        RECT -51.845 -202.125 -51.515 -201.795 ;
        RECT -51.845 -203.485 -51.515 -203.155 ;
        RECT -51.845 -204.845 -51.515 -204.515 ;
        RECT -51.845 -206.555 -51.515 -206.225 ;
        RECT -51.845 -207.565 -51.515 -207.235 ;
        RECT -51.845 -208.925 -51.515 -208.595 ;
        RECT -51.845 -211.645 -51.515 -211.315 ;
        RECT -51.845 -214.365 -51.515 -214.035 ;
        RECT -51.845 -215.725 -51.515 -215.395 ;
        RECT -51.845 -217.085 -51.515 -216.755 ;
        RECT -51.845 -218.445 -51.515 -218.115 ;
        RECT -51.845 -224.09 -51.515 -222.96 ;
        RECT -51.84 -224.205 -51.52 -10.72 ;
    END
    PORT
      LAYER met3 ;
        RECT -50.485 132.52 -50.155 133.65 ;
        RECT -50.485 128.355 -50.155 128.685 ;
        RECT -50.485 126.995 -50.155 127.325 ;
        RECT -50.485 125.635 -50.155 125.965 ;
        RECT -50.485 124.275 -50.155 124.605 ;
        RECT -50.485 122.915 -50.155 123.245 ;
        RECT -50.485 121.555 -50.155 121.885 ;
        RECT -50.485 120.195 -50.155 120.525 ;
        RECT -50.485 118.835 -50.155 119.165 ;
        RECT -50.485 117.475 -50.155 117.805 ;
        RECT -50.485 116.115 -50.155 116.445 ;
        RECT -50.485 114.755 -50.155 115.085 ;
        RECT -50.485 113.395 -50.155 113.725 ;
        RECT -50.485 112.035 -50.155 112.365 ;
        RECT -50.485 110.675 -50.155 111.005 ;
        RECT -50.485 109.315 -50.155 109.645 ;
        RECT -50.485 107.955 -50.155 108.285 ;
        RECT -50.485 106.595 -50.155 106.925 ;
        RECT -50.485 105.235 -50.155 105.565 ;
        RECT -50.485 103.875 -50.155 104.205 ;
        RECT -50.485 102.515 -50.155 102.845 ;
        RECT -50.485 101.155 -50.155 101.485 ;
        RECT -50.485 99.795 -50.155 100.125 ;
        RECT -50.485 98.435 -50.155 98.765 ;
        RECT -50.485 97.075 -50.155 97.405 ;
        RECT -50.485 95.715 -50.155 96.045 ;
        RECT -50.485 94.355 -50.155 94.685 ;
        RECT -50.485 92.995 -50.155 93.325 ;
        RECT -50.485 91.635 -50.155 91.965 ;
        RECT -50.485 90.275 -50.155 90.605 ;
        RECT -50.485 88.915 -50.155 89.245 ;
        RECT -50.485 87.555 -50.155 87.885 ;
        RECT -50.485 86.195 -50.155 86.525 ;
        RECT -50.485 84.835 -50.155 85.165 ;
        RECT -50.485 83.475 -50.155 83.805 ;
        RECT -50.485 82.115 -50.155 82.445 ;
        RECT -50.485 80.755 -50.155 81.085 ;
        RECT -50.485 79.395 -50.155 79.725 ;
        RECT -50.485 78.035 -50.155 78.365 ;
        RECT -50.485 76.675 -50.155 77.005 ;
        RECT -50.485 75.315 -50.155 75.645 ;
        RECT -50.485 73.955 -50.155 74.285 ;
        RECT -50.48 73.28 -50.16 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -50.485 48.115 -50.155 48.445 ;
        RECT -50.485 46.755 -50.155 47.085 ;
        RECT -50.485 45.395 -50.155 45.725 ;
        RECT -50.485 44.035 -50.155 44.365 ;
        RECT -50.485 39.955 -50.155 40.285 ;
        RECT -50.485 38.595 -50.155 38.925 ;
        RECT -50.485 35.875 -50.155 36.205 ;
        RECT -50.485 34.515 -50.155 34.845 ;
        RECT -50.485 33.155 -50.155 33.485 ;
        RECT -50.485 31.795 -50.155 32.125 ;
        RECT -50.485 30.435 -50.155 30.765 ;
        RECT -50.485 29.075 -50.155 29.405 ;
        RECT -50.485 27.715 -50.155 28.045 ;
        RECT -50.485 26.355 -50.155 26.685 ;
        RECT -50.485 24.995 -50.155 25.325 ;
        RECT -50.485 23.635 -50.155 23.965 ;
        RECT -50.485 22.275 -50.155 22.605 ;
        RECT -50.485 20.915 -50.155 21.245 ;
        RECT -50.485 19.555 -50.155 19.885 ;
        RECT -50.485 18.195 -50.155 18.525 ;
        RECT -50.485 16.835 -50.155 17.165 ;
        RECT -50.485 15.475 -50.155 15.805 ;
        RECT -50.485 14.115 -50.155 14.445 ;
        RECT -50.485 12.755 -50.155 13.085 ;
        RECT -50.485 11.395 -50.155 11.725 ;
        RECT -50.485 10.035 -50.155 10.365 ;
        RECT -50.485 8.675 -50.155 9.005 ;
        RECT -50.485 7.315 -50.155 7.645 ;
        RECT -50.485 5.955 -50.155 6.285 ;
        RECT -50.485 4.595 -50.155 4.925 ;
        RECT -50.485 3.235 -50.155 3.565 ;
        RECT -50.485 1.875 -50.155 2.205 ;
        RECT -50.485 0.515 -50.155 0.845 ;
        RECT -50.485 -0.845 -50.155 -0.515 ;
        RECT -50.485 -2.205 -50.155 -1.875 ;
        RECT -50.485 -3.565 -50.155 -3.235 ;
        RECT -50.485 -4.925 -50.155 -4.595 ;
        RECT -50.485 -6.285 -50.155 -5.955 ;
        RECT -50.485 -7.645 -50.155 -7.315 ;
        RECT -50.485 -9.005 -50.155 -8.675 ;
        RECT -50.485 -11.725 -50.155 -11.395 ;
        RECT -50.485 -13.085 -50.155 -12.755 ;
        RECT -50.485 -14.445 -50.155 -14.115 ;
        RECT -50.485 -15.805 -50.155 -15.475 ;
        RECT -50.485 -17.165 -50.155 -16.835 ;
        RECT -50.485 -18.525 -50.155 -18.195 ;
        RECT -50.485 -19.885 -50.155 -19.555 ;
        RECT -50.485 -21.245 -50.155 -20.915 ;
        RECT -50.485 -22.605 -50.155 -22.275 ;
        RECT -50.485 -23.965 -50.155 -23.635 ;
        RECT -50.485 -25.325 -50.155 -24.995 ;
        RECT -50.485 -26.685 -50.155 -26.355 ;
        RECT -50.485 -28.045 -50.155 -27.715 ;
        RECT -50.485 -29.405 -50.155 -29.075 ;
        RECT -50.485 -30.765 -50.155 -30.435 ;
        RECT -50.485 -32.125 -50.155 -31.795 ;
        RECT -50.485 -33.485 -50.155 -33.155 ;
        RECT -50.485 -34.845 -50.155 -34.515 ;
        RECT -50.485 -37.565 -50.155 -37.235 ;
        RECT -50.485 -38.925 -50.155 -38.595 ;
        RECT -50.485 -40.285 -50.155 -39.955 ;
        RECT -50.485 -41.645 -50.155 -41.315 ;
        RECT -50.485 -43.005 -50.155 -42.675 ;
        RECT -50.485 -44.365 -50.155 -44.035 ;
        RECT -50.485 -45.725 -50.155 -45.395 ;
        RECT -50.485 -47.085 -50.155 -46.755 ;
        RECT -50.485 -48.445 -50.155 -48.115 ;
        RECT -50.485 -49.805 -50.155 -49.475 ;
        RECT -50.485 -51.165 -50.155 -50.835 ;
        RECT -50.485 -52.525 -50.155 -52.195 ;
        RECT -50.485 -53.885 -50.155 -53.555 ;
        RECT -50.485 -55.245 -50.155 -54.915 ;
        RECT -50.485 -56.605 -50.155 -56.275 ;
        RECT -50.485 -57.965 -50.155 -57.635 ;
        RECT -50.485 -59.325 -50.155 -58.995 ;
        RECT -50.485 -60.685 -50.155 -60.355 ;
        RECT -50.485 -62.045 -50.155 -61.715 ;
        RECT -50.485 -63.405 -50.155 -63.075 ;
        RECT -50.485 -64.765 -50.155 -64.435 ;
        RECT -50.485 -66.125 -50.155 -65.795 ;
        RECT -50.485 -67.485 -50.155 -67.155 ;
        RECT -50.485 -68.845 -50.155 -68.515 ;
        RECT -50.485 -70.205 -50.155 -69.875 ;
        RECT -50.485 -71.565 -50.155 -71.235 ;
        RECT -50.485 -72.925 -50.155 -72.595 ;
        RECT -50.485 -74.285 -50.155 -73.955 ;
        RECT -50.485 -75.645 -50.155 -75.315 ;
        RECT -50.485 -77.005 -50.155 -76.675 ;
        RECT -50.485 -78.365 -50.155 -78.035 ;
        RECT -50.485 -79.725 -50.155 -79.395 ;
        RECT -50.485 -81.085 -50.155 -80.755 ;
        RECT -50.485 -82.445 -50.155 -82.115 ;
        RECT -50.485 -83.805 -50.155 -83.475 ;
        RECT -50.485 -85.165 -50.155 -84.835 ;
        RECT -50.485 -86.525 -50.155 -86.195 ;
        RECT -50.485 -87.885 -50.155 -87.555 ;
        RECT -50.485 -89.245 -50.155 -88.915 ;
        RECT -50.485 -90.605 -50.155 -90.275 ;
        RECT -50.485 -91.965 -50.155 -91.635 ;
        RECT -50.485 -93.325 -50.155 -92.995 ;
        RECT -50.485 -94.685 -50.155 -94.355 ;
        RECT -50.485 -96.045 -50.155 -95.715 ;
        RECT -50.485 -97.405 -50.155 -97.075 ;
        RECT -50.485 -98.765 -50.155 -98.435 ;
        RECT -50.485 -100.125 -50.155 -99.795 ;
        RECT -50.485 -101.485 -50.155 -101.155 ;
        RECT -50.485 -102.845 -50.155 -102.515 ;
        RECT -50.485 -104.205 -50.155 -103.875 ;
        RECT -50.485 -105.565 -50.155 -105.235 ;
        RECT -50.485 -106.925 -50.155 -106.595 ;
        RECT -50.485 -108.285 -50.155 -107.955 ;
        RECT -50.485 -109.645 -50.155 -109.315 ;
        RECT -50.485 -111.005 -50.155 -110.675 ;
        RECT -50.485 -111.87 -50.155 -111.54 ;
        RECT -50.485 -113.725 -50.155 -113.395 ;
        RECT -50.485 -115.085 -50.155 -114.755 ;
        RECT -50.485 -116.445 -50.155 -116.115 ;
        RECT -50.485 -117.805 -50.155 -117.475 ;
        RECT -50.485 -120.525 -50.155 -120.195 ;
        RECT -50.485 -121.885 -50.155 -121.555 ;
        RECT -50.485 -123.245 -50.155 -122.915 ;
        RECT -50.485 -124.71 -50.155 -124.38 ;
        RECT -50.485 -125.965 -50.155 -125.635 ;
        RECT -50.485 -127.325 -50.155 -126.995 ;
        RECT -50.485 -130.045 -50.155 -129.715 ;
        RECT -50.485 -135.485 -50.155 -135.155 ;
        RECT -50.485 -136.845 -50.155 -136.515 ;
        RECT -50.485 -138.205 -50.155 -137.875 ;
        RECT -50.485 -139.565 -50.155 -139.235 ;
        RECT -50.485 -142.285 -50.155 -141.955 ;
        RECT -50.485 -143.645 -50.155 -143.315 ;
        RECT -50.485 -145.005 -50.155 -144.675 ;
        RECT -50.485 -146.365 -50.155 -146.035 ;
        RECT -50.485 -147.725 -50.155 -147.395 ;
        RECT -50.485 -149.085 -50.155 -148.755 ;
        RECT -50.485 -150.445 -50.155 -150.115 ;
        RECT -50.485 -151.805 -50.155 -151.475 ;
        RECT -50.485 -153.165 -50.155 -152.835 ;
        RECT -50.485 -154.525 -50.155 -154.195 ;
        RECT -50.485 -155.885 -50.155 -155.555 ;
        RECT -50.485 -157.245 -50.155 -156.915 ;
        RECT -50.485 -158.605 -50.155 -158.275 ;
        RECT -50.485 -159.965 -50.155 -159.635 ;
        RECT -50.485 -161.325 -50.155 -160.995 ;
        RECT -50.485 -162.685 -50.155 -162.355 ;
        RECT -50.485 -164.045 -50.155 -163.715 ;
        RECT -50.485 -165.405 -50.155 -165.075 ;
        RECT -50.485 -166.765 -50.155 -166.435 ;
        RECT -50.485 -168.125 -50.155 -167.795 ;
        RECT -50.485 -169.485 -50.155 -169.155 ;
        RECT -50.485 -170.845 -50.155 -170.515 ;
        RECT -50.485 -172.205 -50.155 -171.875 ;
        RECT -50.485 -173.565 -50.155 -173.235 ;
        RECT -50.485 -174.925 -50.155 -174.595 ;
        RECT -50.485 -176.285 -50.155 -175.955 ;
        RECT -50.485 -177.645 -50.155 -177.315 ;
        RECT -50.485 -179.005 -50.155 -178.675 ;
        RECT -50.485 -180.365 -50.155 -180.035 ;
        RECT -50.485 -181.725 -50.155 -181.395 ;
        RECT -50.485 -183.085 -50.155 -182.755 ;
        RECT -50.485 -184.445 -50.155 -184.115 ;
        RECT -50.485 -185.805 -50.155 -185.475 ;
        RECT -50.485 -187.165 -50.155 -186.835 ;
        RECT -50.485 -188.525 -50.155 -188.195 ;
        RECT -50.485 -189.885 -50.155 -189.555 ;
        RECT -50.485 -191.245 -50.155 -190.915 ;
        RECT -50.485 -192.605 -50.155 -192.275 ;
        RECT -50.485 -193.965 -50.155 -193.635 ;
        RECT -50.485 -195.325 -50.155 -194.995 ;
        RECT -50.485 -196.685 -50.155 -196.355 ;
        RECT -50.485 -198.045 -50.155 -197.715 ;
        RECT -50.485 -199.405 -50.155 -199.075 ;
        RECT -50.485 -200.765 -50.155 -200.435 ;
        RECT -50.485 -202.125 -50.155 -201.795 ;
        RECT -50.485 -203.485 -50.155 -203.155 ;
        RECT -50.485 -204.845 -50.155 -204.515 ;
        RECT -50.485 -206.555 -50.155 -206.225 ;
        RECT -50.485 -207.565 -50.155 -207.235 ;
        RECT -50.485 -208.925 -50.155 -208.595 ;
        RECT -50.485 -210.285 -50.155 -209.955 ;
        RECT -50.485 -211.645 -50.155 -211.315 ;
        RECT -50.485 -214.365 -50.155 -214.035 ;
        RECT -50.485 -215.725 -50.155 -215.395 ;
        RECT -50.485 -217.085 -50.155 -216.755 ;
        RECT -50.485 -218.445 -50.155 -218.115 ;
        RECT -50.485 -224.09 -50.155 -222.96 ;
        RECT -50.48 -224.205 -50.16 49.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.125 132.52 -48.795 133.65 ;
        RECT -49.125 128.355 -48.795 128.685 ;
        RECT -49.125 126.995 -48.795 127.325 ;
        RECT -49.125 125.635 -48.795 125.965 ;
        RECT -49.125 124.275 -48.795 124.605 ;
        RECT -49.125 122.915 -48.795 123.245 ;
        RECT -49.125 121.555 -48.795 121.885 ;
        RECT -49.125 120.195 -48.795 120.525 ;
        RECT -49.125 118.835 -48.795 119.165 ;
        RECT -49.125 117.475 -48.795 117.805 ;
        RECT -49.125 116.115 -48.795 116.445 ;
        RECT -49.125 114.755 -48.795 115.085 ;
        RECT -49.125 113.395 -48.795 113.725 ;
        RECT -49.125 112.035 -48.795 112.365 ;
        RECT -49.125 110.675 -48.795 111.005 ;
        RECT -49.125 109.315 -48.795 109.645 ;
        RECT -49.125 107.955 -48.795 108.285 ;
        RECT -49.125 106.595 -48.795 106.925 ;
        RECT -49.125 105.235 -48.795 105.565 ;
        RECT -49.125 103.875 -48.795 104.205 ;
        RECT -49.125 102.515 -48.795 102.845 ;
        RECT -49.125 101.155 -48.795 101.485 ;
        RECT -49.125 99.795 -48.795 100.125 ;
        RECT -49.125 98.435 -48.795 98.765 ;
        RECT -49.125 97.075 -48.795 97.405 ;
        RECT -49.125 95.715 -48.795 96.045 ;
        RECT -49.125 94.355 -48.795 94.685 ;
        RECT -49.125 92.995 -48.795 93.325 ;
        RECT -49.125 91.635 -48.795 91.965 ;
        RECT -49.125 90.275 -48.795 90.605 ;
        RECT -49.125 88.915 -48.795 89.245 ;
        RECT -49.125 87.555 -48.795 87.885 ;
        RECT -49.125 86.195 -48.795 86.525 ;
        RECT -49.125 84.835 -48.795 85.165 ;
        RECT -49.125 83.475 -48.795 83.805 ;
        RECT -49.125 82.115 -48.795 82.445 ;
        RECT -49.125 80.755 -48.795 81.085 ;
        RECT -49.125 79.395 -48.795 79.725 ;
        RECT -49.125 78.035 -48.795 78.365 ;
        RECT -49.125 76.675 -48.795 77.005 ;
        RECT -49.125 75.315 -48.795 75.645 ;
        RECT -49.125 73.955 -48.795 74.285 ;
        RECT -49.12 73.28 -48.8 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.125 -184.445 -48.795 -184.115 ;
        RECT -49.125 -185.805 -48.795 -185.475 ;
        RECT -49.125 -187.165 -48.795 -186.835 ;
        RECT -49.125 -188.525 -48.795 -188.195 ;
        RECT -49.125 -189.885 -48.795 -189.555 ;
        RECT -49.125 -191.245 -48.795 -190.915 ;
        RECT -49.125 -192.605 -48.795 -192.275 ;
        RECT -49.125 -193.965 -48.795 -193.635 ;
        RECT -49.125 -195.325 -48.795 -194.995 ;
        RECT -49.125 -196.685 -48.795 -196.355 ;
        RECT -49.125 -198.045 -48.795 -197.715 ;
        RECT -49.125 -199.405 -48.795 -199.075 ;
        RECT -49.125 -200.765 -48.795 -200.435 ;
        RECT -49.125 -202.125 -48.795 -201.795 ;
        RECT -49.125 -203.485 -48.795 -203.155 ;
        RECT -49.125 -204.845 -48.795 -204.515 ;
        RECT -49.125 -206.555 -48.795 -206.225 ;
        RECT -49.125 -207.565 -48.795 -207.235 ;
        RECT -49.125 -208.925 -48.795 -208.595 ;
        RECT -49.125 -210.285 -48.795 -209.955 ;
        RECT -49.125 -211.645 -48.795 -211.315 ;
        RECT -49.125 -214.365 -48.795 -214.035 ;
        RECT -49.125 -215.725 -48.795 -215.395 ;
        RECT -49.125 -217.085 -48.795 -216.755 ;
        RECT -49.125 -218.445 -48.795 -218.115 ;
        RECT -49.125 -224.09 -48.795 -222.96 ;
        RECT -49.12 -224.205 -48.8 49.12 ;
        RECT -49.125 48.115 -48.795 48.445 ;
        RECT -49.125 46.755 -48.795 47.085 ;
        RECT -49.125 45.395 -48.795 45.725 ;
        RECT -49.125 44.035 -48.795 44.365 ;
        RECT -49.125 39.955 -48.795 40.285 ;
        RECT -49.125 38.595 -48.795 38.925 ;
        RECT -49.125 35.875 -48.795 36.205 ;
        RECT -49.125 34.515 -48.795 34.845 ;
        RECT -49.125 33.155 -48.795 33.485 ;
        RECT -49.125 31.795 -48.795 32.125 ;
        RECT -49.125 30.435 -48.795 30.765 ;
        RECT -49.125 29.075 -48.795 29.405 ;
        RECT -49.125 27.715 -48.795 28.045 ;
        RECT -49.125 26.355 -48.795 26.685 ;
        RECT -49.125 24.995 -48.795 25.325 ;
        RECT -49.125 23.635 -48.795 23.965 ;
        RECT -49.125 22.275 -48.795 22.605 ;
        RECT -49.125 20.915 -48.795 21.245 ;
        RECT -49.125 19.555 -48.795 19.885 ;
        RECT -49.125 18.195 -48.795 18.525 ;
        RECT -49.125 16.835 -48.795 17.165 ;
        RECT -49.125 15.475 -48.795 15.805 ;
        RECT -49.125 14.115 -48.795 14.445 ;
        RECT -49.125 12.755 -48.795 13.085 ;
        RECT -49.125 11.395 -48.795 11.725 ;
        RECT -49.125 10.035 -48.795 10.365 ;
        RECT -49.125 8.675 -48.795 9.005 ;
        RECT -49.125 7.315 -48.795 7.645 ;
        RECT -49.125 5.955 -48.795 6.285 ;
        RECT -49.125 4.595 -48.795 4.925 ;
        RECT -49.125 3.235 -48.795 3.565 ;
        RECT -49.125 1.875 -48.795 2.205 ;
        RECT -49.125 0.515 -48.795 0.845 ;
        RECT -49.125 -0.845 -48.795 -0.515 ;
        RECT -49.125 -2.205 -48.795 -1.875 ;
        RECT -49.125 -3.565 -48.795 -3.235 ;
        RECT -49.125 -4.925 -48.795 -4.595 ;
        RECT -49.125 -6.285 -48.795 -5.955 ;
        RECT -49.125 -7.645 -48.795 -7.315 ;
        RECT -49.125 -9.005 -48.795 -8.675 ;
        RECT -49.125 -11.725 -48.795 -11.395 ;
        RECT -49.125 -13.085 -48.795 -12.755 ;
        RECT -49.125 -14.445 -48.795 -14.115 ;
        RECT -49.125 -15.805 -48.795 -15.475 ;
        RECT -49.125 -17.165 -48.795 -16.835 ;
        RECT -49.125 -18.525 -48.795 -18.195 ;
        RECT -49.125 -19.885 -48.795 -19.555 ;
        RECT -49.125 -21.245 -48.795 -20.915 ;
        RECT -49.125 -22.605 -48.795 -22.275 ;
        RECT -49.125 -23.965 -48.795 -23.635 ;
        RECT -49.125 -25.325 -48.795 -24.995 ;
        RECT -49.125 -26.685 -48.795 -26.355 ;
        RECT -49.125 -28.045 -48.795 -27.715 ;
        RECT -49.125 -29.405 -48.795 -29.075 ;
        RECT -49.125 -30.765 -48.795 -30.435 ;
        RECT -49.125 -32.125 -48.795 -31.795 ;
        RECT -49.125 -33.485 -48.795 -33.155 ;
        RECT -49.125 -34.845 -48.795 -34.515 ;
        RECT -49.125 -37.565 -48.795 -37.235 ;
        RECT -49.125 -38.925 -48.795 -38.595 ;
        RECT -49.125 -40.285 -48.795 -39.955 ;
        RECT -49.125 -41.645 -48.795 -41.315 ;
        RECT -49.125 -43.005 -48.795 -42.675 ;
        RECT -49.125 -44.365 -48.795 -44.035 ;
        RECT -49.125 -45.725 -48.795 -45.395 ;
        RECT -49.125 -47.085 -48.795 -46.755 ;
        RECT -49.125 -48.445 -48.795 -48.115 ;
        RECT -49.125 -49.805 -48.795 -49.475 ;
        RECT -49.125 -51.165 -48.795 -50.835 ;
        RECT -49.125 -52.525 -48.795 -52.195 ;
        RECT -49.125 -53.885 -48.795 -53.555 ;
        RECT -49.125 -55.245 -48.795 -54.915 ;
        RECT -49.125 -56.605 -48.795 -56.275 ;
        RECT -49.125 -57.965 -48.795 -57.635 ;
        RECT -49.125 -59.325 -48.795 -58.995 ;
        RECT -49.125 -60.685 -48.795 -60.355 ;
        RECT -49.125 -62.045 -48.795 -61.715 ;
        RECT -49.125 -63.405 -48.795 -63.075 ;
        RECT -49.125 -64.765 -48.795 -64.435 ;
        RECT -49.125 -66.125 -48.795 -65.795 ;
        RECT -49.125 -67.485 -48.795 -67.155 ;
        RECT -49.125 -68.845 -48.795 -68.515 ;
        RECT -49.125 -70.205 -48.795 -69.875 ;
        RECT -49.125 -71.565 -48.795 -71.235 ;
        RECT -49.125 -72.925 -48.795 -72.595 ;
        RECT -49.125 -74.285 -48.795 -73.955 ;
        RECT -49.125 -75.645 -48.795 -75.315 ;
        RECT -49.125 -77.005 -48.795 -76.675 ;
        RECT -49.125 -78.365 -48.795 -78.035 ;
        RECT -49.125 -79.725 -48.795 -79.395 ;
        RECT -49.125 -81.085 -48.795 -80.755 ;
        RECT -49.125 -82.445 -48.795 -82.115 ;
        RECT -49.125 -83.805 -48.795 -83.475 ;
        RECT -49.125 -85.165 -48.795 -84.835 ;
        RECT -49.125 -86.525 -48.795 -86.195 ;
        RECT -49.125 -87.885 -48.795 -87.555 ;
        RECT -49.125 -89.245 -48.795 -88.915 ;
        RECT -49.125 -90.605 -48.795 -90.275 ;
        RECT -49.125 -91.965 -48.795 -91.635 ;
        RECT -49.125 -93.325 -48.795 -92.995 ;
        RECT -49.125 -94.685 -48.795 -94.355 ;
        RECT -49.125 -96.045 -48.795 -95.715 ;
        RECT -49.125 -97.405 -48.795 -97.075 ;
        RECT -49.125 -98.765 -48.795 -98.435 ;
        RECT -49.125 -100.125 -48.795 -99.795 ;
        RECT -49.125 -101.485 -48.795 -101.155 ;
        RECT -49.125 -102.845 -48.795 -102.515 ;
        RECT -49.125 -104.205 -48.795 -103.875 ;
        RECT -49.125 -105.565 -48.795 -105.235 ;
        RECT -49.125 -106.925 -48.795 -106.595 ;
        RECT -49.125 -108.285 -48.795 -107.955 ;
        RECT -49.125 -109.645 -48.795 -109.315 ;
        RECT -49.125 -111.005 -48.795 -110.675 ;
        RECT -49.125 -111.87 -48.795 -111.54 ;
        RECT -49.125 -113.725 -48.795 -113.395 ;
        RECT -49.125 -115.085 -48.795 -114.755 ;
        RECT -49.125 -116.445 -48.795 -116.115 ;
        RECT -49.125 -117.805 -48.795 -117.475 ;
        RECT -49.125 -120.525 -48.795 -120.195 ;
        RECT -49.125 -121.885 -48.795 -121.555 ;
        RECT -49.125 -123.245 -48.795 -122.915 ;
        RECT -49.125 -124.71 -48.795 -124.38 ;
        RECT -49.125 -125.965 -48.795 -125.635 ;
        RECT -49.125 -127.325 -48.795 -126.995 ;
        RECT -49.125 -130.045 -48.795 -129.715 ;
        RECT -49.125 -135.485 -48.795 -135.155 ;
        RECT -49.125 -136.845 -48.795 -136.515 ;
        RECT -49.125 -138.205 -48.795 -137.875 ;
        RECT -49.125 -139.565 -48.795 -139.235 ;
        RECT -49.125 -142.285 -48.795 -141.955 ;
        RECT -49.125 -143.645 -48.795 -143.315 ;
        RECT -49.125 -145.005 -48.795 -144.675 ;
        RECT -49.125 -146.365 -48.795 -146.035 ;
        RECT -49.125 -147.725 -48.795 -147.395 ;
        RECT -49.125 -149.085 -48.795 -148.755 ;
        RECT -49.125 -150.445 -48.795 -150.115 ;
        RECT -49.125 -151.805 -48.795 -151.475 ;
        RECT -49.125 -153.165 -48.795 -152.835 ;
        RECT -49.125 -154.525 -48.795 -154.195 ;
        RECT -49.125 -155.885 -48.795 -155.555 ;
        RECT -49.125 -157.245 -48.795 -156.915 ;
        RECT -49.125 -158.605 -48.795 -158.275 ;
        RECT -49.125 -159.965 -48.795 -159.635 ;
        RECT -49.125 -161.325 -48.795 -160.995 ;
        RECT -49.125 -162.685 -48.795 -162.355 ;
        RECT -49.125 -164.045 -48.795 -163.715 ;
        RECT -49.125 -165.405 -48.795 -165.075 ;
        RECT -49.125 -166.765 -48.795 -166.435 ;
        RECT -49.125 -168.125 -48.795 -167.795 ;
        RECT -49.125 -169.485 -48.795 -169.155 ;
        RECT -49.125 -170.845 -48.795 -170.515 ;
        RECT -49.125 -172.205 -48.795 -171.875 ;
        RECT -49.125 -173.565 -48.795 -173.235 ;
        RECT -49.125 -174.925 -48.795 -174.595 ;
        RECT -49.125 -176.285 -48.795 -175.955 ;
        RECT -49.125 -177.645 -48.795 -177.315 ;
        RECT -49.125 -179.005 -48.795 -178.675 ;
        RECT -49.125 -180.365 -48.795 -180.035 ;
        RECT -49.125 -181.725 -48.795 -181.395 ;
        RECT -49.125 -183.085 -48.795 -182.755 ;
    END
    PORT
      LAYER met3 ;
        RECT -60.005 132.52 -59.675 133.65 ;
        RECT -60.005 128.355 -59.675 128.685 ;
        RECT -60.005 126.995 -59.675 127.325 ;
        RECT -60.005 125.635 -59.675 125.965 ;
        RECT -60.005 124.275 -59.675 124.605 ;
        RECT -60.005 122.915 -59.675 123.245 ;
        RECT -60.005 121.555 -59.675 121.885 ;
        RECT -60.005 120.195 -59.675 120.525 ;
        RECT -60.005 118.835 -59.675 119.165 ;
        RECT -60.005 117.475 -59.675 117.805 ;
        RECT -60.005 116.115 -59.675 116.445 ;
        RECT -60.005 114.755 -59.675 115.085 ;
        RECT -60.005 113.395 -59.675 113.725 ;
        RECT -60.005 112.035 -59.675 112.365 ;
        RECT -60.005 110.675 -59.675 111.005 ;
        RECT -60.005 109.315 -59.675 109.645 ;
        RECT -60.005 107.955 -59.675 108.285 ;
        RECT -60.005 106.595 -59.675 106.925 ;
        RECT -60.005 105.235 -59.675 105.565 ;
        RECT -60.005 103.875 -59.675 104.205 ;
        RECT -60.005 102.515 -59.675 102.845 ;
        RECT -60.005 101.155 -59.675 101.485 ;
        RECT -60.005 99.795 -59.675 100.125 ;
        RECT -60.005 98.435 -59.675 98.765 ;
        RECT -60.005 97.075 -59.675 97.405 ;
        RECT -60.005 95.715 -59.675 96.045 ;
        RECT -60.005 94.355 -59.675 94.685 ;
        RECT -60.005 92.995 -59.675 93.325 ;
        RECT -60.005 91.635 -59.675 91.965 ;
        RECT -60.005 90.275 -59.675 90.605 ;
        RECT -60.005 88.915 -59.675 89.245 ;
        RECT -60.005 87.555 -59.675 87.885 ;
        RECT -60.005 86.195 -59.675 86.525 ;
        RECT -60.005 84.835 -59.675 85.165 ;
        RECT -60.005 83.475 -59.675 83.805 ;
        RECT -60.005 82.115 -59.675 82.445 ;
        RECT -60.005 80.755 -59.675 81.085 ;
        RECT -60.005 79.395 -59.675 79.725 ;
        RECT -60.005 78.035 -59.675 78.365 ;
        RECT -60.005 76.675 -59.675 77.005 ;
        RECT -60.005 75.315 -59.675 75.645 ;
        RECT -60.005 73.955 -59.675 74.285 ;
        RECT -60.005 72.595 -59.675 72.925 ;
        RECT -60.005 71.235 -59.675 71.565 ;
        RECT -60.005 69.875 -59.675 70.205 ;
        RECT -60.005 68.515 -59.675 68.845 ;
        RECT -60.005 67.155 -59.675 67.485 ;
        RECT -60.005 65.795 -59.675 66.125 ;
        RECT -60.005 64.435 -59.675 64.765 ;
        RECT -60.005 63.075 -59.675 63.405 ;
        RECT -60.005 61.715 -59.675 62.045 ;
        RECT -60.005 60.355 -59.675 60.685 ;
        RECT -60.005 58.995 -59.675 59.325 ;
        RECT -60.005 57.635 -59.675 57.965 ;
        RECT -60.005 56.275 -59.675 56.605 ;
        RECT -60.005 54.915 -59.675 55.245 ;
        RECT -60.005 53.555 -59.675 53.885 ;
        RECT -60.005 52.195 -59.675 52.525 ;
        RECT -60.005 50.835 -59.675 51.165 ;
        RECT -60.005 49.475 -59.675 49.805 ;
        RECT -60.005 48.115 -59.675 48.445 ;
        RECT -60.005 46.755 -59.675 47.085 ;
        RECT -60.005 45.395 -59.675 45.725 ;
        RECT -60.005 44.035 -59.675 44.365 ;
        RECT -60.005 42.675 -59.675 43.005 ;
        RECT -60.005 41.315 -59.675 41.645 ;
        RECT -60.005 39.955 -59.675 40.285 ;
        RECT -60.005 38.595 -59.675 38.925 ;
        RECT -60.005 37.235 -59.675 37.565 ;
        RECT -60.005 35.875 -59.675 36.205 ;
        RECT -60.005 34.515 -59.675 34.845 ;
        RECT -60.005 33.155 -59.675 33.485 ;
        RECT -60.005 31.795 -59.675 32.125 ;
        RECT -60.005 30.435 -59.675 30.765 ;
        RECT -60.005 29.075 -59.675 29.405 ;
        RECT -60.005 27.715 -59.675 28.045 ;
        RECT -60.005 26.355 -59.675 26.685 ;
        RECT -60.005 24.995 -59.675 25.325 ;
        RECT -60.005 23.635 -59.675 23.965 ;
        RECT -60.005 22.275 -59.675 22.605 ;
        RECT -60.005 20.915 -59.675 21.245 ;
        RECT -60.005 19.555 -59.675 19.885 ;
        RECT -60.005 18.195 -59.675 18.525 ;
        RECT -60.005 16.835 -59.675 17.165 ;
        RECT -60.005 15.475 -59.675 15.805 ;
        RECT -60.005 14.115 -59.675 14.445 ;
        RECT -60.005 12.755 -59.675 13.085 ;
        RECT -60.005 11.395 -59.675 11.725 ;
        RECT -60.005 10.035 -59.675 10.365 ;
        RECT -60.005 8.675 -59.675 9.005 ;
        RECT -60.005 7.315 -59.675 7.645 ;
        RECT -60.005 5.955 -59.675 6.285 ;
        RECT -60.005 4.595 -59.675 4.925 ;
        RECT -60.005 3.235 -59.675 3.565 ;
        RECT -60.005 1.875 -59.675 2.205 ;
        RECT -60.005 0.515 -59.675 0.845 ;
        RECT -60.005 -0.845 -59.675 -0.515 ;
        RECT -60.005 -2.205 -59.675 -1.875 ;
        RECT -60.005 -3.565 -59.675 -3.235 ;
        RECT -60.005 -4.925 -59.675 -4.595 ;
        RECT -60.005 -6.285 -59.675 -5.955 ;
        RECT -60.005 -7.645 -59.675 -7.315 ;
        RECT -60.005 -9.005 -59.675 -8.675 ;
        RECT -60.005 -10.365 -59.675 -10.035 ;
        RECT -60.005 -11.725 -59.675 -11.395 ;
        RECT -60.005 -13.085 -59.675 -12.755 ;
        RECT -60.005 -14.445 -59.675 -14.115 ;
        RECT -60.005 -15.805 -59.675 -15.475 ;
        RECT -60.005 -17.165 -59.675 -16.835 ;
        RECT -60.005 -18.525 -59.675 -18.195 ;
        RECT -60.005 -19.885 -59.675 -19.555 ;
        RECT -60.005 -21.245 -59.675 -20.915 ;
        RECT -60.005 -22.605 -59.675 -22.275 ;
        RECT -60.005 -23.965 -59.675 -23.635 ;
        RECT -60.005 -25.325 -59.675 -24.995 ;
        RECT -60.005 -26.685 -59.675 -26.355 ;
        RECT -60.005 -28.045 -59.675 -27.715 ;
        RECT -60.005 -29.405 -59.675 -29.075 ;
        RECT -60.005 -30.765 -59.675 -30.435 ;
        RECT -60.005 -32.125 -59.675 -31.795 ;
        RECT -60.005 -33.485 -59.675 -33.155 ;
        RECT -60.005 -34.845 -59.675 -34.515 ;
        RECT -60.005 -36.205 -59.675 -35.875 ;
        RECT -60.005 -37.565 -59.675 -37.235 ;
        RECT -60.005 -38.925 -59.675 -38.595 ;
        RECT -60.005 -40.285 -59.675 -39.955 ;
        RECT -60.005 -41.645 -59.675 -41.315 ;
        RECT -60.005 -43.005 -59.675 -42.675 ;
        RECT -60.005 -44.365 -59.675 -44.035 ;
        RECT -60.005 -45.725 -59.675 -45.395 ;
        RECT -60.005 -47.085 -59.675 -46.755 ;
        RECT -60.005 -48.445 -59.675 -48.115 ;
        RECT -60.005 -49.805 -59.675 -49.475 ;
        RECT -60.005 -51.165 -59.675 -50.835 ;
        RECT -60.005 -52.525 -59.675 -52.195 ;
        RECT -60.005 -53.885 -59.675 -53.555 ;
        RECT -60.005 -55.245 -59.675 -54.915 ;
        RECT -60.005 -56.605 -59.675 -56.275 ;
        RECT -60.005 -57.965 -59.675 -57.635 ;
        RECT -60.005 -59.325 -59.675 -58.995 ;
        RECT -60.005 -60.685 -59.675 -60.355 ;
        RECT -60.005 -62.045 -59.675 -61.715 ;
        RECT -60.005 -63.405 -59.675 -63.075 ;
        RECT -60.005 -64.765 -59.675 -64.435 ;
        RECT -60.005 -66.125 -59.675 -65.795 ;
        RECT -60.005 -67.485 -59.675 -67.155 ;
        RECT -60.005 -68.845 -59.675 -68.515 ;
        RECT -60.005 -70.205 -59.675 -69.875 ;
        RECT -60.005 -71.565 -59.675 -71.235 ;
        RECT -60.005 -72.925 -59.675 -72.595 ;
        RECT -60.005 -74.285 -59.675 -73.955 ;
        RECT -60.005 -75.645 -59.675 -75.315 ;
        RECT -60.005 -77.005 -59.675 -76.675 ;
        RECT -60.005 -78.365 -59.675 -78.035 ;
        RECT -60.005 -79.725 -59.675 -79.395 ;
        RECT -60.005 -81.085 -59.675 -80.755 ;
        RECT -60.005 -82.445 -59.675 -82.115 ;
        RECT -60.005 -83.805 -59.675 -83.475 ;
        RECT -60.005 -85.165 -59.675 -84.835 ;
        RECT -60.005 -86.525 -59.675 -86.195 ;
        RECT -60.005 -87.885 -59.675 -87.555 ;
        RECT -60.005 -89.245 -59.675 -88.915 ;
        RECT -60.005 -90.605 -59.675 -90.275 ;
        RECT -60.005 -91.965 -59.675 -91.635 ;
        RECT -60.005 -93.325 -59.675 -92.995 ;
        RECT -60.005 -94.685 -59.675 -94.355 ;
        RECT -60.005 -96.045 -59.675 -95.715 ;
        RECT -60.005 -97.405 -59.675 -97.075 ;
        RECT -60.005 -98.765 -59.675 -98.435 ;
        RECT -60.005 -100.125 -59.675 -99.795 ;
        RECT -60.005 -101.485 -59.675 -101.155 ;
        RECT -60.005 -102.845 -59.675 -102.515 ;
        RECT -60.005 -104.205 -59.675 -103.875 ;
        RECT -60.005 -105.565 -59.675 -105.235 ;
        RECT -60.005 -106.925 -59.675 -106.595 ;
        RECT -60.005 -108.285 -59.675 -107.955 ;
        RECT -60.005 -109.645 -59.675 -109.315 ;
        RECT -60.005 -111.005 -59.675 -110.675 ;
        RECT -60.005 -112.365 -59.675 -112.035 ;
        RECT -60.005 -113.725 -59.675 -113.395 ;
        RECT -60.005 -115.085 -59.675 -114.755 ;
        RECT -60.005 -116.445 -59.675 -116.115 ;
        RECT -60.005 -117.805 -59.675 -117.475 ;
        RECT -60.005 -119.165 -59.675 -118.835 ;
        RECT -60.005 -120.525 -59.675 -120.195 ;
        RECT -60.005 -121.885 -59.675 -121.555 ;
        RECT -60.005 -123.245 -59.675 -122.915 ;
        RECT -60.005 -124.605 -59.675 -124.275 ;
        RECT -60.005 -125.965 -59.675 -125.635 ;
        RECT -60.005 -127.325 -59.675 -126.995 ;
        RECT -60.005 -128.685 -59.675 -128.355 ;
        RECT -60.005 -130.045 -59.675 -129.715 ;
        RECT -60.005 -131.405 -59.675 -131.075 ;
        RECT -60 -132.08 -59.68 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -60.005 -214.365 -59.675 -214.035 ;
        RECT -60.005 -215.725 -59.675 -215.395 ;
        RECT -60.005 -217.085 -59.675 -216.755 ;
        RECT -60.005 -218.445 -59.675 -218.115 ;
        RECT -60.005 -224.09 -59.675 -222.96 ;
        RECT -60 -224.205 -59.68 -210.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -58.645 132.52 -58.315 133.65 ;
        RECT -58.645 128.355 -58.315 128.685 ;
        RECT -58.645 126.995 -58.315 127.325 ;
        RECT -58.645 125.635 -58.315 125.965 ;
        RECT -58.645 124.275 -58.315 124.605 ;
        RECT -58.645 122.915 -58.315 123.245 ;
        RECT -58.645 121.555 -58.315 121.885 ;
        RECT -58.645 120.195 -58.315 120.525 ;
        RECT -58.645 118.835 -58.315 119.165 ;
        RECT -58.645 117.475 -58.315 117.805 ;
        RECT -58.645 116.115 -58.315 116.445 ;
        RECT -58.645 114.755 -58.315 115.085 ;
        RECT -58.645 113.395 -58.315 113.725 ;
        RECT -58.645 112.035 -58.315 112.365 ;
        RECT -58.645 110.675 -58.315 111.005 ;
        RECT -58.645 109.315 -58.315 109.645 ;
        RECT -58.645 107.955 -58.315 108.285 ;
        RECT -58.645 106.595 -58.315 106.925 ;
        RECT -58.645 105.235 -58.315 105.565 ;
        RECT -58.645 103.875 -58.315 104.205 ;
        RECT -58.645 102.515 -58.315 102.845 ;
        RECT -58.645 101.155 -58.315 101.485 ;
        RECT -58.645 99.795 -58.315 100.125 ;
        RECT -58.645 98.435 -58.315 98.765 ;
        RECT -58.645 97.075 -58.315 97.405 ;
        RECT -58.645 95.715 -58.315 96.045 ;
        RECT -58.645 94.355 -58.315 94.685 ;
        RECT -58.645 92.995 -58.315 93.325 ;
        RECT -58.645 91.635 -58.315 91.965 ;
        RECT -58.645 90.275 -58.315 90.605 ;
        RECT -58.645 88.915 -58.315 89.245 ;
        RECT -58.645 87.555 -58.315 87.885 ;
        RECT -58.645 86.195 -58.315 86.525 ;
        RECT -58.645 84.835 -58.315 85.165 ;
        RECT -58.645 83.475 -58.315 83.805 ;
        RECT -58.645 82.115 -58.315 82.445 ;
        RECT -58.645 80.755 -58.315 81.085 ;
        RECT -58.645 79.395 -58.315 79.725 ;
        RECT -58.645 78.035 -58.315 78.365 ;
        RECT -58.645 76.675 -58.315 77.005 ;
        RECT -58.645 75.315 -58.315 75.645 ;
        RECT -58.645 73.955 -58.315 74.285 ;
        RECT -58.645 72.595 -58.315 72.925 ;
        RECT -58.645 71.235 -58.315 71.565 ;
        RECT -58.645 69.875 -58.315 70.205 ;
        RECT -58.645 68.515 -58.315 68.845 ;
        RECT -58.645 67.155 -58.315 67.485 ;
        RECT -58.645 65.795 -58.315 66.125 ;
        RECT -58.645 64.435 -58.315 64.765 ;
        RECT -58.645 63.075 -58.315 63.405 ;
        RECT -58.645 61.715 -58.315 62.045 ;
        RECT -58.645 60.355 -58.315 60.685 ;
        RECT -58.645 58.995 -58.315 59.325 ;
        RECT -58.645 57.635 -58.315 57.965 ;
        RECT -58.645 56.275 -58.315 56.605 ;
        RECT -58.645 54.915 -58.315 55.245 ;
        RECT -58.645 53.555 -58.315 53.885 ;
        RECT -58.645 52.195 -58.315 52.525 ;
        RECT -58.645 50.835 -58.315 51.165 ;
        RECT -58.645 49.475 -58.315 49.805 ;
        RECT -58.645 48.115 -58.315 48.445 ;
        RECT -58.645 46.755 -58.315 47.085 ;
        RECT -58.645 45.395 -58.315 45.725 ;
        RECT -58.645 44.035 -58.315 44.365 ;
        RECT -58.645 42.675 -58.315 43.005 ;
        RECT -58.645 41.315 -58.315 41.645 ;
        RECT -58.645 39.955 -58.315 40.285 ;
        RECT -58.645 38.595 -58.315 38.925 ;
        RECT -58.645 37.235 -58.315 37.565 ;
        RECT -58.645 35.875 -58.315 36.205 ;
        RECT -58.645 34.515 -58.315 34.845 ;
        RECT -58.645 33.155 -58.315 33.485 ;
        RECT -58.645 31.795 -58.315 32.125 ;
        RECT -58.645 30.435 -58.315 30.765 ;
        RECT -58.645 29.075 -58.315 29.405 ;
        RECT -58.645 27.715 -58.315 28.045 ;
        RECT -58.645 26.355 -58.315 26.685 ;
        RECT -58.645 24.995 -58.315 25.325 ;
        RECT -58.645 23.635 -58.315 23.965 ;
        RECT -58.645 22.275 -58.315 22.605 ;
        RECT -58.645 20.915 -58.315 21.245 ;
        RECT -58.645 19.555 -58.315 19.885 ;
        RECT -58.645 18.195 -58.315 18.525 ;
        RECT -58.645 16.835 -58.315 17.165 ;
        RECT -58.645 15.475 -58.315 15.805 ;
        RECT -58.645 14.115 -58.315 14.445 ;
        RECT -58.645 12.755 -58.315 13.085 ;
        RECT -58.645 11.395 -58.315 11.725 ;
        RECT -58.645 10.035 -58.315 10.365 ;
        RECT -58.645 8.675 -58.315 9.005 ;
        RECT -58.645 7.315 -58.315 7.645 ;
        RECT -58.645 5.955 -58.315 6.285 ;
        RECT -58.645 4.595 -58.315 4.925 ;
        RECT -58.645 3.235 -58.315 3.565 ;
        RECT -58.645 1.875 -58.315 2.205 ;
        RECT -58.645 0.515 -58.315 0.845 ;
        RECT -58.645 -0.845 -58.315 -0.515 ;
        RECT -58.645 -2.205 -58.315 -1.875 ;
        RECT -58.645 -3.565 -58.315 -3.235 ;
        RECT -58.645 -4.925 -58.315 -4.595 ;
        RECT -58.645 -6.285 -58.315 -5.955 ;
        RECT -58.645 -7.645 -58.315 -7.315 ;
        RECT -58.645 -9.005 -58.315 -8.675 ;
        RECT -58.645 -10.365 -58.315 -10.035 ;
        RECT -58.645 -11.725 -58.315 -11.395 ;
        RECT -58.645 -13.085 -58.315 -12.755 ;
        RECT -58.645 -14.445 -58.315 -14.115 ;
        RECT -58.645 -15.805 -58.315 -15.475 ;
        RECT -58.645 -17.165 -58.315 -16.835 ;
        RECT -58.645 -18.525 -58.315 -18.195 ;
        RECT -58.645 -19.885 -58.315 -19.555 ;
        RECT -58.645 -21.245 -58.315 -20.915 ;
        RECT -58.645 -22.605 -58.315 -22.275 ;
        RECT -58.645 -23.965 -58.315 -23.635 ;
        RECT -58.645 -25.325 -58.315 -24.995 ;
        RECT -58.645 -26.685 -58.315 -26.355 ;
        RECT -58.645 -28.045 -58.315 -27.715 ;
        RECT -58.645 -29.405 -58.315 -29.075 ;
        RECT -58.645 -30.765 -58.315 -30.435 ;
        RECT -58.645 -32.125 -58.315 -31.795 ;
        RECT -58.645 -33.485 -58.315 -33.155 ;
        RECT -58.645 -34.845 -58.315 -34.515 ;
        RECT -58.645 -36.205 -58.315 -35.875 ;
        RECT -58.645 -37.565 -58.315 -37.235 ;
        RECT -58.645 -38.925 -58.315 -38.595 ;
        RECT -58.645 -40.285 -58.315 -39.955 ;
        RECT -58.645 -41.645 -58.315 -41.315 ;
        RECT -58.645 -43.005 -58.315 -42.675 ;
        RECT -58.645 -44.365 -58.315 -44.035 ;
        RECT -58.645 -45.725 -58.315 -45.395 ;
        RECT -58.645 -47.085 -58.315 -46.755 ;
        RECT -58.645 -48.445 -58.315 -48.115 ;
        RECT -58.645 -49.805 -58.315 -49.475 ;
        RECT -58.645 -51.165 -58.315 -50.835 ;
        RECT -58.645 -52.525 -58.315 -52.195 ;
        RECT -58.645 -53.885 -58.315 -53.555 ;
        RECT -58.645 -55.245 -58.315 -54.915 ;
        RECT -58.645 -56.605 -58.315 -56.275 ;
        RECT -58.645 -57.965 -58.315 -57.635 ;
        RECT -58.645 -59.325 -58.315 -58.995 ;
        RECT -58.645 -60.685 -58.315 -60.355 ;
        RECT -58.645 -62.045 -58.315 -61.715 ;
        RECT -58.645 -63.405 -58.315 -63.075 ;
        RECT -58.645 -64.765 -58.315 -64.435 ;
        RECT -58.645 -66.125 -58.315 -65.795 ;
        RECT -58.645 -67.485 -58.315 -67.155 ;
        RECT -58.645 -68.845 -58.315 -68.515 ;
        RECT -58.645 -70.205 -58.315 -69.875 ;
        RECT -58.645 -71.565 -58.315 -71.235 ;
        RECT -58.645 -72.925 -58.315 -72.595 ;
        RECT -58.645 -74.285 -58.315 -73.955 ;
        RECT -58.645 -75.645 -58.315 -75.315 ;
        RECT -58.645 -77.005 -58.315 -76.675 ;
        RECT -58.645 -78.365 -58.315 -78.035 ;
        RECT -58.645 -79.725 -58.315 -79.395 ;
        RECT -58.645 -81.085 -58.315 -80.755 ;
        RECT -58.645 -82.445 -58.315 -82.115 ;
        RECT -58.645 -83.805 -58.315 -83.475 ;
        RECT -58.645 -85.165 -58.315 -84.835 ;
        RECT -58.645 -86.525 -58.315 -86.195 ;
        RECT -58.645 -87.885 -58.315 -87.555 ;
        RECT -58.645 -89.245 -58.315 -88.915 ;
        RECT -58.645 -90.605 -58.315 -90.275 ;
        RECT -58.645 -91.965 -58.315 -91.635 ;
        RECT -58.645 -93.325 -58.315 -92.995 ;
        RECT -58.645 -94.685 -58.315 -94.355 ;
        RECT -58.645 -96.045 -58.315 -95.715 ;
        RECT -58.645 -97.405 -58.315 -97.075 ;
        RECT -58.645 -98.765 -58.315 -98.435 ;
        RECT -58.645 -100.125 -58.315 -99.795 ;
        RECT -58.645 -101.485 -58.315 -101.155 ;
        RECT -58.645 -102.845 -58.315 -102.515 ;
        RECT -58.645 -104.205 -58.315 -103.875 ;
        RECT -58.645 -105.565 -58.315 -105.235 ;
        RECT -58.645 -106.925 -58.315 -106.595 ;
        RECT -58.645 -108.285 -58.315 -107.955 ;
        RECT -58.645 -109.645 -58.315 -109.315 ;
        RECT -58.645 -111.005 -58.315 -110.675 ;
        RECT -58.645 -112.365 -58.315 -112.035 ;
        RECT -58.645 -113.725 -58.315 -113.395 ;
        RECT -58.645 -115.085 -58.315 -114.755 ;
        RECT -58.645 -116.445 -58.315 -116.115 ;
        RECT -58.645 -117.805 -58.315 -117.475 ;
        RECT -58.645 -119.165 -58.315 -118.835 ;
        RECT -58.645 -120.525 -58.315 -120.195 ;
        RECT -58.645 -121.885 -58.315 -121.555 ;
        RECT -58.645 -123.245 -58.315 -122.915 ;
        RECT -58.645 -124.605 -58.315 -124.275 ;
        RECT -58.645 -125.965 -58.315 -125.635 ;
        RECT -58.645 -127.325 -58.315 -126.995 ;
        RECT -58.645 -128.685 -58.315 -128.355 ;
        RECT -58.645 -130.045 -58.315 -129.715 ;
        RECT -58.645 -131.405 -58.315 -131.075 ;
        RECT -58.645 -134.125 -58.315 -133.795 ;
        RECT -58.645 -135.485 -58.315 -135.155 ;
        RECT -58.645 -136.845 -58.315 -136.515 ;
        RECT -58.645 -138.205 -58.315 -137.875 ;
        RECT -58.645 -139.565 -58.315 -139.235 ;
        RECT -58.645 -140.925 -58.315 -140.595 ;
        RECT -58.645 -142.285 -58.315 -141.955 ;
        RECT -58.645 -143.645 -58.315 -143.315 ;
        RECT -58.645 -145.005 -58.315 -144.675 ;
        RECT -58.645 -146.365 -58.315 -146.035 ;
        RECT -58.645 -147.725 -58.315 -147.395 ;
        RECT -58.645 -149.085 -58.315 -148.755 ;
        RECT -58.645 -150.445 -58.315 -150.115 ;
        RECT -58.645 -151.805 -58.315 -151.475 ;
        RECT -58.645 -153.165 -58.315 -152.835 ;
        RECT -58.645 -154.525 -58.315 -154.195 ;
        RECT -58.645 -155.885 -58.315 -155.555 ;
        RECT -58.645 -157.245 -58.315 -156.915 ;
        RECT -58.645 -158.605 -58.315 -158.275 ;
        RECT -58.645 -159.965 -58.315 -159.635 ;
        RECT -58.645 -161.325 -58.315 -160.995 ;
        RECT -58.645 -162.685 -58.315 -162.355 ;
        RECT -58.645 -164.045 -58.315 -163.715 ;
        RECT -58.645 -165.405 -58.315 -165.075 ;
        RECT -58.645 -166.765 -58.315 -166.435 ;
        RECT -58.645 -168.125 -58.315 -167.795 ;
        RECT -58.645 -169.485 -58.315 -169.155 ;
        RECT -58.645 -170.845 -58.315 -170.515 ;
        RECT -58.645 -172.205 -58.315 -171.875 ;
        RECT -58.645 -173.565 -58.315 -173.235 ;
        RECT -58.645 -174.925 -58.315 -174.595 ;
        RECT -58.645 -176.285 -58.315 -175.955 ;
        RECT -58.645 -177.645 -58.315 -177.315 ;
        RECT -58.645 -179.005 -58.315 -178.675 ;
        RECT -58.645 -180.365 -58.315 -180.035 ;
        RECT -58.645 -181.725 -58.315 -181.395 ;
        RECT -58.645 -183.085 -58.315 -182.755 ;
        RECT -58.645 -184.445 -58.315 -184.115 ;
        RECT -58.645 -185.805 -58.315 -185.475 ;
        RECT -58.645 -187.165 -58.315 -186.835 ;
        RECT -58.645 -188.525 -58.315 -188.195 ;
        RECT -58.645 -189.885 -58.315 -189.555 ;
        RECT -58.645 -191.245 -58.315 -190.915 ;
        RECT -58.645 -192.605 -58.315 -192.275 ;
        RECT -58.645 -193.965 -58.315 -193.635 ;
        RECT -58.645 -195.325 -58.315 -194.995 ;
        RECT -58.645 -196.685 -58.315 -196.355 ;
        RECT -58.645 -198.045 -58.315 -197.715 ;
        RECT -58.645 -199.405 -58.315 -199.075 ;
        RECT -58.645 -200.765 -58.315 -200.435 ;
        RECT -58.645 -202.125 -58.315 -201.795 ;
        RECT -58.645 -203.485 -58.315 -203.155 ;
        RECT -58.645 -204.845 -58.315 -204.515 ;
        RECT -58.645 -206.555 -58.315 -206.225 ;
        RECT -58.645 -207.565 -58.315 -207.235 ;
        RECT -58.645 -208.925 -58.315 -208.595 ;
        RECT -58.64 -209.6 -58.32 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -57.285 132.52 -56.955 133.65 ;
        RECT -57.285 128.355 -56.955 128.685 ;
        RECT -57.285 126.995 -56.955 127.325 ;
        RECT -57.285 125.635 -56.955 125.965 ;
        RECT -57.285 124.275 -56.955 124.605 ;
        RECT -57.285 122.915 -56.955 123.245 ;
        RECT -57.285 121.555 -56.955 121.885 ;
        RECT -57.285 120.195 -56.955 120.525 ;
        RECT -57.285 118.835 -56.955 119.165 ;
        RECT -57.285 117.475 -56.955 117.805 ;
        RECT -57.285 116.115 -56.955 116.445 ;
        RECT -57.285 114.755 -56.955 115.085 ;
        RECT -57.285 113.395 -56.955 113.725 ;
        RECT -57.285 112.035 -56.955 112.365 ;
        RECT -57.285 110.675 -56.955 111.005 ;
        RECT -57.285 109.315 -56.955 109.645 ;
        RECT -57.285 107.955 -56.955 108.285 ;
        RECT -57.285 106.595 -56.955 106.925 ;
        RECT -57.285 105.235 -56.955 105.565 ;
        RECT -57.285 103.875 -56.955 104.205 ;
        RECT -57.285 102.515 -56.955 102.845 ;
        RECT -57.285 101.155 -56.955 101.485 ;
        RECT -57.285 99.795 -56.955 100.125 ;
        RECT -57.285 98.435 -56.955 98.765 ;
        RECT -57.285 97.075 -56.955 97.405 ;
        RECT -57.285 95.715 -56.955 96.045 ;
        RECT -57.285 94.355 -56.955 94.685 ;
        RECT -57.285 92.995 -56.955 93.325 ;
        RECT -57.285 91.635 -56.955 91.965 ;
        RECT -57.285 90.275 -56.955 90.605 ;
        RECT -57.285 88.915 -56.955 89.245 ;
        RECT -57.285 87.555 -56.955 87.885 ;
        RECT -57.285 86.195 -56.955 86.525 ;
        RECT -57.285 84.835 -56.955 85.165 ;
        RECT -57.285 83.475 -56.955 83.805 ;
        RECT -57.285 82.115 -56.955 82.445 ;
        RECT -57.285 80.755 -56.955 81.085 ;
        RECT -57.285 79.395 -56.955 79.725 ;
        RECT -57.285 78.035 -56.955 78.365 ;
        RECT -57.285 76.675 -56.955 77.005 ;
        RECT -57.285 75.315 -56.955 75.645 ;
        RECT -57.285 73.955 -56.955 74.285 ;
        RECT -57.285 48.115 -56.955 48.445 ;
        RECT -57.285 46.755 -56.955 47.085 ;
        RECT -57.285 45.395 -56.955 45.725 ;
        RECT -57.285 44.035 -56.955 44.365 ;
        RECT -57.285 42.675 -56.955 43.005 ;
        RECT -57.285 41.315 -56.955 41.645 ;
        RECT -57.285 39.955 -56.955 40.285 ;
        RECT -57.285 38.595 -56.955 38.925 ;
        RECT -57.285 37.235 -56.955 37.565 ;
        RECT -57.285 35.875 -56.955 36.205 ;
        RECT -57.285 34.515 -56.955 34.845 ;
        RECT -57.285 33.155 -56.955 33.485 ;
        RECT -57.285 31.795 -56.955 32.125 ;
        RECT -57.285 30.435 -56.955 30.765 ;
        RECT -57.285 29.075 -56.955 29.405 ;
        RECT -57.285 27.715 -56.955 28.045 ;
        RECT -57.285 26.355 -56.955 26.685 ;
        RECT -57.285 24.995 -56.955 25.325 ;
        RECT -57.285 23.635 -56.955 23.965 ;
        RECT -57.285 22.275 -56.955 22.605 ;
        RECT -57.285 20.915 -56.955 21.245 ;
        RECT -57.285 19.555 -56.955 19.885 ;
        RECT -57.285 18.195 -56.955 18.525 ;
        RECT -57.285 16.835 -56.955 17.165 ;
        RECT -57.285 15.475 -56.955 15.805 ;
        RECT -57.285 14.115 -56.955 14.445 ;
        RECT -57.285 12.755 -56.955 13.085 ;
        RECT -57.285 11.395 -56.955 11.725 ;
        RECT -57.285 10.035 -56.955 10.365 ;
        RECT -57.285 8.675 -56.955 9.005 ;
        RECT -57.285 7.315 -56.955 7.645 ;
        RECT -57.285 5.955 -56.955 6.285 ;
        RECT -57.285 4.595 -56.955 4.925 ;
        RECT -57.285 3.235 -56.955 3.565 ;
        RECT -57.285 1.875 -56.955 2.205 ;
        RECT -57.285 0.515 -56.955 0.845 ;
        RECT -57.285 -0.845 -56.955 -0.515 ;
        RECT -57.285 -2.205 -56.955 -1.875 ;
        RECT -57.285 -3.565 -56.955 -3.235 ;
        RECT -57.285 -4.925 -56.955 -4.595 ;
        RECT -57.285 -6.285 -56.955 -5.955 ;
        RECT -57.285 -7.645 -56.955 -7.315 ;
        RECT -57.285 -9.005 -56.955 -8.675 ;
        RECT -57.285 -10.365 -56.955 -10.035 ;
        RECT -57.285 -11.725 -56.955 -11.395 ;
        RECT -57.285 -13.085 -56.955 -12.755 ;
        RECT -57.285 -14.445 -56.955 -14.115 ;
        RECT -57.285 -15.805 -56.955 -15.475 ;
        RECT -57.285 -17.165 -56.955 -16.835 ;
        RECT -57.285 -18.525 -56.955 -18.195 ;
        RECT -57.285 -19.885 -56.955 -19.555 ;
        RECT -57.285 -21.245 -56.955 -20.915 ;
        RECT -57.285 -22.605 -56.955 -22.275 ;
        RECT -57.285 -23.965 -56.955 -23.635 ;
        RECT -57.285 -25.325 -56.955 -24.995 ;
        RECT -57.285 -26.685 -56.955 -26.355 ;
        RECT -57.285 -28.045 -56.955 -27.715 ;
        RECT -57.285 -29.405 -56.955 -29.075 ;
        RECT -57.285 -30.765 -56.955 -30.435 ;
        RECT -57.285 -32.125 -56.955 -31.795 ;
        RECT -57.285 -33.485 -56.955 -33.155 ;
        RECT -57.285 -34.845 -56.955 -34.515 ;
        RECT -57.285 -36.205 -56.955 -35.875 ;
        RECT -57.285 -37.565 -56.955 -37.235 ;
        RECT -57.285 -38.925 -56.955 -38.595 ;
        RECT -57.285 -40.285 -56.955 -39.955 ;
        RECT -57.285 -41.645 -56.955 -41.315 ;
        RECT -57.285 -43.005 -56.955 -42.675 ;
        RECT -57.285 -44.365 -56.955 -44.035 ;
        RECT -57.285 -45.725 -56.955 -45.395 ;
        RECT -57.285 -47.085 -56.955 -46.755 ;
        RECT -57.285 -48.445 -56.955 -48.115 ;
        RECT -57.285 -49.805 -56.955 -49.475 ;
        RECT -57.285 -51.165 -56.955 -50.835 ;
        RECT -57.285 -52.525 -56.955 -52.195 ;
        RECT -57.285 -53.885 -56.955 -53.555 ;
        RECT -57.285 -55.245 -56.955 -54.915 ;
        RECT -57.285 -56.605 -56.955 -56.275 ;
        RECT -57.285 -57.965 -56.955 -57.635 ;
        RECT -57.285 -59.325 -56.955 -58.995 ;
        RECT -57.285 -60.685 -56.955 -60.355 ;
        RECT -57.285 -62.045 -56.955 -61.715 ;
        RECT -57.285 -63.405 -56.955 -63.075 ;
        RECT -57.285 -64.765 -56.955 -64.435 ;
        RECT -57.285 -66.125 -56.955 -65.795 ;
        RECT -57.285 -67.485 -56.955 -67.155 ;
        RECT -57.285 -68.845 -56.955 -68.515 ;
        RECT -57.285 -70.205 -56.955 -69.875 ;
        RECT -57.285 -71.565 -56.955 -71.235 ;
        RECT -57.285 -72.925 -56.955 -72.595 ;
        RECT -57.285 -74.285 -56.955 -73.955 ;
        RECT -57.285 -75.645 -56.955 -75.315 ;
        RECT -57.285 -77.005 -56.955 -76.675 ;
        RECT -57.285 -78.365 -56.955 -78.035 ;
        RECT -57.285 -79.725 -56.955 -79.395 ;
        RECT -57.285 -81.085 -56.955 -80.755 ;
        RECT -57.285 -82.445 -56.955 -82.115 ;
        RECT -57.285 -83.805 -56.955 -83.475 ;
        RECT -57.285 -85.165 -56.955 -84.835 ;
        RECT -57.285 -86.525 -56.955 -86.195 ;
        RECT -57.285 -87.885 -56.955 -87.555 ;
        RECT -57.285 -89.245 -56.955 -88.915 ;
        RECT -57.285 -90.605 -56.955 -90.275 ;
        RECT -57.285 -91.965 -56.955 -91.635 ;
        RECT -57.285 -93.325 -56.955 -92.995 ;
        RECT -57.285 -94.685 -56.955 -94.355 ;
        RECT -57.285 -96.045 -56.955 -95.715 ;
        RECT -57.285 -97.405 -56.955 -97.075 ;
        RECT -57.285 -98.765 -56.955 -98.435 ;
        RECT -57.285 -100.125 -56.955 -99.795 ;
        RECT -57.285 -101.485 -56.955 -101.155 ;
        RECT -57.285 -102.845 -56.955 -102.515 ;
        RECT -57.285 -104.205 -56.955 -103.875 ;
        RECT -57.285 -105.565 -56.955 -105.235 ;
        RECT -57.285 -106.925 -56.955 -106.595 ;
        RECT -57.285 -108.285 -56.955 -107.955 ;
        RECT -57.285 -109.645 -56.955 -109.315 ;
        RECT -57.285 -111.005 -56.955 -110.675 ;
        RECT -57.285 -112.365 -56.955 -112.035 ;
        RECT -57.285 -113.725 -56.955 -113.395 ;
        RECT -57.285 -115.085 -56.955 -114.755 ;
        RECT -57.285 -116.445 -56.955 -116.115 ;
        RECT -57.285 -117.805 -56.955 -117.475 ;
        RECT -57.285 -119.165 -56.955 -118.835 ;
        RECT -57.285 -120.525 -56.955 -120.195 ;
        RECT -57.285 -121.885 -56.955 -121.555 ;
        RECT -57.285 -123.245 -56.955 -122.915 ;
        RECT -57.285 -124.605 -56.955 -124.275 ;
        RECT -57.285 -125.965 -56.955 -125.635 ;
        RECT -57.285 -127.325 -56.955 -126.995 ;
        RECT -57.285 -128.685 -56.955 -128.355 ;
        RECT -57.285 -130.045 -56.955 -129.715 ;
        RECT -57.285 -131.405 -56.955 -131.075 ;
        RECT -57.285 -134.125 -56.955 -133.795 ;
        RECT -57.285 -135.485 -56.955 -135.155 ;
        RECT -57.285 -136.845 -56.955 -136.515 ;
        RECT -57.285 -138.205 -56.955 -137.875 ;
        RECT -57.285 -139.565 -56.955 -139.235 ;
        RECT -57.285 -140.925 -56.955 -140.595 ;
        RECT -57.285 -142.285 -56.955 -141.955 ;
        RECT -57.285 -143.645 -56.955 -143.315 ;
        RECT -57.285 -145.005 -56.955 -144.675 ;
        RECT -57.285 -146.365 -56.955 -146.035 ;
        RECT -57.285 -147.725 -56.955 -147.395 ;
        RECT -57.285 -149.085 -56.955 -148.755 ;
        RECT -57.285 -150.445 -56.955 -150.115 ;
        RECT -57.285 -151.805 -56.955 -151.475 ;
        RECT -57.285 -153.165 -56.955 -152.835 ;
        RECT -57.285 -154.525 -56.955 -154.195 ;
        RECT -57.285 -155.885 -56.955 -155.555 ;
        RECT -57.285 -157.245 -56.955 -156.915 ;
        RECT -57.285 -158.605 -56.955 -158.275 ;
        RECT -57.285 -159.965 -56.955 -159.635 ;
        RECT -57.285 -161.325 -56.955 -160.995 ;
        RECT -57.285 -162.685 -56.955 -162.355 ;
        RECT -57.285 -164.045 -56.955 -163.715 ;
        RECT -57.285 -165.405 -56.955 -165.075 ;
        RECT -57.285 -166.765 -56.955 -166.435 ;
        RECT -57.285 -168.125 -56.955 -167.795 ;
        RECT -57.285 -169.485 -56.955 -169.155 ;
        RECT -57.285 -170.845 -56.955 -170.515 ;
        RECT -57.285 -172.205 -56.955 -171.875 ;
        RECT -57.285 -173.565 -56.955 -173.235 ;
        RECT -57.285 -174.925 -56.955 -174.595 ;
        RECT -57.285 -176.285 -56.955 -175.955 ;
        RECT -57.285 -177.645 -56.955 -177.315 ;
        RECT -57.285 -179.005 -56.955 -178.675 ;
        RECT -57.285 -180.365 -56.955 -180.035 ;
        RECT -57.285 -181.725 -56.955 -181.395 ;
        RECT -57.285 -183.085 -56.955 -182.755 ;
        RECT -57.285 -184.445 -56.955 -184.115 ;
        RECT -57.285 -185.805 -56.955 -185.475 ;
        RECT -57.285 -187.165 -56.955 -186.835 ;
        RECT -57.285 -188.525 -56.955 -188.195 ;
        RECT -57.285 -189.885 -56.955 -189.555 ;
        RECT -57.285 -191.245 -56.955 -190.915 ;
        RECT -57.285 -192.605 -56.955 -192.275 ;
        RECT -57.285 -193.965 -56.955 -193.635 ;
        RECT -57.285 -195.325 -56.955 -194.995 ;
        RECT -57.285 -196.685 -56.955 -196.355 ;
        RECT -57.285 -198.045 -56.955 -197.715 ;
        RECT -57.285 -199.405 -56.955 -199.075 ;
        RECT -57.285 -200.765 -56.955 -200.435 ;
        RECT -57.285 -202.125 -56.955 -201.795 ;
        RECT -57.285 -203.485 -56.955 -203.155 ;
        RECT -57.285 -204.845 -56.955 -204.515 ;
        RECT -57.285 -206.555 -56.955 -206.225 ;
        RECT -57.285 -207.565 -56.955 -207.235 ;
        RECT -57.285 -208.925 -56.955 -208.595 ;
        RECT -57.285 -211.645 -56.955 -211.315 ;
        RECT -57.285 -214.365 -56.955 -214.035 ;
        RECT -57.285 -215.725 -56.955 -215.395 ;
        RECT -57.285 -217.085 -56.955 -216.755 ;
        RECT -57.285 -218.445 -56.955 -218.115 ;
        RECT -57.285 -224.09 -56.955 -222.96 ;
        RECT -57.28 -224.205 -56.96 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -55.925 -15.805 -55.595 -15.475 ;
        RECT -55.925 -17.165 -55.595 -16.835 ;
        RECT -55.925 -18.525 -55.595 -18.195 ;
        RECT -55.925 -19.885 -55.595 -19.555 ;
        RECT -55.925 -21.245 -55.595 -20.915 ;
        RECT -55.925 -22.605 -55.595 -22.275 ;
        RECT -55.925 -23.965 -55.595 -23.635 ;
        RECT -55.925 -25.325 -55.595 -24.995 ;
        RECT -55.925 -26.685 -55.595 -26.355 ;
        RECT -55.925 -28.045 -55.595 -27.715 ;
        RECT -55.925 -29.405 -55.595 -29.075 ;
        RECT -55.925 -30.765 -55.595 -30.435 ;
        RECT -55.925 -32.125 -55.595 -31.795 ;
        RECT -55.925 -33.485 -55.595 -33.155 ;
        RECT -55.925 -34.845 -55.595 -34.515 ;
        RECT -55.925 -36.205 -55.595 -35.875 ;
        RECT -55.925 -37.565 -55.595 -37.235 ;
        RECT -55.925 -38.925 -55.595 -38.595 ;
        RECT -55.925 -40.285 -55.595 -39.955 ;
        RECT -55.925 -41.645 -55.595 -41.315 ;
        RECT -55.925 -43.005 -55.595 -42.675 ;
        RECT -55.925 -44.365 -55.595 -44.035 ;
        RECT -55.925 -45.725 -55.595 -45.395 ;
        RECT -55.925 -47.085 -55.595 -46.755 ;
        RECT -55.925 -48.445 -55.595 -48.115 ;
        RECT -55.925 -49.805 -55.595 -49.475 ;
        RECT -55.925 -51.165 -55.595 -50.835 ;
        RECT -55.925 -52.525 -55.595 -52.195 ;
        RECT -55.925 -53.885 -55.595 -53.555 ;
        RECT -55.925 -55.245 -55.595 -54.915 ;
        RECT -55.925 -56.605 -55.595 -56.275 ;
        RECT -55.925 -57.965 -55.595 -57.635 ;
        RECT -55.925 -59.325 -55.595 -58.995 ;
        RECT -55.925 -60.685 -55.595 -60.355 ;
        RECT -55.925 -62.045 -55.595 -61.715 ;
        RECT -55.925 -63.405 -55.595 -63.075 ;
        RECT -55.925 -64.765 -55.595 -64.435 ;
        RECT -55.925 -66.125 -55.595 -65.795 ;
        RECT -55.925 -67.485 -55.595 -67.155 ;
        RECT -55.925 -68.845 -55.595 -68.515 ;
        RECT -55.925 -70.205 -55.595 -69.875 ;
        RECT -55.925 -71.565 -55.595 -71.235 ;
        RECT -55.925 -72.925 -55.595 -72.595 ;
        RECT -55.925 -74.285 -55.595 -73.955 ;
        RECT -55.925 -75.645 -55.595 -75.315 ;
        RECT -55.925 -77.005 -55.595 -76.675 ;
        RECT -55.925 -78.365 -55.595 -78.035 ;
        RECT -55.925 -79.725 -55.595 -79.395 ;
        RECT -55.925 -81.085 -55.595 -80.755 ;
        RECT -55.925 -82.445 -55.595 -82.115 ;
        RECT -55.925 -83.805 -55.595 -83.475 ;
        RECT -55.925 -85.165 -55.595 -84.835 ;
        RECT -55.925 -86.525 -55.595 -86.195 ;
        RECT -55.925 -87.885 -55.595 -87.555 ;
        RECT -55.925 -89.245 -55.595 -88.915 ;
        RECT -55.925 -90.605 -55.595 -90.275 ;
        RECT -55.925 -91.965 -55.595 -91.635 ;
        RECT -55.925 -93.325 -55.595 -92.995 ;
        RECT -55.925 -94.685 -55.595 -94.355 ;
        RECT -55.925 -96.045 -55.595 -95.715 ;
        RECT -55.925 -97.405 -55.595 -97.075 ;
        RECT -55.925 -98.765 -55.595 -98.435 ;
        RECT -55.925 -100.125 -55.595 -99.795 ;
        RECT -55.925 -101.485 -55.595 -101.155 ;
        RECT -55.925 -102.845 -55.595 -102.515 ;
        RECT -55.925 -104.205 -55.595 -103.875 ;
        RECT -55.925 -105.565 -55.595 -105.235 ;
        RECT -55.925 -106.925 -55.595 -106.595 ;
        RECT -55.925 -108.285 -55.595 -107.955 ;
        RECT -55.925 -109.645 -55.595 -109.315 ;
        RECT -55.925 -111.005 -55.595 -110.675 ;
        RECT -55.925 -111.87 -55.595 -111.54 ;
        RECT -55.925 -113.725 -55.595 -113.395 ;
        RECT -55.925 -115.085 -55.595 -114.755 ;
        RECT -55.925 -116.445 -55.595 -116.115 ;
        RECT -55.925 -117.805 -55.595 -117.475 ;
        RECT -55.925 -120.525 -55.595 -120.195 ;
        RECT -55.925 -121.885 -55.595 -121.555 ;
        RECT -55.925 -123.245 -55.595 -122.915 ;
        RECT -55.925 -124.71 -55.595 -124.38 ;
        RECT -55.925 -125.965 -55.595 -125.635 ;
        RECT -55.925 -127.325 -55.595 -126.995 ;
        RECT -55.925 -130.045 -55.595 -129.715 ;
        RECT -55.925 -134.125 -55.595 -133.795 ;
        RECT -55.925 -135.485 -55.595 -135.155 ;
        RECT -55.925 -136.845 -55.595 -136.515 ;
        RECT -55.925 -138.205 -55.595 -137.875 ;
        RECT -55.925 -139.565 -55.595 -139.235 ;
        RECT -55.925 -142.285 -55.595 -141.955 ;
        RECT -55.925 -143.645 -55.595 -143.315 ;
        RECT -55.925 -145.005 -55.595 -144.675 ;
        RECT -55.925 -146.365 -55.595 -146.035 ;
        RECT -55.925 -147.725 -55.595 -147.395 ;
        RECT -55.925 -149.085 -55.595 -148.755 ;
        RECT -55.925 -150.445 -55.595 -150.115 ;
        RECT -55.925 -151.805 -55.595 -151.475 ;
        RECT -55.925 -153.165 -55.595 -152.835 ;
        RECT -55.925 -154.525 -55.595 -154.195 ;
        RECT -55.925 -155.885 -55.595 -155.555 ;
        RECT -55.925 -157.245 -55.595 -156.915 ;
        RECT -55.925 -158.605 -55.595 -158.275 ;
        RECT -55.925 -159.965 -55.595 -159.635 ;
        RECT -55.925 -161.325 -55.595 -160.995 ;
        RECT -55.925 -162.685 -55.595 -162.355 ;
        RECT -55.925 -164.045 -55.595 -163.715 ;
        RECT -55.925 -165.405 -55.595 -165.075 ;
        RECT -55.925 -166.765 -55.595 -166.435 ;
        RECT -55.925 -168.125 -55.595 -167.795 ;
        RECT -55.925 -169.485 -55.595 -169.155 ;
        RECT -55.925 -170.845 -55.595 -170.515 ;
        RECT -55.925 -172.205 -55.595 -171.875 ;
        RECT -55.925 -173.565 -55.595 -173.235 ;
        RECT -55.925 -174.925 -55.595 -174.595 ;
        RECT -55.925 -176.285 -55.595 -175.955 ;
        RECT -55.925 -177.645 -55.595 -177.315 ;
        RECT -55.925 -179.005 -55.595 -178.675 ;
        RECT -55.925 -180.365 -55.595 -180.035 ;
        RECT -55.925 -181.725 -55.595 -181.395 ;
        RECT -55.925 -183.085 -55.595 -182.755 ;
        RECT -55.925 -184.445 -55.595 -184.115 ;
        RECT -55.925 -185.805 -55.595 -185.475 ;
        RECT -55.925 -187.165 -55.595 -186.835 ;
        RECT -55.925 -188.525 -55.595 -188.195 ;
        RECT -55.925 -189.885 -55.595 -189.555 ;
        RECT -55.925 -191.245 -55.595 -190.915 ;
        RECT -55.925 -192.605 -55.595 -192.275 ;
        RECT -55.925 -193.965 -55.595 -193.635 ;
        RECT -55.925 -195.325 -55.595 -194.995 ;
        RECT -55.925 -196.685 -55.595 -196.355 ;
        RECT -55.925 -198.045 -55.595 -197.715 ;
        RECT -55.925 -199.405 -55.595 -199.075 ;
        RECT -55.925 -200.765 -55.595 -200.435 ;
        RECT -55.925 -202.125 -55.595 -201.795 ;
        RECT -55.925 -203.485 -55.595 -203.155 ;
        RECT -55.925 -204.845 -55.595 -204.515 ;
        RECT -55.925 -206.555 -55.595 -206.225 ;
        RECT -55.925 -207.565 -55.595 -207.235 ;
        RECT -55.925 -208.925 -55.595 -208.595 ;
        RECT -55.925 -210.285 -55.595 -209.955 ;
        RECT -55.925 -211.645 -55.595 -211.315 ;
        RECT -55.925 -214.365 -55.595 -214.035 ;
        RECT -55.925 -215.725 -55.595 -215.395 ;
        RECT -55.925 -217.085 -55.595 -216.755 ;
        RECT -55.925 -218.445 -55.595 -218.115 ;
        RECT -55.925 -224.09 -55.595 -222.96 ;
        RECT -55.92 -224.205 -55.6 133.765 ;
        RECT -55.925 132.52 -55.595 133.65 ;
        RECT -55.925 128.355 -55.595 128.685 ;
        RECT -55.925 126.995 -55.595 127.325 ;
        RECT -55.925 125.635 -55.595 125.965 ;
        RECT -55.925 124.275 -55.595 124.605 ;
        RECT -55.925 122.915 -55.595 123.245 ;
        RECT -55.925 121.555 -55.595 121.885 ;
        RECT -55.925 120.195 -55.595 120.525 ;
        RECT -55.925 118.835 -55.595 119.165 ;
        RECT -55.925 117.475 -55.595 117.805 ;
        RECT -55.925 116.115 -55.595 116.445 ;
        RECT -55.925 114.755 -55.595 115.085 ;
        RECT -55.925 113.395 -55.595 113.725 ;
        RECT -55.925 112.035 -55.595 112.365 ;
        RECT -55.925 110.675 -55.595 111.005 ;
        RECT -55.925 109.315 -55.595 109.645 ;
        RECT -55.925 107.955 -55.595 108.285 ;
        RECT -55.925 106.595 -55.595 106.925 ;
        RECT -55.925 105.235 -55.595 105.565 ;
        RECT -55.925 103.875 -55.595 104.205 ;
        RECT -55.925 102.515 -55.595 102.845 ;
        RECT -55.925 101.155 -55.595 101.485 ;
        RECT -55.925 99.795 -55.595 100.125 ;
        RECT -55.925 98.435 -55.595 98.765 ;
        RECT -55.925 97.075 -55.595 97.405 ;
        RECT -55.925 95.715 -55.595 96.045 ;
        RECT -55.925 94.355 -55.595 94.685 ;
        RECT -55.925 92.995 -55.595 93.325 ;
        RECT -55.925 91.635 -55.595 91.965 ;
        RECT -55.925 90.275 -55.595 90.605 ;
        RECT -55.925 88.915 -55.595 89.245 ;
        RECT -55.925 87.555 -55.595 87.885 ;
        RECT -55.925 86.195 -55.595 86.525 ;
        RECT -55.925 84.835 -55.595 85.165 ;
        RECT -55.925 83.475 -55.595 83.805 ;
        RECT -55.925 82.115 -55.595 82.445 ;
        RECT -55.925 80.755 -55.595 81.085 ;
        RECT -55.925 79.395 -55.595 79.725 ;
        RECT -55.925 78.035 -55.595 78.365 ;
        RECT -55.925 76.675 -55.595 77.005 ;
        RECT -55.925 75.315 -55.595 75.645 ;
        RECT -55.925 73.955 -55.595 74.285 ;
        RECT -55.925 71.64 -55.595 71.97 ;
        RECT -55.925 69.465 -55.595 69.795 ;
        RECT -55.925 68.615 -55.595 68.945 ;
        RECT -55.925 66.305 -55.595 66.635 ;
        RECT -55.925 65.455 -55.595 65.785 ;
        RECT -55.925 63.145 -55.595 63.475 ;
        RECT -55.925 62.295 -55.595 62.625 ;
        RECT -55.925 59.985 -55.595 60.315 ;
        RECT -55.925 59.135 -55.595 59.465 ;
        RECT -55.925 56.825 -55.595 57.155 ;
        RECT -55.925 55.975 -55.595 56.305 ;
        RECT -55.925 53.665 -55.595 53.995 ;
        RECT -55.925 52.815 -55.595 53.145 ;
        RECT -55.925 50.64 -55.595 50.97 ;
        RECT -55.925 48.115 -55.595 48.445 ;
        RECT -55.925 46.755 -55.595 47.085 ;
        RECT -55.925 45.395 -55.595 45.725 ;
        RECT -55.925 44.035 -55.595 44.365 ;
        RECT -55.925 42.675 -55.595 43.005 ;
        RECT -55.925 41.315 -55.595 41.645 ;
        RECT -55.925 39.955 -55.595 40.285 ;
        RECT -55.925 38.595 -55.595 38.925 ;
        RECT -55.925 37.235 -55.595 37.565 ;
        RECT -55.925 35.875 -55.595 36.205 ;
        RECT -55.925 34.515 -55.595 34.845 ;
        RECT -55.925 33.155 -55.595 33.485 ;
        RECT -55.925 31.795 -55.595 32.125 ;
        RECT -55.925 30.435 -55.595 30.765 ;
        RECT -55.925 29.075 -55.595 29.405 ;
        RECT -55.925 27.715 -55.595 28.045 ;
        RECT -55.925 26.355 -55.595 26.685 ;
        RECT -55.925 24.995 -55.595 25.325 ;
        RECT -55.925 23.635 -55.595 23.965 ;
        RECT -55.925 22.275 -55.595 22.605 ;
        RECT -55.925 20.915 -55.595 21.245 ;
        RECT -55.925 19.555 -55.595 19.885 ;
        RECT -55.925 18.195 -55.595 18.525 ;
        RECT -55.925 16.835 -55.595 17.165 ;
        RECT -55.925 15.475 -55.595 15.805 ;
        RECT -55.925 14.115 -55.595 14.445 ;
        RECT -55.925 12.755 -55.595 13.085 ;
        RECT -55.925 11.395 -55.595 11.725 ;
        RECT -55.925 10.035 -55.595 10.365 ;
        RECT -55.925 8.675 -55.595 9.005 ;
        RECT -55.925 7.315 -55.595 7.645 ;
        RECT -55.925 5.955 -55.595 6.285 ;
        RECT -55.925 4.595 -55.595 4.925 ;
        RECT -55.925 3.235 -55.595 3.565 ;
        RECT -55.925 1.875 -55.595 2.205 ;
        RECT -55.925 0.515 -55.595 0.845 ;
        RECT -55.925 -0.845 -55.595 -0.515 ;
        RECT -55.925 -2.205 -55.595 -1.875 ;
        RECT -55.925 -3.565 -55.595 -3.235 ;
        RECT -55.925 -4.925 -55.595 -4.595 ;
        RECT -55.925 -6.285 -55.595 -5.955 ;
        RECT -55.925 -7.645 -55.595 -7.315 ;
        RECT -55.925 -9.005 -55.595 -8.675 ;
        RECT -55.925 -10.365 -55.595 -10.035 ;
        RECT -55.925 -11.725 -55.595 -11.395 ;
        RECT -55.925 -13.085 -55.595 -12.755 ;
        RECT -55.925 -14.445 -55.595 -14.115 ;
    END
    PORT
      LAYER met3 ;
        RECT -65.445 132.52 -65.115 133.65 ;
        RECT -65.445 128.355 -65.115 128.685 ;
        RECT -65.445 126.995 -65.115 127.325 ;
        RECT -65.445 125.635 -65.115 125.965 ;
        RECT -65.445 124.275 -65.115 124.605 ;
        RECT -65.445 122.915 -65.115 123.245 ;
        RECT -65.445 121.555 -65.115 121.885 ;
        RECT -65.445 120.195 -65.115 120.525 ;
        RECT -65.445 118.835 -65.115 119.165 ;
        RECT -65.445 117.475 -65.115 117.805 ;
        RECT -65.445 116.115 -65.115 116.445 ;
        RECT -65.445 114.755 -65.115 115.085 ;
        RECT -65.445 113.395 -65.115 113.725 ;
        RECT -65.445 112.035 -65.115 112.365 ;
        RECT -65.445 110.675 -65.115 111.005 ;
        RECT -65.445 109.315 -65.115 109.645 ;
        RECT -65.445 107.955 -65.115 108.285 ;
        RECT -65.445 106.595 -65.115 106.925 ;
        RECT -65.445 105.235 -65.115 105.565 ;
        RECT -65.445 103.875 -65.115 104.205 ;
        RECT -65.445 102.515 -65.115 102.845 ;
        RECT -65.445 101.155 -65.115 101.485 ;
        RECT -65.445 99.795 -65.115 100.125 ;
        RECT -65.445 98.435 -65.115 98.765 ;
        RECT -65.445 97.075 -65.115 97.405 ;
        RECT -65.445 95.715 -65.115 96.045 ;
        RECT -65.445 94.355 -65.115 94.685 ;
        RECT -65.445 92.995 -65.115 93.325 ;
        RECT -65.445 91.635 -65.115 91.965 ;
        RECT -65.445 90.275 -65.115 90.605 ;
        RECT -65.445 88.915 -65.115 89.245 ;
        RECT -65.445 87.555 -65.115 87.885 ;
        RECT -65.445 86.195 -65.115 86.525 ;
        RECT -65.445 84.835 -65.115 85.165 ;
        RECT -65.445 83.475 -65.115 83.805 ;
        RECT -65.445 82.115 -65.115 82.445 ;
        RECT -65.445 80.755 -65.115 81.085 ;
        RECT -65.445 79.395 -65.115 79.725 ;
        RECT -65.445 78.035 -65.115 78.365 ;
        RECT -65.445 76.675 -65.115 77.005 ;
        RECT -65.445 75.315 -65.115 75.645 ;
        RECT -65.445 73.955 -65.115 74.285 ;
        RECT -65.445 72.595 -65.115 72.925 ;
        RECT -65.445 71.235 -65.115 71.565 ;
        RECT -65.445 69.875 -65.115 70.205 ;
        RECT -65.445 68.515 -65.115 68.845 ;
        RECT -65.445 67.155 -65.115 67.485 ;
        RECT -65.445 65.795 -65.115 66.125 ;
        RECT -65.445 64.435 -65.115 64.765 ;
        RECT -65.445 63.075 -65.115 63.405 ;
        RECT -65.445 61.715 -65.115 62.045 ;
        RECT -65.445 60.355 -65.115 60.685 ;
        RECT -65.445 58.995 -65.115 59.325 ;
        RECT -65.445 57.635 -65.115 57.965 ;
        RECT -65.445 56.275 -65.115 56.605 ;
        RECT -65.445 54.915 -65.115 55.245 ;
        RECT -65.445 53.555 -65.115 53.885 ;
        RECT -65.445 52.195 -65.115 52.525 ;
        RECT -65.445 50.835 -65.115 51.165 ;
        RECT -65.445 49.475 -65.115 49.805 ;
        RECT -65.445 48.115 -65.115 48.445 ;
        RECT -65.445 46.755 -65.115 47.085 ;
        RECT -65.445 45.395 -65.115 45.725 ;
        RECT -65.445 44.035 -65.115 44.365 ;
        RECT -65.445 42.675 -65.115 43.005 ;
        RECT -65.445 41.315 -65.115 41.645 ;
        RECT -65.445 39.955 -65.115 40.285 ;
        RECT -65.445 38.595 -65.115 38.925 ;
        RECT -65.445 37.235 -65.115 37.565 ;
        RECT -65.445 35.875 -65.115 36.205 ;
        RECT -65.445 34.515 -65.115 34.845 ;
        RECT -65.445 33.155 -65.115 33.485 ;
        RECT -65.445 31.795 -65.115 32.125 ;
        RECT -65.445 30.435 -65.115 30.765 ;
        RECT -65.445 29.075 -65.115 29.405 ;
        RECT -65.445 27.715 -65.115 28.045 ;
        RECT -65.445 26.355 -65.115 26.685 ;
        RECT -65.445 24.995 -65.115 25.325 ;
        RECT -65.445 23.635 -65.115 23.965 ;
        RECT -65.445 22.275 -65.115 22.605 ;
        RECT -65.445 20.915 -65.115 21.245 ;
        RECT -65.445 19.555 -65.115 19.885 ;
        RECT -65.445 18.195 -65.115 18.525 ;
        RECT -65.445 16.835 -65.115 17.165 ;
        RECT -65.445 15.475 -65.115 15.805 ;
        RECT -65.445 14.115 -65.115 14.445 ;
        RECT -65.445 12.755 -65.115 13.085 ;
        RECT -65.445 11.395 -65.115 11.725 ;
        RECT -65.445 10.035 -65.115 10.365 ;
        RECT -65.445 8.675 -65.115 9.005 ;
        RECT -65.445 7.315 -65.115 7.645 ;
        RECT -65.445 5.955 -65.115 6.285 ;
        RECT -65.445 4.595 -65.115 4.925 ;
        RECT -65.445 3.235 -65.115 3.565 ;
        RECT -65.445 1.875 -65.115 2.205 ;
        RECT -65.445 0.515 -65.115 0.845 ;
        RECT -65.445 -0.845 -65.115 -0.515 ;
        RECT -65.445 -2.205 -65.115 -1.875 ;
        RECT -65.445 -3.565 -65.115 -3.235 ;
        RECT -65.445 -4.925 -65.115 -4.595 ;
        RECT -65.445 -6.285 -65.115 -5.955 ;
        RECT -65.445 -7.645 -65.115 -7.315 ;
        RECT -65.445 -9.005 -65.115 -8.675 ;
        RECT -65.445 -10.365 -65.115 -10.035 ;
        RECT -65.445 -11.725 -65.115 -11.395 ;
        RECT -65.445 -13.085 -65.115 -12.755 ;
        RECT -65.445 -14.445 -65.115 -14.115 ;
        RECT -65.445 -15.805 -65.115 -15.475 ;
        RECT -65.445 -17.165 -65.115 -16.835 ;
        RECT -65.445 -18.525 -65.115 -18.195 ;
        RECT -65.445 -19.885 -65.115 -19.555 ;
        RECT -65.445 -21.245 -65.115 -20.915 ;
        RECT -65.445 -22.605 -65.115 -22.275 ;
        RECT -65.445 -23.965 -65.115 -23.635 ;
        RECT -65.445 -25.325 -65.115 -24.995 ;
        RECT -65.445 -26.685 -65.115 -26.355 ;
        RECT -65.445 -28.045 -65.115 -27.715 ;
        RECT -65.445 -29.405 -65.115 -29.075 ;
        RECT -65.445 -30.765 -65.115 -30.435 ;
        RECT -65.445 -32.125 -65.115 -31.795 ;
        RECT -65.445 -33.485 -65.115 -33.155 ;
        RECT -65.445 -34.845 -65.115 -34.515 ;
        RECT -65.445 -36.205 -65.115 -35.875 ;
        RECT -65.445 -37.565 -65.115 -37.235 ;
        RECT -65.445 -38.925 -65.115 -38.595 ;
        RECT -65.445 -40.285 -65.115 -39.955 ;
        RECT -65.445 -41.645 -65.115 -41.315 ;
        RECT -65.445 -43.005 -65.115 -42.675 ;
        RECT -65.445 -44.365 -65.115 -44.035 ;
        RECT -65.445 -45.725 -65.115 -45.395 ;
        RECT -65.445 -47.085 -65.115 -46.755 ;
        RECT -65.445 -48.445 -65.115 -48.115 ;
        RECT -65.445 -49.805 -65.115 -49.475 ;
        RECT -65.445 -51.165 -65.115 -50.835 ;
        RECT -65.445 -52.525 -65.115 -52.195 ;
        RECT -65.445 -53.885 -65.115 -53.555 ;
        RECT -65.445 -55.245 -65.115 -54.915 ;
        RECT -65.445 -56.605 -65.115 -56.275 ;
        RECT -65.445 -57.965 -65.115 -57.635 ;
        RECT -65.445 -59.325 -65.115 -58.995 ;
        RECT -65.445 -60.685 -65.115 -60.355 ;
        RECT -65.445 -62.045 -65.115 -61.715 ;
        RECT -65.445 -63.405 -65.115 -63.075 ;
        RECT -65.445 -64.765 -65.115 -64.435 ;
        RECT -65.445 -66.125 -65.115 -65.795 ;
        RECT -65.445 -67.485 -65.115 -67.155 ;
        RECT -65.445 -68.845 -65.115 -68.515 ;
        RECT -65.445 -70.205 -65.115 -69.875 ;
        RECT -65.445 -71.565 -65.115 -71.235 ;
        RECT -65.445 -72.925 -65.115 -72.595 ;
        RECT -65.445 -74.285 -65.115 -73.955 ;
        RECT -65.445 -75.645 -65.115 -75.315 ;
        RECT -65.445 -77.005 -65.115 -76.675 ;
        RECT -65.445 -78.365 -65.115 -78.035 ;
        RECT -65.445 -79.725 -65.115 -79.395 ;
        RECT -65.445 -81.085 -65.115 -80.755 ;
        RECT -65.445 -82.445 -65.115 -82.115 ;
        RECT -65.445 -83.805 -65.115 -83.475 ;
        RECT -65.445 -85.165 -65.115 -84.835 ;
        RECT -65.445 -86.525 -65.115 -86.195 ;
        RECT -65.445 -87.885 -65.115 -87.555 ;
        RECT -65.445 -89.245 -65.115 -88.915 ;
        RECT -65.445 -90.605 -65.115 -90.275 ;
        RECT -65.445 -91.965 -65.115 -91.635 ;
        RECT -65.445 -93.325 -65.115 -92.995 ;
        RECT -65.445 -94.685 -65.115 -94.355 ;
        RECT -65.445 -96.045 -65.115 -95.715 ;
        RECT -65.445 -97.405 -65.115 -97.075 ;
        RECT -65.445 -98.765 -65.115 -98.435 ;
        RECT -65.445 -100.125 -65.115 -99.795 ;
        RECT -65.445 -101.485 -65.115 -101.155 ;
        RECT -65.445 -102.845 -65.115 -102.515 ;
        RECT -65.445 -104.205 -65.115 -103.875 ;
        RECT -65.445 -105.565 -65.115 -105.235 ;
        RECT -65.445 -106.925 -65.115 -106.595 ;
        RECT -65.445 -108.285 -65.115 -107.955 ;
        RECT -65.445 -109.645 -65.115 -109.315 ;
        RECT -65.445 -111.005 -65.115 -110.675 ;
        RECT -65.445 -112.365 -65.115 -112.035 ;
        RECT -65.445 -113.725 -65.115 -113.395 ;
        RECT -65.445 -115.085 -65.115 -114.755 ;
        RECT -65.445 -116.445 -65.115 -116.115 ;
        RECT -65.445 -117.805 -65.115 -117.475 ;
        RECT -65.445 -119.165 -65.115 -118.835 ;
        RECT -65.445 -120.525 -65.115 -120.195 ;
        RECT -65.445 -121.885 -65.115 -121.555 ;
        RECT -65.445 -123.245 -65.115 -122.915 ;
        RECT -65.445 -124.605 -65.115 -124.275 ;
        RECT -65.445 -125.965 -65.115 -125.635 ;
        RECT -65.445 -127.325 -65.115 -126.995 ;
        RECT -65.445 -128.685 -65.115 -128.355 ;
        RECT -65.445 -130.045 -65.115 -129.715 ;
        RECT -65.445 -131.405 -65.115 -131.075 ;
        RECT -65.445 -132.765 -65.115 -132.435 ;
        RECT -65.445 -134.125 -65.115 -133.795 ;
        RECT -65.445 -135.485 -65.115 -135.155 ;
        RECT -65.445 -136.845 -65.115 -136.515 ;
        RECT -65.445 -138.205 -65.115 -137.875 ;
        RECT -65.445 -139.565 -65.115 -139.235 ;
        RECT -65.445 -140.925 -65.115 -140.595 ;
        RECT -65.445 -142.285 -65.115 -141.955 ;
        RECT -65.445 -143.645 -65.115 -143.315 ;
        RECT -65.445 -145.005 -65.115 -144.675 ;
        RECT -65.445 -146.365 -65.115 -146.035 ;
        RECT -65.445 -147.725 -65.115 -147.395 ;
        RECT -65.445 -149.085 -65.115 -148.755 ;
        RECT -65.445 -150.445 -65.115 -150.115 ;
        RECT -65.445 -151.805 -65.115 -151.475 ;
        RECT -65.445 -153.165 -65.115 -152.835 ;
        RECT -65.445 -154.525 -65.115 -154.195 ;
        RECT -65.445 -155.885 -65.115 -155.555 ;
        RECT -65.445 -157.245 -65.115 -156.915 ;
        RECT -65.445 -158.605 -65.115 -158.275 ;
        RECT -65.445 -159.965 -65.115 -159.635 ;
        RECT -65.445 -161.325 -65.115 -160.995 ;
        RECT -65.445 -162.685 -65.115 -162.355 ;
        RECT -65.445 -164.045 -65.115 -163.715 ;
        RECT -65.445 -165.405 -65.115 -165.075 ;
        RECT -65.445 -166.765 -65.115 -166.435 ;
        RECT -65.445 -168.125 -65.115 -167.795 ;
        RECT -65.445 -169.485 -65.115 -169.155 ;
        RECT -65.445 -170.845 -65.115 -170.515 ;
        RECT -65.445 -172.205 -65.115 -171.875 ;
        RECT -65.445 -173.565 -65.115 -173.235 ;
        RECT -65.445 -174.925 -65.115 -174.595 ;
        RECT -65.445 -176.285 -65.115 -175.955 ;
        RECT -65.445 -177.645 -65.115 -177.315 ;
        RECT -65.445 -179.005 -65.115 -178.675 ;
        RECT -65.445 -180.365 -65.115 -180.035 ;
        RECT -65.445 -181.725 -65.115 -181.395 ;
        RECT -65.445 -183.085 -65.115 -182.755 ;
        RECT -65.445 -184.445 -65.115 -184.115 ;
        RECT -65.445 -185.805 -65.115 -185.475 ;
        RECT -65.445 -187.165 -65.115 -186.835 ;
        RECT -65.445 -188.525 -65.115 -188.195 ;
        RECT -65.445 -189.885 -65.115 -189.555 ;
        RECT -65.445 -191.245 -65.115 -190.915 ;
        RECT -65.445 -192.605 -65.115 -192.275 ;
        RECT -65.445 -193.965 -65.115 -193.635 ;
        RECT -65.445 -195.325 -65.115 -194.995 ;
        RECT -65.445 -196.685 -65.115 -196.355 ;
        RECT -65.445 -198.045 -65.115 -197.715 ;
        RECT -65.445 -199.405 -65.115 -199.075 ;
        RECT -65.445 -200.765 -65.115 -200.435 ;
        RECT -65.445 -202.125 -65.115 -201.795 ;
        RECT -65.445 -203.485 -65.115 -203.155 ;
        RECT -65.445 -204.845 -65.115 -204.515 ;
        RECT -65.445 -206.555 -65.115 -206.225 ;
        RECT -65.445 -207.565 -65.115 -207.235 ;
        RECT -65.445 -208.925 -65.115 -208.595 ;
        RECT -65.445 -211.645 -65.115 -211.315 ;
        RECT -65.445 -214.365 -65.115 -214.035 ;
        RECT -65.445 -215.725 -65.115 -215.395 ;
        RECT -65.445 -217.085 -65.115 -216.755 ;
        RECT -65.445 -218.445 -65.115 -218.115 ;
        RECT -65.445 -224.09 -65.115 -222.96 ;
        RECT -65.44 -224.205 -65.12 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -64.085 132.52 -63.755 133.65 ;
        RECT -64.085 128.355 -63.755 128.685 ;
        RECT -64.085 126.995 -63.755 127.325 ;
        RECT -64.085 125.635 -63.755 125.965 ;
        RECT -64.085 124.275 -63.755 124.605 ;
        RECT -64.085 122.915 -63.755 123.245 ;
        RECT -64.085 121.555 -63.755 121.885 ;
        RECT -64.085 120.195 -63.755 120.525 ;
        RECT -64.085 118.835 -63.755 119.165 ;
        RECT -64.085 117.475 -63.755 117.805 ;
        RECT -64.085 116.115 -63.755 116.445 ;
        RECT -64.085 114.755 -63.755 115.085 ;
        RECT -64.085 113.395 -63.755 113.725 ;
        RECT -64.085 112.035 -63.755 112.365 ;
        RECT -64.085 110.675 -63.755 111.005 ;
        RECT -64.085 109.315 -63.755 109.645 ;
        RECT -64.085 107.955 -63.755 108.285 ;
        RECT -64.085 106.595 -63.755 106.925 ;
        RECT -64.085 105.235 -63.755 105.565 ;
        RECT -64.085 103.875 -63.755 104.205 ;
        RECT -64.085 102.515 -63.755 102.845 ;
        RECT -64.085 101.155 -63.755 101.485 ;
        RECT -64.085 99.795 -63.755 100.125 ;
        RECT -64.085 98.435 -63.755 98.765 ;
        RECT -64.085 97.075 -63.755 97.405 ;
        RECT -64.085 95.715 -63.755 96.045 ;
        RECT -64.085 94.355 -63.755 94.685 ;
        RECT -64.085 92.995 -63.755 93.325 ;
        RECT -64.085 91.635 -63.755 91.965 ;
        RECT -64.085 90.275 -63.755 90.605 ;
        RECT -64.085 88.915 -63.755 89.245 ;
        RECT -64.085 87.555 -63.755 87.885 ;
        RECT -64.085 86.195 -63.755 86.525 ;
        RECT -64.085 84.835 -63.755 85.165 ;
        RECT -64.085 83.475 -63.755 83.805 ;
        RECT -64.085 82.115 -63.755 82.445 ;
        RECT -64.085 80.755 -63.755 81.085 ;
        RECT -64.085 79.395 -63.755 79.725 ;
        RECT -64.085 78.035 -63.755 78.365 ;
        RECT -64.085 76.675 -63.755 77.005 ;
        RECT -64.085 75.315 -63.755 75.645 ;
        RECT -64.085 73.955 -63.755 74.285 ;
        RECT -64.085 72.595 -63.755 72.925 ;
        RECT -64.085 71.235 -63.755 71.565 ;
        RECT -64.085 69.875 -63.755 70.205 ;
        RECT -64.085 68.515 -63.755 68.845 ;
        RECT -64.085 67.155 -63.755 67.485 ;
        RECT -64.085 65.795 -63.755 66.125 ;
        RECT -64.085 64.435 -63.755 64.765 ;
        RECT -64.085 63.075 -63.755 63.405 ;
        RECT -64.085 61.715 -63.755 62.045 ;
        RECT -64.085 60.355 -63.755 60.685 ;
        RECT -64.085 58.995 -63.755 59.325 ;
        RECT -64.085 57.635 -63.755 57.965 ;
        RECT -64.085 56.275 -63.755 56.605 ;
        RECT -64.085 54.915 -63.755 55.245 ;
        RECT -64.085 53.555 -63.755 53.885 ;
        RECT -64.085 52.195 -63.755 52.525 ;
        RECT -64.085 50.835 -63.755 51.165 ;
        RECT -64.085 49.475 -63.755 49.805 ;
        RECT -64.085 48.115 -63.755 48.445 ;
        RECT -64.085 46.755 -63.755 47.085 ;
        RECT -64.085 45.395 -63.755 45.725 ;
        RECT -64.085 44.035 -63.755 44.365 ;
        RECT -64.085 42.675 -63.755 43.005 ;
        RECT -64.085 41.315 -63.755 41.645 ;
        RECT -64.085 39.955 -63.755 40.285 ;
        RECT -64.085 38.595 -63.755 38.925 ;
        RECT -64.085 37.235 -63.755 37.565 ;
        RECT -64.085 35.875 -63.755 36.205 ;
        RECT -64.085 34.515 -63.755 34.845 ;
        RECT -64.085 33.155 -63.755 33.485 ;
        RECT -64.085 31.795 -63.755 32.125 ;
        RECT -64.085 30.435 -63.755 30.765 ;
        RECT -64.085 29.075 -63.755 29.405 ;
        RECT -64.085 27.715 -63.755 28.045 ;
        RECT -64.085 26.355 -63.755 26.685 ;
        RECT -64.085 24.995 -63.755 25.325 ;
        RECT -64.085 23.635 -63.755 23.965 ;
        RECT -64.085 22.275 -63.755 22.605 ;
        RECT -64.085 20.915 -63.755 21.245 ;
        RECT -64.085 19.555 -63.755 19.885 ;
        RECT -64.085 18.195 -63.755 18.525 ;
        RECT -64.085 16.835 -63.755 17.165 ;
        RECT -64.085 15.475 -63.755 15.805 ;
        RECT -64.085 14.115 -63.755 14.445 ;
        RECT -64.085 12.755 -63.755 13.085 ;
        RECT -64.085 11.395 -63.755 11.725 ;
        RECT -64.085 10.035 -63.755 10.365 ;
        RECT -64.085 8.675 -63.755 9.005 ;
        RECT -64.085 7.315 -63.755 7.645 ;
        RECT -64.085 5.955 -63.755 6.285 ;
        RECT -64.085 4.595 -63.755 4.925 ;
        RECT -64.085 3.235 -63.755 3.565 ;
        RECT -64.085 1.875 -63.755 2.205 ;
        RECT -64.085 0.515 -63.755 0.845 ;
        RECT -64.085 -0.845 -63.755 -0.515 ;
        RECT -64.085 -2.205 -63.755 -1.875 ;
        RECT -64.085 -3.565 -63.755 -3.235 ;
        RECT -64.085 -4.925 -63.755 -4.595 ;
        RECT -64.085 -6.285 -63.755 -5.955 ;
        RECT -64.085 -7.645 -63.755 -7.315 ;
        RECT -64.085 -9.005 -63.755 -8.675 ;
        RECT -64.085 -10.365 -63.755 -10.035 ;
        RECT -64.085 -11.725 -63.755 -11.395 ;
        RECT -64.085 -13.085 -63.755 -12.755 ;
        RECT -64.085 -14.445 -63.755 -14.115 ;
        RECT -64.085 -15.805 -63.755 -15.475 ;
        RECT -64.085 -17.165 -63.755 -16.835 ;
        RECT -64.085 -18.525 -63.755 -18.195 ;
        RECT -64.085 -19.885 -63.755 -19.555 ;
        RECT -64.085 -21.245 -63.755 -20.915 ;
        RECT -64.085 -22.605 -63.755 -22.275 ;
        RECT -64.085 -23.965 -63.755 -23.635 ;
        RECT -64.085 -25.325 -63.755 -24.995 ;
        RECT -64.085 -26.685 -63.755 -26.355 ;
        RECT -64.085 -28.045 -63.755 -27.715 ;
        RECT -64.085 -29.405 -63.755 -29.075 ;
        RECT -64.085 -30.765 -63.755 -30.435 ;
        RECT -64.085 -32.125 -63.755 -31.795 ;
        RECT -64.085 -33.485 -63.755 -33.155 ;
        RECT -64.085 -34.845 -63.755 -34.515 ;
        RECT -64.085 -36.205 -63.755 -35.875 ;
        RECT -64.085 -37.565 -63.755 -37.235 ;
        RECT -64.085 -38.925 -63.755 -38.595 ;
        RECT -64.085 -40.285 -63.755 -39.955 ;
        RECT -64.085 -41.645 -63.755 -41.315 ;
        RECT -64.085 -43.005 -63.755 -42.675 ;
        RECT -64.085 -44.365 -63.755 -44.035 ;
        RECT -64.085 -45.725 -63.755 -45.395 ;
        RECT -64.085 -47.085 -63.755 -46.755 ;
        RECT -64.085 -48.445 -63.755 -48.115 ;
        RECT -64.085 -49.805 -63.755 -49.475 ;
        RECT -64.085 -51.165 -63.755 -50.835 ;
        RECT -64.085 -52.525 -63.755 -52.195 ;
        RECT -64.085 -53.885 -63.755 -53.555 ;
        RECT -64.085 -55.245 -63.755 -54.915 ;
        RECT -64.085 -56.605 -63.755 -56.275 ;
        RECT -64.085 -57.965 -63.755 -57.635 ;
        RECT -64.085 -59.325 -63.755 -58.995 ;
        RECT -64.085 -60.685 -63.755 -60.355 ;
        RECT -64.085 -62.045 -63.755 -61.715 ;
        RECT -64.085 -63.405 -63.755 -63.075 ;
        RECT -64.085 -64.765 -63.755 -64.435 ;
        RECT -64.085 -66.125 -63.755 -65.795 ;
        RECT -64.085 -67.485 -63.755 -67.155 ;
        RECT -64.085 -68.845 -63.755 -68.515 ;
        RECT -64.085 -70.205 -63.755 -69.875 ;
        RECT -64.085 -71.565 -63.755 -71.235 ;
        RECT -64.085 -72.925 -63.755 -72.595 ;
        RECT -64.085 -74.285 -63.755 -73.955 ;
        RECT -64.085 -75.645 -63.755 -75.315 ;
        RECT -64.085 -77.005 -63.755 -76.675 ;
        RECT -64.085 -78.365 -63.755 -78.035 ;
        RECT -64.085 -79.725 -63.755 -79.395 ;
        RECT -64.085 -81.085 -63.755 -80.755 ;
        RECT -64.085 -82.445 -63.755 -82.115 ;
        RECT -64.085 -83.805 -63.755 -83.475 ;
        RECT -64.085 -85.165 -63.755 -84.835 ;
        RECT -64.085 -86.525 -63.755 -86.195 ;
        RECT -64.085 -87.885 -63.755 -87.555 ;
        RECT -64.085 -89.245 -63.755 -88.915 ;
        RECT -64.085 -90.605 -63.755 -90.275 ;
        RECT -64.085 -91.965 -63.755 -91.635 ;
        RECT -64.085 -93.325 -63.755 -92.995 ;
        RECT -64.085 -94.685 -63.755 -94.355 ;
        RECT -64.085 -96.045 -63.755 -95.715 ;
        RECT -64.085 -97.405 -63.755 -97.075 ;
        RECT -64.085 -98.765 -63.755 -98.435 ;
        RECT -64.085 -100.125 -63.755 -99.795 ;
        RECT -64.085 -101.485 -63.755 -101.155 ;
        RECT -64.085 -102.845 -63.755 -102.515 ;
        RECT -64.085 -104.205 -63.755 -103.875 ;
        RECT -64.085 -105.565 -63.755 -105.235 ;
        RECT -64.085 -106.925 -63.755 -106.595 ;
        RECT -64.085 -108.285 -63.755 -107.955 ;
        RECT -64.085 -109.645 -63.755 -109.315 ;
        RECT -64.085 -111.005 -63.755 -110.675 ;
        RECT -64.085 -112.365 -63.755 -112.035 ;
        RECT -64.085 -113.725 -63.755 -113.395 ;
        RECT -64.085 -115.085 -63.755 -114.755 ;
        RECT -64.085 -116.445 -63.755 -116.115 ;
        RECT -64.085 -117.805 -63.755 -117.475 ;
        RECT -64.085 -119.165 -63.755 -118.835 ;
        RECT -64.085 -120.525 -63.755 -120.195 ;
        RECT -64.085 -121.885 -63.755 -121.555 ;
        RECT -64.085 -123.245 -63.755 -122.915 ;
        RECT -64.085 -124.605 -63.755 -124.275 ;
        RECT -64.085 -125.965 -63.755 -125.635 ;
        RECT -64.085 -127.325 -63.755 -126.995 ;
        RECT -64.085 -128.685 -63.755 -128.355 ;
        RECT -64.085 -130.045 -63.755 -129.715 ;
        RECT -64.085 -131.405 -63.755 -131.075 ;
        RECT -64.085 -132.765 -63.755 -132.435 ;
        RECT -64.085 -134.125 -63.755 -133.795 ;
        RECT -64.085 -135.485 -63.755 -135.155 ;
        RECT -64.085 -136.845 -63.755 -136.515 ;
        RECT -64.085 -138.205 -63.755 -137.875 ;
        RECT -64.085 -139.565 -63.755 -139.235 ;
        RECT -64.085 -140.925 -63.755 -140.595 ;
        RECT -64.085 -142.285 -63.755 -141.955 ;
        RECT -64.085 -143.645 -63.755 -143.315 ;
        RECT -64.085 -145.005 -63.755 -144.675 ;
        RECT -64.085 -146.365 -63.755 -146.035 ;
        RECT -64.085 -147.725 -63.755 -147.395 ;
        RECT -64.085 -149.085 -63.755 -148.755 ;
        RECT -64.085 -150.445 -63.755 -150.115 ;
        RECT -64.085 -151.805 -63.755 -151.475 ;
        RECT -64.085 -153.165 -63.755 -152.835 ;
        RECT -64.085 -154.525 -63.755 -154.195 ;
        RECT -64.085 -155.885 -63.755 -155.555 ;
        RECT -64.085 -157.245 -63.755 -156.915 ;
        RECT -64.085 -158.605 -63.755 -158.275 ;
        RECT -64.085 -159.965 -63.755 -159.635 ;
        RECT -64.085 -161.325 -63.755 -160.995 ;
        RECT -64.085 -162.685 -63.755 -162.355 ;
        RECT -64.085 -164.045 -63.755 -163.715 ;
        RECT -64.085 -165.405 -63.755 -165.075 ;
        RECT -64.085 -166.765 -63.755 -166.435 ;
        RECT -64.085 -168.125 -63.755 -167.795 ;
        RECT -64.085 -169.485 -63.755 -169.155 ;
        RECT -64.085 -170.845 -63.755 -170.515 ;
        RECT -64.085 -172.205 -63.755 -171.875 ;
        RECT -64.085 -173.565 -63.755 -173.235 ;
        RECT -64.085 -174.925 -63.755 -174.595 ;
        RECT -64.085 -176.285 -63.755 -175.955 ;
        RECT -64.085 -177.645 -63.755 -177.315 ;
        RECT -64.085 -179.005 -63.755 -178.675 ;
        RECT -64.085 -180.365 -63.755 -180.035 ;
        RECT -64.085 -181.725 -63.755 -181.395 ;
        RECT -64.085 -183.085 -63.755 -182.755 ;
        RECT -64.085 -184.445 -63.755 -184.115 ;
        RECT -64.085 -185.805 -63.755 -185.475 ;
        RECT -64.085 -187.165 -63.755 -186.835 ;
        RECT -64.085 -188.525 -63.755 -188.195 ;
        RECT -64.085 -189.885 -63.755 -189.555 ;
        RECT -64.085 -191.245 -63.755 -190.915 ;
        RECT -64.085 -192.605 -63.755 -192.275 ;
        RECT -64.085 -193.965 -63.755 -193.635 ;
        RECT -64.085 -195.325 -63.755 -194.995 ;
        RECT -64.085 -196.685 -63.755 -196.355 ;
        RECT -64.085 -198.045 -63.755 -197.715 ;
        RECT -64.085 -199.405 -63.755 -199.075 ;
        RECT -64.085 -200.765 -63.755 -200.435 ;
        RECT -64.085 -202.125 -63.755 -201.795 ;
        RECT -64.085 -203.485 -63.755 -203.155 ;
        RECT -64.085 -204.845 -63.755 -204.515 ;
        RECT -64.085 -206.555 -63.755 -206.225 ;
        RECT -64.085 -207.565 -63.755 -207.235 ;
        RECT -64.085 -208.925 -63.755 -208.595 ;
        RECT -64.085 -211.645 -63.755 -211.315 ;
        RECT -64.085 -214.365 -63.755 -214.035 ;
        RECT -64.085 -215.725 -63.755 -215.395 ;
        RECT -64.085 -217.085 -63.755 -216.755 ;
        RECT -64.085 -218.445 -63.755 -218.115 ;
        RECT -64.085 -224.09 -63.755 -222.96 ;
        RECT -64.08 -224.205 -63.76 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -62.725 132.52 -62.395 133.65 ;
        RECT -62.725 128.355 -62.395 128.685 ;
        RECT -62.725 126.995 -62.395 127.325 ;
        RECT -62.725 125.635 -62.395 125.965 ;
        RECT -62.725 124.275 -62.395 124.605 ;
        RECT -62.725 122.915 -62.395 123.245 ;
        RECT -62.725 121.555 -62.395 121.885 ;
        RECT -62.725 120.195 -62.395 120.525 ;
        RECT -62.725 118.835 -62.395 119.165 ;
        RECT -62.725 117.475 -62.395 117.805 ;
        RECT -62.725 116.115 -62.395 116.445 ;
        RECT -62.725 114.755 -62.395 115.085 ;
        RECT -62.725 113.395 -62.395 113.725 ;
        RECT -62.725 112.035 -62.395 112.365 ;
        RECT -62.725 110.675 -62.395 111.005 ;
        RECT -62.725 109.315 -62.395 109.645 ;
        RECT -62.725 107.955 -62.395 108.285 ;
        RECT -62.725 106.595 -62.395 106.925 ;
        RECT -62.725 105.235 -62.395 105.565 ;
        RECT -62.725 103.875 -62.395 104.205 ;
        RECT -62.725 102.515 -62.395 102.845 ;
        RECT -62.725 101.155 -62.395 101.485 ;
        RECT -62.725 99.795 -62.395 100.125 ;
        RECT -62.725 98.435 -62.395 98.765 ;
        RECT -62.725 97.075 -62.395 97.405 ;
        RECT -62.725 95.715 -62.395 96.045 ;
        RECT -62.725 94.355 -62.395 94.685 ;
        RECT -62.725 92.995 -62.395 93.325 ;
        RECT -62.725 91.635 -62.395 91.965 ;
        RECT -62.725 90.275 -62.395 90.605 ;
        RECT -62.725 88.915 -62.395 89.245 ;
        RECT -62.725 87.555 -62.395 87.885 ;
        RECT -62.725 86.195 -62.395 86.525 ;
        RECT -62.725 84.835 -62.395 85.165 ;
        RECT -62.725 83.475 -62.395 83.805 ;
        RECT -62.725 82.115 -62.395 82.445 ;
        RECT -62.725 80.755 -62.395 81.085 ;
        RECT -62.725 79.395 -62.395 79.725 ;
        RECT -62.725 78.035 -62.395 78.365 ;
        RECT -62.725 76.675 -62.395 77.005 ;
        RECT -62.725 75.315 -62.395 75.645 ;
        RECT -62.725 73.955 -62.395 74.285 ;
        RECT -62.725 72.595 -62.395 72.925 ;
        RECT -62.725 71.235 -62.395 71.565 ;
        RECT -62.725 69.875 -62.395 70.205 ;
        RECT -62.725 68.515 -62.395 68.845 ;
        RECT -62.725 67.155 -62.395 67.485 ;
        RECT -62.725 65.795 -62.395 66.125 ;
        RECT -62.725 64.435 -62.395 64.765 ;
        RECT -62.725 63.075 -62.395 63.405 ;
        RECT -62.725 61.715 -62.395 62.045 ;
        RECT -62.725 60.355 -62.395 60.685 ;
        RECT -62.725 58.995 -62.395 59.325 ;
        RECT -62.725 57.635 -62.395 57.965 ;
        RECT -62.725 56.275 -62.395 56.605 ;
        RECT -62.725 54.915 -62.395 55.245 ;
        RECT -62.725 53.555 -62.395 53.885 ;
        RECT -62.725 52.195 -62.395 52.525 ;
        RECT -62.725 50.835 -62.395 51.165 ;
        RECT -62.725 49.475 -62.395 49.805 ;
        RECT -62.725 48.115 -62.395 48.445 ;
        RECT -62.725 46.755 -62.395 47.085 ;
        RECT -62.725 45.395 -62.395 45.725 ;
        RECT -62.725 44.035 -62.395 44.365 ;
        RECT -62.725 42.675 -62.395 43.005 ;
        RECT -62.725 41.315 -62.395 41.645 ;
        RECT -62.725 39.955 -62.395 40.285 ;
        RECT -62.725 38.595 -62.395 38.925 ;
        RECT -62.725 37.235 -62.395 37.565 ;
        RECT -62.725 35.875 -62.395 36.205 ;
        RECT -62.725 34.515 -62.395 34.845 ;
        RECT -62.725 33.155 -62.395 33.485 ;
        RECT -62.725 31.795 -62.395 32.125 ;
        RECT -62.725 30.435 -62.395 30.765 ;
        RECT -62.725 29.075 -62.395 29.405 ;
        RECT -62.725 27.715 -62.395 28.045 ;
        RECT -62.725 26.355 -62.395 26.685 ;
        RECT -62.725 24.995 -62.395 25.325 ;
        RECT -62.725 23.635 -62.395 23.965 ;
        RECT -62.725 22.275 -62.395 22.605 ;
        RECT -62.725 20.915 -62.395 21.245 ;
        RECT -62.725 19.555 -62.395 19.885 ;
        RECT -62.725 18.195 -62.395 18.525 ;
        RECT -62.725 16.835 -62.395 17.165 ;
        RECT -62.725 15.475 -62.395 15.805 ;
        RECT -62.725 14.115 -62.395 14.445 ;
        RECT -62.725 12.755 -62.395 13.085 ;
        RECT -62.725 11.395 -62.395 11.725 ;
        RECT -62.725 10.035 -62.395 10.365 ;
        RECT -62.725 8.675 -62.395 9.005 ;
        RECT -62.725 7.315 -62.395 7.645 ;
        RECT -62.725 5.955 -62.395 6.285 ;
        RECT -62.725 4.595 -62.395 4.925 ;
        RECT -62.725 3.235 -62.395 3.565 ;
        RECT -62.725 1.875 -62.395 2.205 ;
        RECT -62.725 0.515 -62.395 0.845 ;
        RECT -62.725 -0.845 -62.395 -0.515 ;
        RECT -62.725 -2.205 -62.395 -1.875 ;
        RECT -62.725 -3.565 -62.395 -3.235 ;
        RECT -62.725 -4.925 -62.395 -4.595 ;
        RECT -62.725 -6.285 -62.395 -5.955 ;
        RECT -62.725 -7.645 -62.395 -7.315 ;
        RECT -62.725 -9.005 -62.395 -8.675 ;
        RECT -62.725 -10.365 -62.395 -10.035 ;
        RECT -62.725 -11.725 -62.395 -11.395 ;
        RECT -62.725 -13.085 -62.395 -12.755 ;
        RECT -62.725 -14.445 -62.395 -14.115 ;
        RECT -62.725 -15.805 -62.395 -15.475 ;
        RECT -62.725 -17.165 -62.395 -16.835 ;
        RECT -62.725 -18.525 -62.395 -18.195 ;
        RECT -62.725 -19.885 -62.395 -19.555 ;
        RECT -62.725 -21.245 -62.395 -20.915 ;
        RECT -62.725 -22.605 -62.395 -22.275 ;
        RECT -62.725 -23.965 -62.395 -23.635 ;
        RECT -62.725 -25.325 -62.395 -24.995 ;
        RECT -62.725 -26.685 -62.395 -26.355 ;
        RECT -62.725 -28.045 -62.395 -27.715 ;
        RECT -62.725 -29.405 -62.395 -29.075 ;
        RECT -62.725 -30.765 -62.395 -30.435 ;
        RECT -62.725 -32.125 -62.395 -31.795 ;
        RECT -62.725 -33.485 -62.395 -33.155 ;
        RECT -62.725 -34.845 -62.395 -34.515 ;
        RECT -62.725 -36.205 -62.395 -35.875 ;
        RECT -62.725 -37.565 -62.395 -37.235 ;
        RECT -62.725 -38.925 -62.395 -38.595 ;
        RECT -62.725 -40.285 -62.395 -39.955 ;
        RECT -62.725 -41.645 -62.395 -41.315 ;
        RECT -62.725 -43.005 -62.395 -42.675 ;
        RECT -62.725 -44.365 -62.395 -44.035 ;
        RECT -62.725 -45.725 -62.395 -45.395 ;
        RECT -62.725 -47.085 -62.395 -46.755 ;
        RECT -62.725 -48.445 -62.395 -48.115 ;
        RECT -62.725 -49.805 -62.395 -49.475 ;
        RECT -62.725 -51.165 -62.395 -50.835 ;
        RECT -62.725 -52.525 -62.395 -52.195 ;
        RECT -62.725 -53.885 -62.395 -53.555 ;
        RECT -62.725 -55.245 -62.395 -54.915 ;
        RECT -62.725 -56.605 -62.395 -56.275 ;
        RECT -62.725 -57.965 -62.395 -57.635 ;
        RECT -62.725 -59.325 -62.395 -58.995 ;
        RECT -62.725 -60.685 -62.395 -60.355 ;
        RECT -62.725 -62.045 -62.395 -61.715 ;
        RECT -62.725 -63.405 -62.395 -63.075 ;
        RECT -62.725 -64.765 -62.395 -64.435 ;
        RECT -62.725 -66.125 -62.395 -65.795 ;
        RECT -62.725 -67.485 -62.395 -67.155 ;
        RECT -62.725 -68.845 -62.395 -68.515 ;
        RECT -62.725 -70.205 -62.395 -69.875 ;
        RECT -62.725 -71.565 -62.395 -71.235 ;
        RECT -62.725 -72.925 -62.395 -72.595 ;
        RECT -62.725 -74.285 -62.395 -73.955 ;
        RECT -62.725 -75.645 -62.395 -75.315 ;
        RECT -62.725 -77.005 -62.395 -76.675 ;
        RECT -62.725 -78.365 -62.395 -78.035 ;
        RECT -62.725 -79.725 -62.395 -79.395 ;
        RECT -62.725 -81.085 -62.395 -80.755 ;
        RECT -62.725 -82.445 -62.395 -82.115 ;
        RECT -62.725 -83.805 -62.395 -83.475 ;
        RECT -62.725 -85.165 -62.395 -84.835 ;
        RECT -62.725 -86.525 -62.395 -86.195 ;
        RECT -62.725 -87.885 -62.395 -87.555 ;
        RECT -62.725 -89.245 -62.395 -88.915 ;
        RECT -62.725 -90.605 -62.395 -90.275 ;
        RECT -62.725 -91.965 -62.395 -91.635 ;
        RECT -62.725 -93.325 -62.395 -92.995 ;
        RECT -62.725 -94.685 -62.395 -94.355 ;
        RECT -62.725 -96.045 -62.395 -95.715 ;
        RECT -62.725 -97.405 -62.395 -97.075 ;
        RECT -62.725 -98.765 -62.395 -98.435 ;
        RECT -62.725 -100.125 -62.395 -99.795 ;
        RECT -62.725 -101.485 -62.395 -101.155 ;
        RECT -62.725 -102.845 -62.395 -102.515 ;
        RECT -62.725 -104.205 -62.395 -103.875 ;
        RECT -62.725 -105.565 -62.395 -105.235 ;
        RECT -62.725 -106.925 -62.395 -106.595 ;
        RECT -62.725 -108.285 -62.395 -107.955 ;
        RECT -62.725 -109.645 -62.395 -109.315 ;
        RECT -62.725 -111.005 -62.395 -110.675 ;
        RECT -62.725 -112.365 -62.395 -112.035 ;
        RECT -62.725 -113.725 -62.395 -113.395 ;
        RECT -62.725 -115.085 -62.395 -114.755 ;
        RECT -62.725 -116.445 -62.395 -116.115 ;
        RECT -62.725 -117.805 -62.395 -117.475 ;
        RECT -62.725 -119.165 -62.395 -118.835 ;
        RECT -62.725 -120.525 -62.395 -120.195 ;
        RECT -62.725 -121.885 -62.395 -121.555 ;
        RECT -62.725 -123.245 -62.395 -122.915 ;
        RECT -62.725 -124.605 -62.395 -124.275 ;
        RECT -62.725 -125.965 -62.395 -125.635 ;
        RECT -62.725 -127.325 -62.395 -126.995 ;
        RECT -62.725 -128.685 -62.395 -128.355 ;
        RECT -62.725 -130.045 -62.395 -129.715 ;
        RECT -62.725 -131.405 -62.395 -131.075 ;
        RECT -62.725 -132.765 -62.395 -132.435 ;
        RECT -62.725 -134.125 -62.395 -133.795 ;
        RECT -62.725 -135.485 -62.395 -135.155 ;
        RECT -62.725 -136.845 -62.395 -136.515 ;
        RECT -62.725 -138.205 -62.395 -137.875 ;
        RECT -62.725 -139.565 -62.395 -139.235 ;
        RECT -62.725 -140.925 -62.395 -140.595 ;
        RECT -62.725 -142.285 -62.395 -141.955 ;
        RECT -62.725 -143.645 -62.395 -143.315 ;
        RECT -62.725 -145.005 -62.395 -144.675 ;
        RECT -62.725 -146.365 -62.395 -146.035 ;
        RECT -62.725 -147.725 -62.395 -147.395 ;
        RECT -62.725 -149.085 -62.395 -148.755 ;
        RECT -62.725 -150.445 -62.395 -150.115 ;
        RECT -62.725 -151.805 -62.395 -151.475 ;
        RECT -62.725 -153.165 -62.395 -152.835 ;
        RECT -62.725 -154.525 -62.395 -154.195 ;
        RECT -62.725 -155.885 -62.395 -155.555 ;
        RECT -62.725 -157.245 -62.395 -156.915 ;
        RECT -62.725 -158.605 -62.395 -158.275 ;
        RECT -62.725 -159.965 -62.395 -159.635 ;
        RECT -62.725 -161.325 -62.395 -160.995 ;
        RECT -62.725 -162.685 -62.395 -162.355 ;
        RECT -62.725 -164.045 -62.395 -163.715 ;
        RECT -62.725 -165.405 -62.395 -165.075 ;
        RECT -62.725 -166.765 -62.395 -166.435 ;
        RECT -62.725 -168.125 -62.395 -167.795 ;
        RECT -62.725 -169.485 -62.395 -169.155 ;
        RECT -62.725 -170.845 -62.395 -170.515 ;
        RECT -62.725 -172.205 -62.395 -171.875 ;
        RECT -62.725 -173.565 -62.395 -173.235 ;
        RECT -62.725 -174.925 -62.395 -174.595 ;
        RECT -62.725 -176.285 -62.395 -175.955 ;
        RECT -62.725 -177.645 -62.395 -177.315 ;
        RECT -62.725 -179.005 -62.395 -178.675 ;
        RECT -62.725 -180.365 -62.395 -180.035 ;
        RECT -62.725 -181.725 -62.395 -181.395 ;
        RECT -62.725 -183.085 -62.395 -182.755 ;
        RECT -62.725 -184.445 -62.395 -184.115 ;
        RECT -62.725 -185.805 -62.395 -185.475 ;
        RECT -62.725 -187.165 -62.395 -186.835 ;
        RECT -62.725 -188.525 -62.395 -188.195 ;
        RECT -62.725 -189.885 -62.395 -189.555 ;
        RECT -62.725 -191.245 -62.395 -190.915 ;
        RECT -62.725 -192.605 -62.395 -192.275 ;
        RECT -62.725 -193.965 -62.395 -193.635 ;
        RECT -62.725 -195.325 -62.395 -194.995 ;
        RECT -62.725 -196.685 -62.395 -196.355 ;
        RECT -62.725 -198.045 -62.395 -197.715 ;
        RECT -62.725 -199.405 -62.395 -199.075 ;
        RECT -62.725 -200.765 -62.395 -200.435 ;
        RECT -62.725 -202.125 -62.395 -201.795 ;
        RECT -62.725 -203.485 -62.395 -203.155 ;
        RECT -62.725 -204.845 -62.395 -204.515 ;
        RECT -62.725 -206.555 -62.395 -206.225 ;
        RECT -62.725 -207.565 -62.395 -207.235 ;
        RECT -62.725 -208.925 -62.395 -208.595 ;
        RECT -62.725 -210.285 -62.395 -209.955 ;
        RECT -62.725 -211.645 -62.395 -211.315 ;
        RECT -62.725 -214.365 -62.395 -214.035 ;
        RECT -62.725 -215.725 -62.395 -215.395 ;
        RECT -62.725 -217.085 -62.395 -216.755 ;
        RECT -62.725 -218.445 -62.395 -218.115 ;
        RECT -62.725 -224.09 -62.395 -222.96 ;
        RECT -62.72 -224.205 -62.4 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -61.365 -96.045 -61.035 -95.715 ;
        RECT -61.365 -97.405 -61.035 -97.075 ;
        RECT -61.365 -98.765 -61.035 -98.435 ;
        RECT -61.365 -100.125 -61.035 -99.795 ;
        RECT -61.365 -101.485 -61.035 -101.155 ;
        RECT -61.365 -102.845 -61.035 -102.515 ;
        RECT -61.365 -104.205 -61.035 -103.875 ;
        RECT -61.365 -105.565 -61.035 -105.235 ;
        RECT -61.365 -106.925 -61.035 -106.595 ;
        RECT -61.365 -108.285 -61.035 -107.955 ;
        RECT -61.365 -109.645 -61.035 -109.315 ;
        RECT -61.365 -111.005 -61.035 -110.675 ;
        RECT -61.365 -112.365 -61.035 -112.035 ;
        RECT -61.365 -113.725 -61.035 -113.395 ;
        RECT -61.365 -115.085 -61.035 -114.755 ;
        RECT -61.365 -116.445 -61.035 -116.115 ;
        RECT -61.365 -117.805 -61.035 -117.475 ;
        RECT -61.365 -119.165 -61.035 -118.835 ;
        RECT -61.365 -120.525 -61.035 -120.195 ;
        RECT -61.365 -121.885 -61.035 -121.555 ;
        RECT -61.365 -123.245 -61.035 -122.915 ;
        RECT -61.365 -124.605 -61.035 -124.275 ;
        RECT -61.365 -125.965 -61.035 -125.635 ;
        RECT -61.365 -127.325 -61.035 -126.995 ;
        RECT -61.365 -128.685 -61.035 -128.355 ;
        RECT -61.365 -130.045 -61.035 -129.715 ;
        RECT -61.365 -131.405 -61.035 -131.075 ;
        RECT -61.365 -132.765 -61.035 -132.435 ;
        RECT -61.365 -134.125 -61.035 -133.795 ;
        RECT -61.365 -135.485 -61.035 -135.155 ;
        RECT -61.365 -136.845 -61.035 -136.515 ;
        RECT -61.365 -138.205 -61.035 -137.875 ;
        RECT -61.365 -139.565 -61.035 -139.235 ;
        RECT -61.365 -140.925 -61.035 -140.595 ;
        RECT -61.365 -142.285 -61.035 -141.955 ;
        RECT -61.365 -143.645 -61.035 -143.315 ;
        RECT -61.365 -145.005 -61.035 -144.675 ;
        RECT -61.365 -146.365 -61.035 -146.035 ;
        RECT -61.365 -147.725 -61.035 -147.395 ;
        RECT -61.365 -149.085 -61.035 -148.755 ;
        RECT -61.365 -150.445 -61.035 -150.115 ;
        RECT -61.365 -151.805 -61.035 -151.475 ;
        RECT -61.365 -153.165 -61.035 -152.835 ;
        RECT -61.365 -154.525 -61.035 -154.195 ;
        RECT -61.365 -155.885 -61.035 -155.555 ;
        RECT -61.365 -157.245 -61.035 -156.915 ;
        RECT -61.365 -158.605 -61.035 -158.275 ;
        RECT -61.365 -159.965 -61.035 -159.635 ;
        RECT -61.365 -161.325 -61.035 -160.995 ;
        RECT -61.365 -162.685 -61.035 -162.355 ;
        RECT -61.365 -164.045 -61.035 -163.715 ;
        RECT -61.365 -165.405 -61.035 -165.075 ;
        RECT -61.365 -166.765 -61.035 -166.435 ;
        RECT -61.365 -168.125 -61.035 -167.795 ;
        RECT -61.365 -169.485 -61.035 -169.155 ;
        RECT -61.365 -170.845 -61.035 -170.515 ;
        RECT -61.365 -172.205 -61.035 -171.875 ;
        RECT -61.365 -173.565 -61.035 -173.235 ;
        RECT -61.365 -174.925 -61.035 -174.595 ;
        RECT -61.365 -176.285 -61.035 -175.955 ;
        RECT -61.365 -177.645 -61.035 -177.315 ;
        RECT -61.365 -179.005 -61.035 -178.675 ;
        RECT -61.365 -180.365 -61.035 -180.035 ;
        RECT -61.365 -181.725 -61.035 -181.395 ;
        RECT -61.365 -183.085 -61.035 -182.755 ;
        RECT -61.365 -184.445 -61.035 -184.115 ;
        RECT -61.365 -185.805 -61.035 -185.475 ;
        RECT -61.365 -187.165 -61.035 -186.835 ;
        RECT -61.365 -188.525 -61.035 -188.195 ;
        RECT -61.365 -189.885 -61.035 -189.555 ;
        RECT -61.365 -191.245 -61.035 -190.915 ;
        RECT -61.365 -192.605 -61.035 -192.275 ;
        RECT -61.365 -193.965 -61.035 -193.635 ;
        RECT -61.365 -195.325 -61.035 -194.995 ;
        RECT -61.365 -196.685 -61.035 -196.355 ;
        RECT -61.365 -198.045 -61.035 -197.715 ;
        RECT -61.365 -199.405 -61.035 -199.075 ;
        RECT -61.365 -200.765 -61.035 -200.435 ;
        RECT -61.365 -202.125 -61.035 -201.795 ;
        RECT -61.365 -203.485 -61.035 -203.155 ;
        RECT -61.365 -204.845 -61.035 -204.515 ;
        RECT -61.365 -206.555 -61.035 -206.225 ;
        RECT -61.365 -207.565 -61.035 -207.235 ;
        RECT -61.365 -208.925 -61.035 -208.595 ;
        RECT -61.365 -210.285 -61.035 -209.955 ;
        RECT -61.365 -211.645 -61.035 -211.315 ;
        RECT -61.365 -214.365 -61.035 -214.035 ;
        RECT -61.365 -215.725 -61.035 -215.395 ;
        RECT -61.365 -217.085 -61.035 -216.755 ;
        RECT -61.365 -218.445 -61.035 -218.115 ;
        RECT -61.365 -224.09 -61.035 -222.96 ;
        RECT -61.36 -224.205 -61.04 133.765 ;
        RECT -61.365 132.52 -61.035 133.65 ;
        RECT -61.365 128.355 -61.035 128.685 ;
        RECT -61.365 126.995 -61.035 127.325 ;
        RECT -61.365 125.635 -61.035 125.965 ;
        RECT -61.365 124.275 -61.035 124.605 ;
        RECT -61.365 122.915 -61.035 123.245 ;
        RECT -61.365 121.555 -61.035 121.885 ;
        RECT -61.365 120.195 -61.035 120.525 ;
        RECT -61.365 118.835 -61.035 119.165 ;
        RECT -61.365 117.475 -61.035 117.805 ;
        RECT -61.365 116.115 -61.035 116.445 ;
        RECT -61.365 114.755 -61.035 115.085 ;
        RECT -61.365 113.395 -61.035 113.725 ;
        RECT -61.365 112.035 -61.035 112.365 ;
        RECT -61.365 110.675 -61.035 111.005 ;
        RECT -61.365 109.315 -61.035 109.645 ;
        RECT -61.365 107.955 -61.035 108.285 ;
        RECT -61.365 106.595 -61.035 106.925 ;
        RECT -61.365 105.235 -61.035 105.565 ;
        RECT -61.365 103.875 -61.035 104.205 ;
        RECT -61.365 102.515 -61.035 102.845 ;
        RECT -61.365 101.155 -61.035 101.485 ;
        RECT -61.365 99.795 -61.035 100.125 ;
        RECT -61.365 98.435 -61.035 98.765 ;
        RECT -61.365 97.075 -61.035 97.405 ;
        RECT -61.365 95.715 -61.035 96.045 ;
        RECT -61.365 94.355 -61.035 94.685 ;
        RECT -61.365 92.995 -61.035 93.325 ;
        RECT -61.365 91.635 -61.035 91.965 ;
        RECT -61.365 90.275 -61.035 90.605 ;
        RECT -61.365 88.915 -61.035 89.245 ;
        RECT -61.365 87.555 -61.035 87.885 ;
        RECT -61.365 86.195 -61.035 86.525 ;
        RECT -61.365 84.835 -61.035 85.165 ;
        RECT -61.365 83.475 -61.035 83.805 ;
        RECT -61.365 82.115 -61.035 82.445 ;
        RECT -61.365 80.755 -61.035 81.085 ;
        RECT -61.365 79.395 -61.035 79.725 ;
        RECT -61.365 78.035 -61.035 78.365 ;
        RECT -61.365 76.675 -61.035 77.005 ;
        RECT -61.365 75.315 -61.035 75.645 ;
        RECT -61.365 73.955 -61.035 74.285 ;
        RECT -61.365 72.595 -61.035 72.925 ;
        RECT -61.365 71.235 -61.035 71.565 ;
        RECT -61.365 69.875 -61.035 70.205 ;
        RECT -61.365 68.515 -61.035 68.845 ;
        RECT -61.365 67.155 -61.035 67.485 ;
        RECT -61.365 65.795 -61.035 66.125 ;
        RECT -61.365 64.435 -61.035 64.765 ;
        RECT -61.365 63.075 -61.035 63.405 ;
        RECT -61.365 61.715 -61.035 62.045 ;
        RECT -61.365 60.355 -61.035 60.685 ;
        RECT -61.365 58.995 -61.035 59.325 ;
        RECT -61.365 57.635 -61.035 57.965 ;
        RECT -61.365 56.275 -61.035 56.605 ;
        RECT -61.365 54.915 -61.035 55.245 ;
        RECT -61.365 53.555 -61.035 53.885 ;
        RECT -61.365 52.195 -61.035 52.525 ;
        RECT -61.365 50.835 -61.035 51.165 ;
        RECT -61.365 49.475 -61.035 49.805 ;
        RECT -61.365 48.115 -61.035 48.445 ;
        RECT -61.365 46.755 -61.035 47.085 ;
        RECT -61.365 45.395 -61.035 45.725 ;
        RECT -61.365 44.035 -61.035 44.365 ;
        RECT -61.365 42.675 -61.035 43.005 ;
        RECT -61.365 41.315 -61.035 41.645 ;
        RECT -61.365 39.955 -61.035 40.285 ;
        RECT -61.365 38.595 -61.035 38.925 ;
        RECT -61.365 37.235 -61.035 37.565 ;
        RECT -61.365 35.875 -61.035 36.205 ;
        RECT -61.365 34.515 -61.035 34.845 ;
        RECT -61.365 33.155 -61.035 33.485 ;
        RECT -61.365 31.795 -61.035 32.125 ;
        RECT -61.365 30.435 -61.035 30.765 ;
        RECT -61.365 29.075 -61.035 29.405 ;
        RECT -61.365 27.715 -61.035 28.045 ;
        RECT -61.365 26.355 -61.035 26.685 ;
        RECT -61.365 24.995 -61.035 25.325 ;
        RECT -61.365 23.635 -61.035 23.965 ;
        RECT -61.365 22.275 -61.035 22.605 ;
        RECT -61.365 20.915 -61.035 21.245 ;
        RECT -61.365 19.555 -61.035 19.885 ;
        RECT -61.365 18.195 -61.035 18.525 ;
        RECT -61.365 16.835 -61.035 17.165 ;
        RECT -61.365 15.475 -61.035 15.805 ;
        RECT -61.365 14.115 -61.035 14.445 ;
        RECT -61.365 12.755 -61.035 13.085 ;
        RECT -61.365 11.395 -61.035 11.725 ;
        RECT -61.365 10.035 -61.035 10.365 ;
        RECT -61.365 8.675 -61.035 9.005 ;
        RECT -61.365 7.315 -61.035 7.645 ;
        RECT -61.365 5.955 -61.035 6.285 ;
        RECT -61.365 4.595 -61.035 4.925 ;
        RECT -61.365 3.235 -61.035 3.565 ;
        RECT -61.365 1.875 -61.035 2.205 ;
        RECT -61.365 0.515 -61.035 0.845 ;
        RECT -61.365 -0.845 -61.035 -0.515 ;
        RECT -61.365 -2.205 -61.035 -1.875 ;
        RECT -61.365 -3.565 -61.035 -3.235 ;
        RECT -61.365 -4.925 -61.035 -4.595 ;
        RECT -61.365 -6.285 -61.035 -5.955 ;
        RECT -61.365 -7.645 -61.035 -7.315 ;
        RECT -61.365 -9.005 -61.035 -8.675 ;
        RECT -61.365 -10.365 -61.035 -10.035 ;
        RECT -61.365 -11.725 -61.035 -11.395 ;
        RECT -61.365 -13.085 -61.035 -12.755 ;
        RECT -61.365 -14.445 -61.035 -14.115 ;
        RECT -61.365 -15.805 -61.035 -15.475 ;
        RECT -61.365 -17.165 -61.035 -16.835 ;
        RECT -61.365 -18.525 -61.035 -18.195 ;
        RECT -61.365 -19.885 -61.035 -19.555 ;
        RECT -61.365 -21.245 -61.035 -20.915 ;
        RECT -61.365 -22.605 -61.035 -22.275 ;
        RECT -61.365 -23.965 -61.035 -23.635 ;
        RECT -61.365 -25.325 -61.035 -24.995 ;
        RECT -61.365 -26.685 -61.035 -26.355 ;
        RECT -61.365 -28.045 -61.035 -27.715 ;
        RECT -61.365 -29.405 -61.035 -29.075 ;
        RECT -61.365 -30.765 -61.035 -30.435 ;
        RECT -61.365 -32.125 -61.035 -31.795 ;
        RECT -61.365 -33.485 -61.035 -33.155 ;
        RECT -61.365 -34.845 -61.035 -34.515 ;
        RECT -61.365 -36.205 -61.035 -35.875 ;
        RECT -61.365 -37.565 -61.035 -37.235 ;
        RECT -61.365 -38.925 -61.035 -38.595 ;
        RECT -61.365 -40.285 -61.035 -39.955 ;
        RECT -61.365 -41.645 -61.035 -41.315 ;
        RECT -61.365 -43.005 -61.035 -42.675 ;
        RECT -61.365 -44.365 -61.035 -44.035 ;
        RECT -61.365 -45.725 -61.035 -45.395 ;
        RECT -61.365 -47.085 -61.035 -46.755 ;
        RECT -61.365 -48.445 -61.035 -48.115 ;
        RECT -61.365 -49.805 -61.035 -49.475 ;
        RECT -61.365 -51.165 -61.035 -50.835 ;
        RECT -61.365 -52.525 -61.035 -52.195 ;
        RECT -61.365 -53.885 -61.035 -53.555 ;
        RECT -61.365 -55.245 -61.035 -54.915 ;
        RECT -61.365 -56.605 -61.035 -56.275 ;
        RECT -61.365 -57.965 -61.035 -57.635 ;
        RECT -61.365 -59.325 -61.035 -58.995 ;
        RECT -61.365 -60.685 -61.035 -60.355 ;
        RECT -61.365 -62.045 -61.035 -61.715 ;
        RECT -61.365 -63.405 -61.035 -63.075 ;
        RECT -61.365 -64.765 -61.035 -64.435 ;
        RECT -61.365 -66.125 -61.035 -65.795 ;
        RECT -61.365 -67.485 -61.035 -67.155 ;
        RECT -61.365 -68.845 -61.035 -68.515 ;
        RECT -61.365 -70.205 -61.035 -69.875 ;
        RECT -61.365 -71.565 -61.035 -71.235 ;
        RECT -61.365 -72.925 -61.035 -72.595 ;
        RECT -61.365 -74.285 -61.035 -73.955 ;
        RECT -61.365 -75.645 -61.035 -75.315 ;
        RECT -61.365 -77.005 -61.035 -76.675 ;
        RECT -61.365 -78.365 -61.035 -78.035 ;
        RECT -61.365 -79.725 -61.035 -79.395 ;
        RECT -61.365 -81.085 -61.035 -80.755 ;
        RECT -61.365 -82.445 -61.035 -82.115 ;
        RECT -61.365 -83.805 -61.035 -83.475 ;
        RECT -61.365 -85.165 -61.035 -84.835 ;
        RECT -61.365 -86.525 -61.035 -86.195 ;
        RECT -61.365 -87.885 -61.035 -87.555 ;
        RECT -61.365 -89.245 -61.035 -88.915 ;
        RECT -61.365 -90.605 -61.035 -90.275 ;
        RECT -61.365 -91.965 -61.035 -91.635 ;
        RECT -61.365 -93.325 -61.035 -92.995 ;
        RECT -61.365 -94.685 -61.035 -94.355 ;
    END
    PORT
      LAYER met3 ;
        RECT -70.885 132.52 -70.555 133.65 ;
        RECT -70.885 128.355 -70.555 128.685 ;
        RECT -70.885 126.995 -70.555 127.325 ;
        RECT -70.885 125.635 -70.555 125.965 ;
        RECT -70.885 124.275 -70.555 124.605 ;
        RECT -70.885 122.915 -70.555 123.245 ;
        RECT -70.885 121.555 -70.555 121.885 ;
        RECT -70.885 120.195 -70.555 120.525 ;
        RECT -70.885 118.835 -70.555 119.165 ;
        RECT -70.885 117.475 -70.555 117.805 ;
        RECT -70.885 116.115 -70.555 116.445 ;
        RECT -70.885 114.755 -70.555 115.085 ;
        RECT -70.885 113.395 -70.555 113.725 ;
        RECT -70.885 112.035 -70.555 112.365 ;
        RECT -70.885 110.675 -70.555 111.005 ;
        RECT -70.885 109.315 -70.555 109.645 ;
        RECT -70.885 107.955 -70.555 108.285 ;
        RECT -70.885 106.595 -70.555 106.925 ;
        RECT -70.885 105.235 -70.555 105.565 ;
        RECT -70.885 103.875 -70.555 104.205 ;
        RECT -70.885 102.515 -70.555 102.845 ;
        RECT -70.885 101.155 -70.555 101.485 ;
        RECT -70.885 99.795 -70.555 100.125 ;
        RECT -70.885 98.435 -70.555 98.765 ;
        RECT -70.885 97.075 -70.555 97.405 ;
        RECT -70.885 95.715 -70.555 96.045 ;
        RECT -70.885 94.355 -70.555 94.685 ;
        RECT -70.885 92.995 -70.555 93.325 ;
        RECT -70.885 91.635 -70.555 91.965 ;
        RECT -70.885 90.275 -70.555 90.605 ;
        RECT -70.885 88.915 -70.555 89.245 ;
        RECT -70.885 87.555 -70.555 87.885 ;
        RECT -70.885 86.195 -70.555 86.525 ;
        RECT -70.885 84.835 -70.555 85.165 ;
        RECT -70.885 83.475 -70.555 83.805 ;
        RECT -70.885 82.115 -70.555 82.445 ;
        RECT -70.885 80.755 -70.555 81.085 ;
        RECT -70.885 79.395 -70.555 79.725 ;
        RECT -70.885 78.035 -70.555 78.365 ;
        RECT -70.885 76.675 -70.555 77.005 ;
        RECT -70.885 75.315 -70.555 75.645 ;
        RECT -70.885 73.955 -70.555 74.285 ;
        RECT -70.885 72.595 -70.555 72.925 ;
        RECT -70.885 71.235 -70.555 71.565 ;
        RECT -70.885 69.875 -70.555 70.205 ;
        RECT -70.885 68.515 -70.555 68.845 ;
        RECT -70.885 67.155 -70.555 67.485 ;
        RECT -70.885 65.795 -70.555 66.125 ;
        RECT -70.885 64.435 -70.555 64.765 ;
        RECT -70.885 63.075 -70.555 63.405 ;
        RECT -70.885 61.715 -70.555 62.045 ;
        RECT -70.885 60.355 -70.555 60.685 ;
        RECT -70.885 58.995 -70.555 59.325 ;
        RECT -70.885 57.635 -70.555 57.965 ;
        RECT -70.885 56.275 -70.555 56.605 ;
        RECT -70.885 54.915 -70.555 55.245 ;
        RECT -70.885 53.555 -70.555 53.885 ;
        RECT -70.885 52.195 -70.555 52.525 ;
        RECT -70.885 50.835 -70.555 51.165 ;
        RECT -70.885 49.475 -70.555 49.805 ;
        RECT -70.885 48.115 -70.555 48.445 ;
        RECT -70.885 46.755 -70.555 47.085 ;
        RECT -70.885 45.395 -70.555 45.725 ;
        RECT -70.885 44.035 -70.555 44.365 ;
        RECT -70.885 42.675 -70.555 43.005 ;
        RECT -70.885 41.315 -70.555 41.645 ;
        RECT -70.885 39.955 -70.555 40.285 ;
        RECT -70.885 38.595 -70.555 38.925 ;
        RECT -70.885 37.235 -70.555 37.565 ;
        RECT -70.885 35.875 -70.555 36.205 ;
        RECT -70.885 34.515 -70.555 34.845 ;
        RECT -70.885 33.155 -70.555 33.485 ;
        RECT -70.885 31.795 -70.555 32.125 ;
        RECT -70.885 30.435 -70.555 30.765 ;
        RECT -70.885 29.075 -70.555 29.405 ;
        RECT -70.885 27.715 -70.555 28.045 ;
        RECT -70.885 26.355 -70.555 26.685 ;
        RECT -70.885 24.995 -70.555 25.325 ;
        RECT -70.885 23.635 -70.555 23.965 ;
        RECT -70.885 22.275 -70.555 22.605 ;
        RECT -70.885 20.915 -70.555 21.245 ;
        RECT -70.885 19.555 -70.555 19.885 ;
        RECT -70.885 18.195 -70.555 18.525 ;
        RECT -70.885 16.835 -70.555 17.165 ;
        RECT -70.885 15.475 -70.555 15.805 ;
        RECT -70.885 14.115 -70.555 14.445 ;
        RECT -70.885 12.755 -70.555 13.085 ;
        RECT -70.885 11.395 -70.555 11.725 ;
        RECT -70.885 10.035 -70.555 10.365 ;
        RECT -70.885 8.675 -70.555 9.005 ;
        RECT -70.885 7.315 -70.555 7.645 ;
        RECT -70.885 5.955 -70.555 6.285 ;
        RECT -70.885 4.595 -70.555 4.925 ;
        RECT -70.885 3.235 -70.555 3.565 ;
        RECT -70.885 1.875 -70.555 2.205 ;
        RECT -70.885 0.515 -70.555 0.845 ;
        RECT -70.885 -0.845 -70.555 -0.515 ;
        RECT -70.885 -2.205 -70.555 -1.875 ;
        RECT -70.885 -3.565 -70.555 -3.235 ;
        RECT -70.885 -4.925 -70.555 -4.595 ;
        RECT -70.885 -6.285 -70.555 -5.955 ;
        RECT -70.885 -7.645 -70.555 -7.315 ;
        RECT -70.885 -9.005 -70.555 -8.675 ;
        RECT -70.885 -10.365 -70.555 -10.035 ;
        RECT -70.885 -11.725 -70.555 -11.395 ;
        RECT -70.885 -13.085 -70.555 -12.755 ;
        RECT -70.885 -14.445 -70.555 -14.115 ;
        RECT -70.885 -15.805 -70.555 -15.475 ;
        RECT -70.885 -17.165 -70.555 -16.835 ;
        RECT -70.885 -18.525 -70.555 -18.195 ;
        RECT -70.885 -19.885 -70.555 -19.555 ;
        RECT -70.885 -21.245 -70.555 -20.915 ;
        RECT -70.885 -22.605 -70.555 -22.275 ;
        RECT -70.885 -23.965 -70.555 -23.635 ;
        RECT -70.885 -25.325 -70.555 -24.995 ;
        RECT -70.885 -26.685 -70.555 -26.355 ;
        RECT -70.885 -28.045 -70.555 -27.715 ;
        RECT -70.885 -29.405 -70.555 -29.075 ;
        RECT -70.885 -30.765 -70.555 -30.435 ;
        RECT -70.885 -32.125 -70.555 -31.795 ;
        RECT -70.885 -33.485 -70.555 -33.155 ;
        RECT -70.885 -34.845 -70.555 -34.515 ;
        RECT -70.885 -36.205 -70.555 -35.875 ;
        RECT -70.885 -37.565 -70.555 -37.235 ;
        RECT -70.885 -38.925 -70.555 -38.595 ;
        RECT -70.885 -40.285 -70.555 -39.955 ;
        RECT -70.885 -41.645 -70.555 -41.315 ;
        RECT -70.885 -43.005 -70.555 -42.675 ;
        RECT -70.885 -44.365 -70.555 -44.035 ;
        RECT -70.885 -45.725 -70.555 -45.395 ;
        RECT -70.885 -47.085 -70.555 -46.755 ;
        RECT -70.885 -48.445 -70.555 -48.115 ;
        RECT -70.885 -49.805 -70.555 -49.475 ;
        RECT -70.885 -51.165 -70.555 -50.835 ;
        RECT -70.885 -52.525 -70.555 -52.195 ;
        RECT -70.885 -53.885 -70.555 -53.555 ;
        RECT -70.885 -55.245 -70.555 -54.915 ;
        RECT -70.885 -56.605 -70.555 -56.275 ;
        RECT -70.885 -57.965 -70.555 -57.635 ;
        RECT -70.885 -59.325 -70.555 -58.995 ;
        RECT -70.885 -60.685 -70.555 -60.355 ;
        RECT -70.885 -62.045 -70.555 -61.715 ;
        RECT -70.885 -63.405 -70.555 -63.075 ;
        RECT -70.885 -64.765 -70.555 -64.435 ;
        RECT -70.885 -66.125 -70.555 -65.795 ;
        RECT -70.885 -67.485 -70.555 -67.155 ;
        RECT -70.885 -68.845 -70.555 -68.515 ;
        RECT -70.885 -70.205 -70.555 -69.875 ;
        RECT -70.885 -71.565 -70.555 -71.235 ;
        RECT -70.885 -72.925 -70.555 -72.595 ;
        RECT -70.885 -74.285 -70.555 -73.955 ;
        RECT -70.885 -75.645 -70.555 -75.315 ;
        RECT -70.885 -77.005 -70.555 -76.675 ;
        RECT -70.885 -78.365 -70.555 -78.035 ;
        RECT -70.885 -79.725 -70.555 -79.395 ;
        RECT -70.885 -81.085 -70.555 -80.755 ;
        RECT -70.885 -82.445 -70.555 -82.115 ;
        RECT -70.885 -83.805 -70.555 -83.475 ;
        RECT -70.885 -85.165 -70.555 -84.835 ;
        RECT -70.885 -86.525 -70.555 -86.195 ;
        RECT -70.885 -87.885 -70.555 -87.555 ;
        RECT -70.885 -89.245 -70.555 -88.915 ;
        RECT -70.885 -90.605 -70.555 -90.275 ;
        RECT -70.885 -91.965 -70.555 -91.635 ;
        RECT -70.885 -93.325 -70.555 -92.995 ;
        RECT -70.885 -94.685 -70.555 -94.355 ;
        RECT -70.885 -96.045 -70.555 -95.715 ;
        RECT -70.885 -97.405 -70.555 -97.075 ;
        RECT -70.885 -98.765 -70.555 -98.435 ;
        RECT -70.885 -100.125 -70.555 -99.795 ;
        RECT -70.885 -101.485 -70.555 -101.155 ;
        RECT -70.885 -102.845 -70.555 -102.515 ;
        RECT -70.885 -104.205 -70.555 -103.875 ;
        RECT -70.885 -105.565 -70.555 -105.235 ;
        RECT -70.885 -106.925 -70.555 -106.595 ;
        RECT -70.885 -108.285 -70.555 -107.955 ;
        RECT -70.885 -109.645 -70.555 -109.315 ;
        RECT -70.885 -111.005 -70.555 -110.675 ;
        RECT -70.885 -112.365 -70.555 -112.035 ;
        RECT -70.885 -113.725 -70.555 -113.395 ;
        RECT -70.885 -115.085 -70.555 -114.755 ;
        RECT -70.885 -116.445 -70.555 -116.115 ;
        RECT -70.885 -117.805 -70.555 -117.475 ;
        RECT -70.885 -119.165 -70.555 -118.835 ;
        RECT -70.885 -120.525 -70.555 -120.195 ;
        RECT -70.885 -121.885 -70.555 -121.555 ;
        RECT -70.885 -123.245 -70.555 -122.915 ;
        RECT -70.885 -124.605 -70.555 -124.275 ;
        RECT -70.885 -125.965 -70.555 -125.635 ;
        RECT -70.885 -127.325 -70.555 -126.995 ;
        RECT -70.885 -128.685 -70.555 -128.355 ;
        RECT -70.885 -130.045 -70.555 -129.715 ;
        RECT -70.885 -131.405 -70.555 -131.075 ;
        RECT -70.885 -132.765 -70.555 -132.435 ;
        RECT -70.885 -134.125 -70.555 -133.795 ;
        RECT -70.885 -135.485 -70.555 -135.155 ;
        RECT -70.885 -136.845 -70.555 -136.515 ;
        RECT -70.885 -138.205 -70.555 -137.875 ;
        RECT -70.885 -139.565 -70.555 -139.235 ;
        RECT -70.885 -140.925 -70.555 -140.595 ;
        RECT -70.885 -142.285 -70.555 -141.955 ;
        RECT -70.885 -143.645 -70.555 -143.315 ;
        RECT -70.885 -145.005 -70.555 -144.675 ;
        RECT -70.885 -146.365 -70.555 -146.035 ;
        RECT -70.885 -147.725 -70.555 -147.395 ;
        RECT -70.885 -149.085 -70.555 -148.755 ;
        RECT -70.885 -150.445 -70.555 -150.115 ;
        RECT -70.885 -151.805 -70.555 -151.475 ;
        RECT -70.885 -153.165 -70.555 -152.835 ;
        RECT -70.885 -154.525 -70.555 -154.195 ;
        RECT -70.885 -155.885 -70.555 -155.555 ;
        RECT -70.885 -157.245 -70.555 -156.915 ;
        RECT -70.885 -158.605 -70.555 -158.275 ;
        RECT -70.885 -159.965 -70.555 -159.635 ;
        RECT -70.885 -161.325 -70.555 -160.995 ;
        RECT -70.885 -162.685 -70.555 -162.355 ;
        RECT -70.885 -164.045 -70.555 -163.715 ;
        RECT -70.885 -165.405 -70.555 -165.075 ;
        RECT -70.885 -166.765 -70.555 -166.435 ;
        RECT -70.885 -168.125 -70.555 -167.795 ;
        RECT -70.885 -169.485 -70.555 -169.155 ;
        RECT -70.885 -170.845 -70.555 -170.515 ;
        RECT -70.885 -172.205 -70.555 -171.875 ;
        RECT -70.885 -173.565 -70.555 -173.235 ;
        RECT -70.885 -174.925 -70.555 -174.595 ;
        RECT -70.885 -176.285 -70.555 -175.955 ;
        RECT -70.885 -177.645 -70.555 -177.315 ;
        RECT -70.885 -179.005 -70.555 -178.675 ;
        RECT -70.885 -180.365 -70.555 -180.035 ;
        RECT -70.885 -181.725 -70.555 -181.395 ;
        RECT -70.885 -183.085 -70.555 -182.755 ;
        RECT -70.885 -184.445 -70.555 -184.115 ;
        RECT -70.885 -185.805 -70.555 -185.475 ;
        RECT -70.885 -187.165 -70.555 -186.835 ;
        RECT -70.885 -188.525 -70.555 -188.195 ;
        RECT -70.885 -189.885 -70.555 -189.555 ;
        RECT -70.885 -191.245 -70.555 -190.915 ;
        RECT -70.885 -192.605 -70.555 -192.275 ;
        RECT -70.885 -193.965 -70.555 -193.635 ;
        RECT -70.885 -195.325 -70.555 -194.995 ;
        RECT -70.885 -196.685 -70.555 -196.355 ;
        RECT -70.885 -198.045 -70.555 -197.715 ;
        RECT -70.885 -199.405 -70.555 -199.075 ;
        RECT -70.885 -200.765 -70.555 -200.435 ;
        RECT -70.885 -202.125 -70.555 -201.795 ;
        RECT -70.885 -203.485 -70.555 -203.155 ;
        RECT -70.885 -204.845 -70.555 -204.515 ;
        RECT -70.885 -206.205 -70.555 -205.875 ;
        RECT -70.885 -207.565 -70.555 -207.235 ;
        RECT -70.885 -208.925 -70.555 -208.595 ;
        RECT -70.885 -210.285 -70.555 -209.955 ;
        RECT -70.885 -211.645 -70.555 -211.315 ;
        RECT -70.885 -213.005 -70.555 -212.675 ;
        RECT -70.885 -214.365 -70.555 -214.035 ;
        RECT -70.885 -215.725 -70.555 -215.395 ;
        RECT -70.885 -217.085 -70.555 -216.755 ;
        RECT -70.885 -218.445 -70.555 -218.115 ;
        RECT -70.885 -224.09 -70.555 -222.96 ;
        RECT -70.88 -224.205 -70.56 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -69.525 132.52 -69.195 133.65 ;
        RECT -69.525 128.355 -69.195 128.685 ;
        RECT -69.525 126.995 -69.195 127.325 ;
        RECT -69.525 125.635 -69.195 125.965 ;
        RECT -69.525 124.275 -69.195 124.605 ;
        RECT -69.525 122.915 -69.195 123.245 ;
        RECT -69.525 121.555 -69.195 121.885 ;
        RECT -69.525 120.195 -69.195 120.525 ;
        RECT -69.525 118.835 -69.195 119.165 ;
        RECT -69.525 117.475 -69.195 117.805 ;
        RECT -69.525 116.115 -69.195 116.445 ;
        RECT -69.525 114.755 -69.195 115.085 ;
        RECT -69.525 113.395 -69.195 113.725 ;
        RECT -69.525 112.035 -69.195 112.365 ;
        RECT -69.525 110.675 -69.195 111.005 ;
        RECT -69.525 109.315 -69.195 109.645 ;
        RECT -69.525 107.955 -69.195 108.285 ;
        RECT -69.525 106.595 -69.195 106.925 ;
        RECT -69.525 105.235 -69.195 105.565 ;
        RECT -69.525 103.875 -69.195 104.205 ;
        RECT -69.525 102.515 -69.195 102.845 ;
        RECT -69.525 101.155 -69.195 101.485 ;
        RECT -69.525 99.795 -69.195 100.125 ;
        RECT -69.525 98.435 -69.195 98.765 ;
        RECT -69.525 97.075 -69.195 97.405 ;
        RECT -69.525 95.715 -69.195 96.045 ;
        RECT -69.525 94.355 -69.195 94.685 ;
        RECT -69.525 92.995 -69.195 93.325 ;
        RECT -69.525 91.635 -69.195 91.965 ;
        RECT -69.525 90.275 -69.195 90.605 ;
        RECT -69.525 88.915 -69.195 89.245 ;
        RECT -69.525 87.555 -69.195 87.885 ;
        RECT -69.525 86.195 -69.195 86.525 ;
        RECT -69.525 84.835 -69.195 85.165 ;
        RECT -69.525 83.475 -69.195 83.805 ;
        RECT -69.525 82.115 -69.195 82.445 ;
        RECT -69.525 80.755 -69.195 81.085 ;
        RECT -69.525 79.395 -69.195 79.725 ;
        RECT -69.525 78.035 -69.195 78.365 ;
        RECT -69.525 76.675 -69.195 77.005 ;
        RECT -69.525 75.315 -69.195 75.645 ;
        RECT -69.525 73.955 -69.195 74.285 ;
        RECT -69.525 72.595 -69.195 72.925 ;
        RECT -69.525 71.235 -69.195 71.565 ;
        RECT -69.525 69.875 -69.195 70.205 ;
        RECT -69.525 68.515 -69.195 68.845 ;
        RECT -69.525 67.155 -69.195 67.485 ;
        RECT -69.525 65.795 -69.195 66.125 ;
        RECT -69.525 64.435 -69.195 64.765 ;
        RECT -69.525 63.075 -69.195 63.405 ;
        RECT -69.525 61.715 -69.195 62.045 ;
        RECT -69.525 60.355 -69.195 60.685 ;
        RECT -69.525 58.995 -69.195 59.325 ;
        RECT -69.525 57.635 -69.195 57.965 ;
        RECT -69.525 56.275 -69.195 56.605 ;
        RECT -69.525 54.915 -69.195 55.245 ;
        RECT -69.525 53.555 -69.195 53.885 ;
        RECT -69.525 52.195 -69.195 52.525 ;
        RECT -69.525 50.835 -69.195 51.165 ;
        RECT -69.525 49.475 -69.195 49.805 ;
        RECT -69.525 48.115 -69.195 48.445 ;
        RECT -69.525 46.755 -69.195 47.085 ;
        RECT -69.525 45.395 -69.195 45.725 ;
        RECT -69.525 44.035 -69.195 44.365 ;
        RECT -69.525 42.675 -69.195 43.005 ;
        RECT -69.525 41.315 -69.195 41.645 ;
        RECT -69.525 39.955 -69.195 40.285 ;
        RECT -69.525 38.595 -69.195 38.925 ;
        RECT -69.525 37.235 -69.195 37.565 ;
        RECT -69.525 35.875 -69.195 36.205 ;
        RECT -69.525 34.515 -69.195 34.845 ;
        RECT -69.525 33.155 -69.195 33.485 ;
        RECT -69.525 31.795 -69.195 32.125 ;
        RECT -69.525 30.435 -69.195 30.765 ;
        RECT -69.525 29.075 -69.195 29.405 ;
        RECT -69.525 27.715 -69.195 28.045 ;
        RECT -69.525 26.355 -69.195 26.685 ;
        RECT -69.525 24.995 -69.195 25.325 ;
        RECT -69.525 23.635 -69.195 23.965 ;
        RECT -69.525 22.275 -69.195 22.605 ;
        RECT -69.525 20.915 -69.195 21.245 ;
        RECT -69.525 19.555 -69.195 19.885 ;
        RECT -69.525 18.195 -69.195 18.525 ;
        RECT -69.525 16.835 -69.195 17.165 ;
        RECT -69.525 15.475 -69.195 15.805 ;
        RECT -69.525 14.115 -69.195 14.445 ;
        RECT -69.525 12.755 -69.195 13.085 ;
        RECT -69.525 11.395 -69.195 11.725 ;
        RECT -69.525 10.035 -69.195 10.365 ;
        RECT -69.525 8.675 -69.195 9.005 ;
        RECT -69.525 7.315 -69.195 7.645 ;
        RECT -69.525 5.955 -69.195 6.285 ;
        RECT -69.525 4.595 -69.195 4.925 ;
        RECT -69.525 3.235 -69.195 3.565 ;
        RECT -69.525 1.875 -69.195 2.205 ;
        RECT -69.525 0.515 -69.195 0.845 ;
        RECT -69.525 -0.845 -69.195 -0.515 ;
        RECT -69.525 -2.205 -69.195 -1.875 ;
        RECT -69.525 -3.565 -69.195 -3.235 ;
        RECT -69.525 -4.925 -69.195 -4.595 ;
        RECT -69.525 -6.285 -69.195 -5.955 ;
        RECT -69.525 -7.645 -69.195 -7.315 ;
        RECT -69.525 -9.005 -69.195 -8.675 ;
        RECT -69.525 -10.365 -69.195 -10.035 ;
        RECT -69.525 -11.725 -69.195 -11.395 ;
        RECT -69.525 -13.085 -69.195 -12.755 ;
        RECT -69.525 -14.445 -69.195 -14.115 ;
        RECT -69.525 -15.805 -69.195 -15.475 ;
        RECT -69.525 -17.165 -69.195 -16.835 ;
        RECT -69.525 -18.525 -69.195 -18.195 ;
        RECT -69.525 -19.885 -69.195 -19.555 ;
        RECT -69.525 -21.245 -69.195 -20.915 ;
        RECT -69.525 -22.605 -69.195 -22.275 ;
        RECT -69.525 -23.965 -69.195 -23.635 ;
        RECT -69.525 -25.325 -69.195 -24.995 ;
        RECT -69.525 -26.685 -69.195 -26.355 ;
        RECT -69.525 -28.045 -69.195 -27.715 ;
        RECT -69.525 -29.405 -69.195 -29.075 ;
        RECT -69.525 -30.765 -69.195 -30.435 ;
        RECT -69.525 -32.125 -69.195 -31.795 ;
        RECT -69.525 -33.485 -69.195 -33.155 ;
        RECT -69.525 -34.845 -69.195 -34.515 ;
        RECT -69.525 -36.205 -69.195 -35.875 ;
        RECT -69.525 -37.565 -69.195 -37.235 ;
        RECT -69.525 -38.925 -69.195 -38.595 ;
        RECT -69.525 -40.285 -69.195 -39.955 ;
        RECT -69.525 -41.645 -69.195 -41.315 ;
        RECT -69.525 -43.005 -69.195 -42.675 ;
        RECT -69.525 -44.365 -69.195 -44.035 ;
        RECT -69.525 -45.725 -69.195 -45.395 ;
        RECT -69.525 -47.085 -69.195 -46.755 ;
        RECT -69.525 -48.445 -69.195 -48.115 ;
        RECT -69.525 -49.805 -69.195 -49.475 ;
        RECT -69.525 -51.165 -69.195 -50.835 ;
        RECT -69.525 -52.525 -69.195 -52.195 ;
        RECT -69.525 -53.885 -69.195 -53.555 ;
        RECT -69.525 -55.245 -69.195 -54.915 ;
        RECT -69.525 -56.605 -69.195 -56.275 ;
        RECT -69.525 -57.965 -69.195 -57.635 ;
        RECT -69.525 -59.325 -69.195 -58.995 ;
        RECT -69.525 -60.685 -69.195 -60.355 ;
        RECT -69.525 -62.045 -69.195 -61.715 ;
        RECT -69.525 -63.405 -69.195 -63.075 ;
        RECT -69.525 -64.765 -69.195 -64.435 ;
        RECT -69.525 -66.125 -69.195 -65.795 ;
        RECT -69.525 -67.485 -69.195 -67.155 ;
        RECT -69.525 -68.845 -69.195 -68.515 ;
        RECT -69.525 -70.205 -69.195 -69.875 ;
        RECT -69.525 -71.565 -69.195 -71.235 ;
        RECT -69.525 -72.925 -69.195 -72.595 ;
        RECT -69.525 -74.285 -69.195 -73.955 ;
        RECT -69.525 -75.645 -69.195 -75.315 ;
        RECT -69.525 -77.005 -69.195 -76.675 ;
        RECT -69.525 -78.365 -69.195 -78.035 ;
        RECT -69.525 -79.725 -69.195 -79.395 ;
        RECT -69.525 -81.085 -69.195 -80.755 ;
        RECT -69.525 -82.445 -69.195 -82.115 ;
        RECT -69.525 -83.805 -69.195 -83.475 ;
        RECT -69.525 -85.165 -69.195 -84.835 ;
        RECT -69.525 -86.525 -69.195 -86.195 ;
        RECT -69.525 -87.885 -69.195 -87.555 ;
        RECT -69.525 -89.245 -69.195 -88.915 ;
        RECT -69.525 -90.605 -69.195 -90.275 ;
        RECT -69.525 -91.965 -69.195 -91.635 ;
        RECT -69.525 -93.325 -69.195 -92.995 ;
        RECT -69.525 -94.685 -69.195 -94.355 ;
        RECT -69.525 -96.045 -69.195 -95.715 ;
        RECT -69.525 -97.405 -69.195 -97.075 ;
        RECT -69.525 -98.765 -69.195 -98.435 ;
        RECT -69.525 -100.125 -69.195 -99.795 ;
        RECT -69.525 -101.485 -69.195 -101.155 ;
        RECT -69.525 -102.845 -69.195 -102.515 ;
        RECT -69.525 -104.205 -69.195 -103.875 ;
        RECT -69.525 -105.565 -69.195 -105.235 ;
        RECT -69.525 -106.925 -69.195 -106.595 ;
        RECT -69.525 -108.285 -69.195 -107.955 ;
        RECT -69.525 -109.645 -69.195 -109.315 ;
        RECT -69.525 -111.005 -69.195 -110.675 ;
        RECT -69.525 -112.365 -69.195 -112.035 ;
        RECT -69.525 -113.725 -69.195 -113.395 ;
        RECT -69.525 -115.085 -69.195 -114.755 ;
        RECT -69.525 -116.445 -69.195 -116.115 ;
        RECT -69.525 -117.805 -69.195 -117.475 ;
        RECT -69.525 -119.165 -69.195 -118.835 ;
        RECT -69.525 -120.525 -69.195 -120.195 ;
        RECT -69.525 -121.885 -69.195 -121.555 ;
        RECT -69.525 -123.245 -69.195 -122.915 ;
        RECT -69.525 -124.605 -69.195 -124.275 ;
        RECT -69.525 -125.965 -69.195 -125.635 ;
        RECT -69.525 -127.325 -69.195 -126.995 ;
        RECT -69.525 -128.685 -69.195 -128.355 ;
        RECT -69.525 -130.045 -69.195 -129.715 ;
        RECT -69.525 -131.405 -69.195 -131.075 ;
        RECT -69.525 -132.765 -69.195 -132.435 ;
        RECT -69.525 -134.125 -69.195 -133.795 ;
        RECT -69.525 -135.485 -69.195 -135.155 ;
        RECT -69.525 -136.845 -69.195 -136.515 ;
        RECT -69.525 -138.205 -69.195 -137.875 ;
        RECT -69.525 -139.565 -69.195 -139.235 ;
        RECT -69.525 -140.925 -69.195 -140.595 ;
        RECT -69.525 -142.285 -69.195 -141.955 ;
        RECT -69.525 -143.645 -69.195 -143.315 ;
        RECT -69.525 -145.005 -69.195 -144.675 ;
        RECT -69.525 -146.365 -69.195 -146.035 ;
        RECT -69.525 -147.725 -69.195 -147.395 ;
        RECT -69.525 -149.085 -69.195 -148.755 ;
        RECT -69.525 -150.445 -69.195 -150.115 ;
        RECT -69.525 -151.805 -69.195 -151.475 ;
        RECT -69.525 -153.165 -69.195 -152.835 ;
        RECT -69.525 -154.525 -69.195 -154.195 ;
        RECT -69.525 -155.885 -69.195 -155.555 ;
        RECT -69.525 -157.245 -69.195 -156.915 ;
        RECT -69.525 -158.605 -69.195 -158.275 ;
        RECT -69.525 -159.965 -69.195 -159.635 ;
        RECT -69.525 -161.325 -69.195 -160.995 ;
        RECT -69.525 -162.685 -69.195 -162.355 ;
        RECT -69.525 -164.045 -69.195 -163.715 ;
        RECT -69.525 -165.405 -69.195 -165.075 ;
        RECT -69.525 -166.765 -69.195 -166.435 ;
        RECT -69.525 -168.125 -69.195 -167.795 ;
        RECT -69.525 -169.485 -69.195 -169.155 ;
        RECT -69.525 -170.845 -69.195 -170.515 ;
        RECT -69.525 -172.205 -69.195 -171.875 ;
        RECT -69.525 -173.565 -69.195 -173.235 ;
        RECT -69.525 -174.925 -69.195 -174.595 ;
        RECT -69.525 -176.285 -69.195 -175.955 ;
        RECT -69.525 -177.645 -69.195 -177.315 ;
        RECT -69.525 -179.005 -69.195 -178.675 ;
        RECT -69.525 -180.365 -69.195 -180.035 ;
        RECT -69.525 -181.725 -69.195 -181.395 ;
        RECT -69.525 -183.085 -69.195 -182.755 ;
        RECT -69.525 -184.445 -69.195 -184.115 ;
        RECT -69.525 -185.805 -69.195 -185.475 ;
        RECT -69.525 -187.165 -69.195 -186.835 ;
        RECT -69.525 -188.525 -69.195 -188.195 ;
        RECT -69.525 -189.885 -69.195 -189.555 ;
        RECT -69.525 -191.245 -69.195 -190.915 ;
        RECT -69.525 -192.605 -69.195 -192.275 ;
        RECT -69.525 -193.965 -69.195 -193.635 ;
        RECT -69.525 -195.325 -69.195 -194.995 ;
        RECT -69.525 -196.685 -69.195 -196.355 ;
        RECT -69.525 -198.045 -69.195 -197.715 ;
        RECT -69.525 -199.405 -69.195 -199.075 ;
        RECT -69.525 -200.765 -69.195 -200.435 ;
        RECT -69.525 -202.125 -69.195 -201.795 ;
        RECT -69.525 -203.485 -69.195 -203.155 ;
        RECT -69.525 -204.845 -69.195 -204.515 ;
        RECT -69.525 -206.205 -69.195 -205.875 ;
        RECT -69.525 -207.565 -69.195 -207.235 ;
        RECT -69.525 -208.925 -69.195 -208.595 ;
        RECT -69.525 -210.285 -69.195 -209.955 ;
        RECT -69.525 -211.645 -69.195 -211.315 ;
        RECT -69.525 -213.005 -69.195 -212.675 ;
        RECT -69.525 -214.365 -69.195 -214.035 ;
        RECT -69.525 -215.725 -69.195 -215.395 ;
        RECT -69.525 -217.085 -69.195 -216.755 ;
        RECT -69.525 -218.445 -69.195 -218.115 ;
        RECT -69.525 -224.09 -69.195 -222.96 ;
        RECT -69.52 -224.205 -69.2 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -68.165 132.52 -67.835 133.65 ;
        RECT -68.165 128.355 -67.835 128.685 ;
        RECT -68.165 126.995 -67.835 127.325 ;
        RECT -68.165 125.635 -67.835 125.965 ;
        RECT -68.165 124.275 -67.835 124.605 ;
        RECT -68.165 122.915 -67.835 123.245 ;
        RECT -68.165 121.555 -67.835 121.885 ;
        RECT -68.165 120.195 -67.835 120.525 ;
        RECT -68.165 118.835 -67.835 119.165 ;
        RECT -68.165 117.475 -67.835 117.805 ;
        RECT -68.165 116.115 -67.835 116.445 ;
        RECT -68.165 114.755 -67.835 115.085 ;
        RECT -68.165 113.395 -67.835 113.725 ;
        RECT -68.165 112.035 -67.835 112.365 ;
        RECT -68.165 110.675 -67.835 111.005 ;
        RECT -68.165 109.315 -67.835 109.645 ;
        RECT -68.165 107.955 -67.835 108.285 ;
        RECT -68.165 106.595 -67.835 106.925 ;
        RECT -68.165 105.235 -67.835 105.565 ;
        RECT -68.165 103.875 -67.835 104.205 ;
        RECT -68.165 102.515 -67.835 102.845 ;
        RECT -68.165 101.155 -67.835 101.485 ;
        RECT -68.165 99.795 -67.835 100.125 ;
        RECT -68.165 98.435 -67.835 98.765 ;
        RECT -68.165 97.075 -67.835 97.405 ;
        RECT -68.165 95.715 -67.835 96.045 ;
        RECT -68.165 94.355 -67.835 94.685 ;
        RECT -68.165 92.995 -67.835 93.325 ;
        RECT -68.165 91.635 -67.835 91.965 ;
        RECT -68.165 90.275 -67.835 90.605 ;
        RECT -68.165 88.915 -67.835 89.245 ;
        RECT -68.165 87.555 -67.835 87.885 ;
        RECT -68.165 86.195 -67.835 86.525 ;
        RECT -68.165 84.835 -67.835 85.165 ;
        RECT -68.165 83.475 -67.835 83.805 ;
        RECT -68.165 82.115 -67.835 82.445 ;
        RECT -68.165 80.755 -67.835 81.085 ;
        RECT -68.165 79.395 -67.835 79.725 ;
        RECT -68.165 78.035 -67.835 78.365 ;
        RECT -68.165 76.675 -67.835 77.005 ;
        RECT -68.165 75.315 -67.835 75.645 ;
        RECT -68.165 73.955 -67.835 74.285 ;
        RECT -68.165 72.595 -67.835 72.925 ;
        RECT -68.165 71.235 -67.835 71.565 ;
        RECT -68.165 69.875 -67.835 70.205 ;
        RECT -68.165 68.515 -67.835 68.845 ;
        RECT -68.165 67.155 -67.835 67.485 ;
        RECT -68.165 65.795 -67.835 66.125 ;
        RECT -68.165 64.435 -67.835 64.765 ;
        RECT -68.165 63.075 -67.835 63.405 ;
        RECT -68.165 61.715 -67.835 62.045 ;
        RECT -68.165 60.355 -67.835 60.685 ;
        RECT -68.165 58.995 -67.835 59.325 ;
        RECT -68.165 57.635 -67.835 57.965 ;
        RECT -68.165 56.275 -67.835 56.605 ;
        RECT -68.165 54.915 -67.835 55.245 ;
        RECT -68.165 53.555 -67.835 53.885 ;
        RECT -68.165 52.195 -67.835 52.525 ;
        RECT -68.165 50.835 -67.835 51.165 ;
        RECT -68.165 49.475 -67.835 49.805 ;
        RECT -68.165 48.115 -67.835 48.445 ;
        RECT -68.165 46.755 -67.835 47.085 ;
        RECT -68.165 45.395 -67.835 45.725 ;
        RECT -68.165 44.035 -67.835 44.365 ;
        RECT -68.165 42.675 -67.835 43.005 ;
        RECT -68.165 41.315 -67.835 41.645 ;
        RECT -68.165 39.955 -67.835 40.285 ;
        RECT -68.165 38.595 -67.835 38.925 ;
        RECT -68.165 37.235 -67.835 37.565 ;
        RECT -68.165 35.875 -67.835 36.205 ;
        RECT -68.165 34.515 -67.835 34.845 ;
        RECT -68.165 33.155 -67.835 33.485 ;
        RECT -68.165 31.795 -67.835 32.125 ;
        RECT -68.165 30.435 -67.835 30.765 ;
        RECT -68.165 29.075 -67.835 29.405 ;
        RECT -68.165 27.715 -67.835 28.045 ;
        RECT -68.165 26.355 -67.835 26.685 ;
        RECT -68.165 24.995 -67.835 25.325 ;
        RECT -68.165 23.635 -67.835 23.965 ;
        RECT -68.165 22.275 -67.835 22.605 ;
        RECT -68.165 20.915 -67.835 21.245 ;
        RECT -68.165 19.555 -67.835 19.885 ;
        RECT -68.165 18.195 -67.835 18.525 ;
        RECT -68.165 16.835 -67.835 17.165 ;
        RECT -68.165 15.475 -67.835 15.805 ;
        RECT -68.165 14.115 -67.835 14.445 ;
        RECT -68.165 12.755 -67.835 13.085 ;
        RECT -68.165 11.395 -67.835 11.725 ;
        RECT -68.165 10.035 -67.835 10.365 ;
        RECT -68.165 8.675 -67.835 9.005 ;
        RECT -68.165 7.315 -67.835 7.645 ;
        RECT -68.165 5.955 -67.835 6.285 ;
        RECT -68.165 4.595 -67.835 4.925 ;
        RECT -68.165 3.235 -67.835 3.565 ;
        RECT -68.165 1.875 -67.835 2.205 ;
        RECT -68.165 0.515 -67.835 0.845 ;
        RECT -68.165 -0.845 -67.835 -0.515 ;
        RECT -68.165 -2.205 -67.835 -1.875 ;
        RECT -68.165 -3.565 -67.835 -3.235 ;
        RECT -68.165 -4.925 -67.835 -4.595 ;
        RECT -68.165 -6.285 -67.835 -5.955 ;
        RECT -68.165 -7.645 -67.835 -7.315 ;
        RECT -68.165 -9.005 -67.835 -8.675 ;
        RECT -68.165 -10.365 -67.835 -10.035 ;
        RECT -68.165 -11.725 -67.835 -11.395 ;
        RECT -68.165 -13.085 -67.835 -12.755 ;
        RECT -68.165 -14.445 -67.835 -14.115 ;
        RECT -68.165 -15.805 -67.835 -15.475 ;
        RECT -68.165 -17.165 -67.835 -16.835 ;
        RECT -68.165 -18.525 -67.835 -18.195 ;
        RECT -68.165 -19.885 -67.835 -19.555 ;
        RECT -68.165 -21.245 -67.835 -20.915 ;
        RECT -68.165 -22.605 -67.835 -22.275 ;
        RECT -68.165 -23.965 -67.835 -23.635 ;
        RECT -68.165 -25.325 -67.835 -24.995 ;
        RECT -68.165 -26.685 -67.835 -26.355 ;
        RECT -68.165 -28.045 -67.835 -27.715 ;
        RECT -68.165 -29.405 -67.835 -29.075 ;
        RECT -68.165 -30.765 -67.835 -30.435 ;
        RECT -68.165 -32.125 -67.835 -31.795 ;
        RECT -68.165 -33.485 -67.835 -33.155 ;
        RECT -68.165 -34.845 -67.835 -34.515 ;
        RECT -68.165 -36.205 -67.835 -35.875 ;
        RECT -68.165 -37.565 -67.835 -37.235 ;
        RECT -68.165 -38.925 -67.835 -38.595 ;
        RECT -68.165 -40.285 -67.835 -39.955 ;
        RECT -68.165 -41.645 -67.835 -41.315 ;
        RECT -68.165 -43.005 -67.835 -42.675 ;
        RECT -68.165 -44.365 -67.835 -44.035 ;
        RECT -68.165 -45.725 -67.835 -45.395 ;
        RECT -68.165 -47.085 -67.835 -46.755 ;
        RECT -68.165 -48.445 -67.835 -48.115 ;
        RECT -68.165 -49.805 -67.835 -49.475 ;
        RECT -68.165 -51.165 -67.835 -50.835 ;
        RECT -68.165 -52.525 -67.835 -52.195 ;
        RECT -68.165 -53.885 -67.835 -53.555 ;
        RECT -68.165 -55.245 -67.835 -54.915 ;
        RECT -68.165 -56.605 -67.835 -56.275 ;
        RECT -68.165 -57.965 -67.835 -57.635 ;
        RECT -68.165 -59.325 -67.835 -58.995 ;
        RECT -68.165 -60.685 -67.835 -60.355 ;
        RECT -68.165 -62.045 -67.835 -61.715 ;
        RECT -68.165 -63.405 -67.835 -63.075 ;
        RECT -68.165 -64.765 -67.835 -64.435 ;
        RECT -68.165 -66.125 -67.835 -65.795 ;
        RECT -68.165 -67.485 -67.835 -67.155 ;
        RECT -68.165 -68.845 -67.835 -68.515 ;
        RECT -68.165 -70.205 -67.835 -69.875 ;
        RECT -68.165 -71.565 -67.835 -71.235 ;
        RECT -68.165 -72.925 -67.835 -72.595 ;
        RECT -68.165 -74.285 -67.835 -73.955 ;
        RECT -68.165 -75.645 -67.835 -75.315 ;
        RECT -68.165 -77.005 -67.835 -76.675 ;
        RECT -68.165 -78.365 -67.835 -78.035 ;
        RECT -68.165 -79.725 -67.835 -79.395 ;
        RECT -68.165 -81.085 -67.835 -80.755 ;
        RECT -68.165 -82.445 -67.835 -82.115 ;
        RECT -68.165 -83.805 -67.835 -83.475 ;
        RECT -68.165 -85.165 -67.835 -84.835 ;
        RECT -68.165 -86.525 -67.835 -86.195 ;
        RECT -68.165 -87.885 -67.835 -87.555 ;
        RECT -68.165 -89.245 -67.835 -88.915 ;
        RECT -68.165 -90.605 -67.835 -90.275 ;
        RECT -68.165 -91.965 -67.835 -91.635 ;
        RECT -68.165 -93.325 -67.835 -92.995 ;
        RECT -68.165 -94.685 -67.835 -94.355 ;
        RECT -68.165 -96.045 -67.835 -95.715 ;
        RECT -68.165 -97.405 -67.835 -97.075 ;
        RECT -68.165 -98.765 -67.835 -98.435 ;
        RECT -68.165 -100.125 -67.835 -99.795 ;
        RECT -68.165 -101.485 -67.835 -101.155 ;
        RECT -68.165 -102.845 -67.835 -102.515 ;
        RECT -68.165 -104.205 -67.835 -103.875 ;
        RECT -68.165 -105.565 -67.835 -105.235 ;
        RECT -68.165 -106.925 -67.835 -106.595 ;
        RECT -68.165 -108.285 -67.835 -107.955 ;
        RECT -68.165 -109.645 -67.835 -109.315 ;
        RECT -68.165 -111.005 -67.835 -110.675 ;
        RECT -68.165 -112.365 -67.835 -112.035 ;
        RECT -68.165 -113.725 -67.835 -113.395 ;
        RECT -68.165 -115.085 -67.835 -114.755 ;
        RECT -68.165 -116.445 -67.835 -116.115 ;
        RECT -68.165 -117.805 -67.835 -117.475 ;
        RECT -68.165 -119.165 -67.835 -118.835 ;
        RECT -68.165 -120.525 -67.835 -120.195 ;
        RECT -68.165 -121.885 -67.835 -121.555 ;
        RECT -68.165 -123.245 -67.835 -122.915 ;
        RECT -68.165 -124.605 -67.835 -124.275 ;
        RECT -68.165 -125.965 -67.835 -125.635 ;
        RECT -68.165 -127.325 -67.835 -126.995 ;
        RECT -68.165 -128.685 -67.835 -128.355 ;
        RECT -68.165 -130.045 -67.835 -129.715 ;
        RECT -68.165 -131.405 -67.835 -131.075 ;
        RECT -68.165 -132.765 -67.835 -132.435 ;
        RECT -68.165 -134.125 -67.835 -133.795 ;
        RECT -68.165 -135.485 -67.835 -135.155 ;
        RECT -68.165 -136.845 -67.835 -136.515 ;
        RECT -68.165 -138.205 -67.835 -137.875 ;
        RECT -68.165 -139.565 -67.835 -139.235 ;
        RECT -68.165 -140.925 -67.835 -140.595 ;
        RECT -68.165 -142.285 -67.835 -141.955 ;
        RECT -68.165 -143.645 -67.835 -143.315 ;
        RECT -68.165 -145.005 -67.835 -144.675 ;
        RECT -68.165 -146.365 -67.835 -146.035 ;
        RECT -68.165 -147.725 -67.835 -147.395 ;
        RECT -68.165 -149.085 -67.835 -148.755 ;
        RECT -68.165 -150.445 -67.835 -150.115 ;
        RECT -68.165 -151.805 -67.835 -151.475 ;
        RECT -68.165 -153.165 -67.835 -152.835 ;
        RECT -68.165 -154.525 -67.835 -154.195 ;
        RECT -68.165 -155.885 -67.835 -155.555 ;
        RECT -68.165 -157.245 -67.835 -156.915 ;
        RECT -68.165 -158.605 -67.835 -158.275 ;
        RECT -68.165 -159.965 -67.835 -159.635 ;
        RECT -68.165 -161.325 -67.835 -160.995 ;
        RECT -68.165 -162.685 -67.835 -162.355 ;
        RECT -68.165 -164.045 -67.835 -163.715 ;
        RECT -68.165 -165.405 -67.835 -165.075 ;
        RECT -68.165 -166.765 -67.835 -166.435 ;
        RECT -68.165 -168.125 -67.835 -167.795 ;
        RECT -68.165 -169.485 -67.835 -169.155 ;
        RECT -68.165 -170.845 -67.835 -170.515 ;
        RECT -68.165 -172.205 -67.835 -171.875 ;
        RECT -68.165 -173.565 -67.835 -173.235 ;
        RECT -68.165 -174.925 -67.835 -174.595 ;
        RECT -68.165 -176.285 -67.835 -175.955 ;
        RECT -68.165 -177.645 -67.835 -177.315 ;
        RECT -68.165 -179.005 -67.835 -178.675 ;
        RECT -68.165 -180.365 -67.835 -180.035 ;
        RECT -68.165 -181.725 -67.835 -181.395 ;
        RECT -68.165 -183.085 -67.835 -182.755 ;
        RECT -68.165 -184.445 -67.835 -184.115 ;
        RECT -68.165 -185.805 -67.835 -185.475 ;
        RECT -68.165 -187.165 -67.835 -186.835 ;
        RECT -68.165 -188.525 -67.835 -188.195 ;
        RECT -68.165 -189.885 -67.835 -189.555 ;
        RECT -68.165 -191.245 -67.835 -190.915 ;
        RECT -68.165 -192.605 -67.835 -192.275 ;
        RECT -68.165 -193.965 -67.835 -193.635 ;
        RECT -68.165 -195.325 -67.835 -194.995 ;
        RECT -68.165 -196.685 -67.835 -196.355 ;
        RECT -68.165 -198.045 -67.835 -197.715 ;
        RECT -68.165 -199.405 -67.835 -199.075 ;
        RECT -68.165 -200.765 -67.835 -200.435 ;
        RECT -68.165 -202.125 -67.835 -201.795 ;
        RECT -68.165 -203.485 -67.835 -203.155 ;
        RECT -68.165 -204.845 -67.835 -204.515 ;
        RECT -68.165 -206.205 -67.835 -205.875 ;
        RECT -68.165 -207.565 -67.835 -207.235 ;
        RECT -68.165 -208.925 -67.835 -208.595 ;
        RECT -68.165 -210.285 -67.835 -209.955 ;
        RECT -68.165 -211.645 -67.835 -211.315 ;
        RECT -68.165 -213.005 -67.835 -212.675 ;
        RECT -68.165 -214.365 -67.835 -214.035 ;
        RECT -68.165 -215.725 -67.835 -215.395 ;
        RECT -68.165 -217.085 -67.835 -216.755 ;
        RECT -68.165 -218.445 -67.835 -218.115 ;
        RECT -68.165 -224.09 -67.835 -222.96 ;
        RECT -68.16 -224.205 -67.84 133.765 ;
    END
    PORT
      LAYER met3 ;
        RECT -66.805 -55.245 -66.475 -54.915 ;
        RECT -66.805 -56.605 -66.475 -56.275 ;
        RECT -66.805 -57.965 -66.475 -57.635 ;
        RECT -66.805 -59.325 -66.475 -58.995 ;
        RECT -66.805 -60.685 -66.475 -60.355 ;
        RECT -66.805 -62.045 -66.475 -61.715 ;
        RECT -66.805 -63.405 -66.475 -63.075 ;
        RECT -66.805 -64.765 -66.475 -64.435 ;
        RECT -66.805 -66.125 -66.475 -65.795 ;
        RECT -66.805 -67.485 -66.475 -67.155 ;
        RECT -66.805 -68.845 -66.475 -68.515 ;
        RECT -66.805 -70.205 -66.475 -69.875 ;
        RECT -66.805 -71.565 -66.475 -71.235 ;
        RECT -66.805 -72.925 -66.475 -72.595 ;
        RECT -66.805 -74.285 -66.475 -73.955 ;
        RECT -66.805 -75.645 -66.475 -75.315 ;
        RECT -66.805 -77.005 -66.475 -76.675 ;
        RECT -66.805 -78.365 -66.475 -78.035 ;
        RECT -66.805 -79.725 -66.475 -79.395 ;
        RECT -66.805 -81.085 -66.475 -80.755 ;
        RECT -66.805 -82.445 -66.475 -82.115 ;
        RECT -66.805 -83.805 -66.475 -83.475 ;
        RECT -66.805 -85.165 -66.475 -84.835 ;
        RECT -66.805 -86.525 -66.475 -86.195 ;
        RECT -66.805 -87.885 -66.475 -87.555 ;
        RECT -66.805 -89.245 -66.475 -88.915 ;
        RECT -66.805 -90.605 -66.475 -90.275 ;
        RECT -66.805 -91.965 -66.475 -91.635 ;
        RECT -66.805 -93.325 -66.475 -92.995 ;
        RECT -66.805 -94.685 -66.475 -94.355 ;
        RECT -66.805 -96.045 -66.475 -95.715 ;
        RECT -66.805 -97.405 -66.475 -97.075 ;
        RECT -66.805 -98.765 -66.475 -98.435 ;
        RECT -66.805 -100.125 -66.475 -99.795 ;
        RECT -66.805 -101.485 -66.475 -101.155 ;
        RECT -66.805 -102.845 -66.475 -102.515 ;
        RECT -66.805 -104.205 -66.475 -103.875 ;
        RECT -66.805 -105.565 -66.475 -105.235 ;
        RECT -66.805 -106.925 -66.475 -106.595 ;
        RECT -66.805 -108.285 -66.475 -107.955 ;
        RECT -66.805 -109.645 -66.475 -109.315 ;
        RECT -66.805 -111.005 -66.475 -110.675 ;
        RECT -66.805 -112.365 -66.475 -112.035 ;
        RECT -66.805 -113.725 -66.475 -113.395 ;
        RECT -66.805 -115.085 -66.475 -114.755 ;
        RECT -66.805 -116.445 -66.475 -116.115 ;
        RECT -66.805 -117.805 -66.475 -117.475 ;
        RECT -66.805 -119.165 -66.475 -118.835 ;
        RECT -66.805 -120.525 -66.475 -120.195 ;
        RECT -66.805 -121.885 -66.475 -121.555 ;
        RECT -66.805 -123.245 -66.475 -122.915 ;
        RECT -66.805 -124.605 -66.475 -124.275 ;
        RECT -66.805 -125.965 -66.475 -125.635 ;
        RECT -66.805 -127.325 -66.475 -126.995 ;
        RECT -66.805 -128.685 -66.475 -128.355 ;
        RECT -66.805 -130.045 -66.475 -129.715 ;
        RECT -66.805 -131.405 -66.475 -131.075 ;
        RECT -66.805 -132.765 -66.475 -132.435 ;
        RECT -66.805 -134.125 -66.475 -133.795 ;
        RECT -66.805 -135.485 -66.475 -135.155 ;
        RECT -66.805 -136.845 -66.475 -136.515 ;
        RECT -66.805 -138.205 -66.475 -137.875 ;
        RECT -66.805 -139.565 -66.475 -139.235 ;
        RECT -66.805 -140.925 -66.475 -140.595 ;
        RECT -66.805 -142.285 -66.475 -141.955 ;
        RECT -66.805 -143.645 -66.475 -143.315 ;
        RECT -66.805 -145.005 -66.475 -144.675 ;
        RECT -66.805 -146.365 -66.475 -146.035 ;
        RECT -66.805 -147.725 -66.475 -147.395 ;
        RECT -66.805 -149.085 -66.475 -148.755 ;
        RECT -66.805 -150.445 -66.475 -150.115 ;
        RECT -66.805 -151.805 -66.475 -151.475 ;
        RECT -66.805 -153.165 -66.475 -152.835 ;
        RECT -66.805 -154.525 -66.475 -154.195 ;
        RECT -66.805 -155.885 -66.475 -155.555 ;
        RECT -66.805 -157.245 -66.475 -156.915 ;
        RECT -66.805 -158.605 -66.475 -158.275 ;
        RECT -66.805 -159.965 -66.475 -159.635 ;
        RECT -66.805 -161.325 -66.475 -160.995 ;
        RECT -66.805 -162.685 -66.475 -162.355 ;
        RECT -66.805 -164.045 -66.475 -163.715 ;
        RECT -66.805 -165.405 -66.475 -165.075 ;
        RECT -66.805 -166.765 -66.475 -166.435 ;
        RECT -66.805 -168.125 -66.475 -167.795 ;
        RECT -66.805 -169.485 -66.475 -169.155 ;
        RECT -66.805 -170.845 -66.475 -170.515 ;
        RECT -66.805 -172.205 -66.475 -171.875 ;
        RECT -66.805 -173.565 -66.475 -173.235 ;
        RECT -66.805 -174.925 -66.475 -174.595 ;
        RECT -66.805 -176.285 -66.475 -175.955 ;
        RECT -66.805 -177.645 -66.475 -177.315 ;
        RECT -66.805 -179.005 -66.475 -178.675 ;
        RECT -66.805 -180.365 -66.475 -180.035 ;
        RECT -66.805 -181.725 -66.475 -181.395 ;
        RECT -66.805 -183.085 -66.475 -182.755 ;
        RECT -66.805 -184.445 -66.475 -184.115 ;
        RECT -66.805 -185.805 -66.475 -185.475 ;
        RECT -66.805 -187.165 -66.475 -186.835 ;
        RECT -66.805 -188.525 -66.475 -188.195 ;
        RECT -66.805 -189.885 -66.475 -189.555 ;
        RECT -66.805 -191.245 -66.475 -190.915 ;
        RECT -66.805 -192.605 -66.475 -192.275 ;
        RECT -66.805 -193.965 -66.475 -193.635 ;
        RECT -66.805 -195.325 -66.475 -194.995 ;
        RECT -66.805 -196.685 -66.475 -196.355 ;
        RECT -66.805 -198.045 -66.475 -197.715 ;
        RECT -66.805 -199.405 -66.475 -199.075 ;
        RECT -66.805 -200.765 -66.475 -200.435 ;
        RECT -66.805 -202.125 -66.475 -201.795 ;
        RECT -66.805 -203.485 -66.475 -203.155 ;
        RECT -66.805 -204.845 -66.475 -204.515 ;
        RECT -66.805 -206.205 -66.475 -205.875 ;
        RECT -66.805 -207.565 -66.475 -207.235 ;
        RECT -66.805 -208.925 -66.475 -208.595 ;
        RECT -66.805 -210.285 -66.475 -209.955 ;
        RECT -66.805 -211.645 -66.475 -211.315 ;
        RECT -66.805 -213.005 -66.475 -212.675 ;
        RECT -66.805 -214.365 -66.475 -214.035 ;
        RECT -66.805 -215.725 -66.475 -215.395 ;
        RECT -66.805 -217.085 -66.475 -216.755 ;
        RECT -66.805 -218.445 -66.475 -218.115 ;
        RECT -66.805 -224.09 -66.475 -222.96 ;
        RECT -66.8 -224.205 -66.48 133.765 ;
        RECT -66.805 132.52 -66.475 133.65 ;
        RECT -66.805 128.355 -66.475 128.685 ;
        RECT -66.805 126.995 -66.475 127.325 ;
        RECT -66.805 125.635 -66.475 125.965 ;
        RECT -66.805 124.275 -66.475 124.605 ;
        RECT -66.805 122.915 -66.475 123.245 ;
        RECT -66.805 121.555 -66.475 121.885 ;
        RECT -66.805 120.195 -66.475 120.525 ;
        RECT -66.805 118.835 -66.475 119.165 ;
        RECT -66.805 117.475 -66.475 117.805 ;
        RECT -66.805 116.115 -66.475 116.445 ;
        RECT -66.805 114.755 -66.475 115.085 ;
        RECT -66.805 113.395 -66.475 113.725 ;
        RECT -66.805 112.035 -66.475 112.365 ;
        RECT -66.805 110.675 -66.475 111.005 ;
        RECT -66.805 109.315 -66.475 109.645 ;
        RECT -66.805 107.955 -66.475 108.285 ;
        RECT -66.805 106.595 -66.475 106.925 ;
        RECT -66.805 105.235 -66.475 105.565 ;
        RECT -66.805 103.875 -66.475 104.205 ;
        RECT -66.805 102.515 -66.475 102.845 ;
        RECT -66.805 101.155 -66.475 101.485 ;
        RECT -66.805 99.795 -66.475 100.125 ;
        RECT -66.805 98.435 -66.475 98.765 ;
        RECT -66.805 97.075 -66.475 97.405 ;
        RECT -66.805 95.715 -66.475 96.045 ;
        RECT -66.805 94.355 -66.475 94.685 ;
        RECT -66.805 92.995 -66.475 93.325 ;
        RECT -66.805 91.635 -66.475 91.965 ;
        RECT -66.805 90.275 -66.475 90.605 ;
        RECT -66.805 88.915 -66.475 89.245 ;
        RECT -66.805 87.555 -66.475 87.885 ;
        RECT -66.805 86.195 -66.475 86.525 ;
        RECT -66.805 84.835 -66.475 85.165 ;
        RECT -66.805 83.475 -66.475 83.805 ;
        RECT -66.805 82.115 -66.475 82.445 ;
        RECT -66.805 80.755 -66.475 81.085 ;
        RECT -66.805 79.395 -66.475 79.725 ;
        RECT -66.805 78.035 -66.475 78.365 ;
        RECT -66.805 76.675 -66.475 77.005 ;
        RECT -66.805 75.315 -66.475 75.645 ;
        RECT -66.805 73.955 -66.475 74.285 ;
        RECT -66.805 72.595 -66.475 72.925 ;
        RECT -66.805 71.235 -66.475 71.565 ;
        RECT -66.805 69.875 -66.475 70.205 ;
        RECT -66.805 68.515 -66.475 68.845 ;
        RECT -66.805 67.155 -66.475 67.485 ;
        RECT -66.805 65.795 -66.475 66.125 ;
        RECT -66.805 64.435 -66.475 64.765 ;
        RECT -66.805 63.075 -66.475 63.405 ;
        RECT -66.805 61.715 -66.475 62.045 ;
        RECT -66.805 60.355 -66.475 60.685 ;
        RECT -66.805 58.995 -66.475 59.325 ;
        RECT -66.805 57.635 -66.475 57.965 ;
        RECT -66.805 56.275 -66.475 56.605 ;
        RECT -66.805 54.915 -66.475 55.245 ;
        RECT -66.805 53.555 -66.475 53.885 ;
        RECT -66.805 52.195 -66.475 52.525 ;
        RECT -66.805 50.835 -66.475 51.165 ;
        RECT -66.805 49.475 -66.475 49.805 ;
        RECT -66.805 48.115 -66.475 48.445 ;
        RECT -66.805 46.755 -66.475 47.085 ;
        RECT -66.805 45.395 -66.475 45.725 ;
        RECT -66.805 44.035 -66.475 44.365 ;
        RECT -66.805 42.675 -66.475 43.005 ;
        RECT -66.805 41.315 -66.475 41.645 ;
        RECT -66.805 39.955 -66.475 40.285 ;
        RECT -66.805 38.595 -66.475 38.925 ;
        RECT -66.805 37.235 -66.475 37.565 ;
        RECT -66.805 35.875 -66.475 36.205 ;
        RECT -66.805 34.515 -66.475 34.845 ;
        RECT -66.805 33.155 -66.475 33.485 ;
        RECT -66.805 31.795 -66.475 32.125 ;
        RECT -66.805 30.435 -66.475 30.765 ;
        RECT -66.805 29.075 -66.475 29.405 ;
        RECT -66.805 27.715 -66.475 28.045 ;
        RECT -66.805 26.355 -66.475 26.685 ;
        RECT -66.805 24.995 -66.475 25.325 ;
        RECT -66.805 23.635 -66.475 23.965 ;
        RECT -66.805 22.275 -66.475 22.605 ;
        RECT -66.805 20.915 -66.475 21.245 ;
        RECT -66.805 19.555 -66.475 19.885 ;
        RECT -66.805 18.195 -66.475 18.525 ;
        RECT -66.805 16.835 -66.475 17.165 ;
        RECT -66.805 15.475 -66.475 15.805 ;
        RECT -66.805 14.115 -66.475 14.445 ;
        RECT -66.805 12.755 -66.475 13.085 ;
        RECT -66.805 11.395 -66.475 11.725 ;
        RECT -66.805 10.035 -66.475 10.365 ;
        RECT -66.805 8.675 -66.475 9.005 ;
        RECT -66.805 7.315 -66.475 7.645 ;
        RECT -66.805 5.955 -66.475 6.285 ;
        RECT -66.805 4.595 -66.475 4.925 ;
        RECT -66.805 3.235 -66.475 3.565 ;
        RECT -66.805 1.875 -66.475 2.205 ;
        RECT -66.805 0.515 -66.475 0.845 ;
        RECT -66.805 -0.845 -66.475 -0.515 ;
        RECT -66.805 -2.205 -66.475 -1.875 ;
        RECT -66.805 -3.565 -66.475 -3.235 ;
        RECT -66.805 -4.925 -66.475 -4.595 ;
        RECT -66.805 -6.285 -66.475 -5.955 ;
        RECT -66.805 -7.645 -66.475 -7.315 ;
        RECT -66.805 -9.005 -66.475 -8.675 ;
        RECT -66.805 -10.365 -66.475 -10.035 ;
        RECT -66.805 -11.725 -66.475 -11.395 ;
        RECT -66.805 -13.085 -66.475 -12.755 ;
        RECT -66.805 -14.445 -66.475 -14.115 ;
        RECT -66.805 -15.805 -66.475 -15.475 ;
        RECT -66.805 -17.165 -66.475 -16.835 ;
        RECT -66.805 -18.525 -66.475 -18.195 ;
        RECT -66.805 -19.885 -66.475 -19.555 ;
        RECT -66.805 -21.245 -66.475 -20.915 ;
        RECT -66.805 -22.605 -66.475 -22.275 ;
        RECT -66.805 -23.965 -66.475 -23.635 ;
        RECT -66.805 -25.325 -66.475 -24.995 ;
        RECT -66.805 -26.685 -66.475 -26.355 ;
        RECT -66.805 -28.045 -66.475 -27.715 ;
        RECT -66.805 -29.405 -66.475 -29.075 ;
        RECT -66.805 -30.765 -66.475 -30.435 ;
        RECT -66.805 -32.125 -66.475 -31.795 ;
        RECT -66.805 -33.485 -66.475 -33.155 ;
        RECT -66.805 -34.845 -66.475 -34.515 ;
        RECT -66.805 -36.205 -66.475 -35.875 ;
        RECT -66.805 -37.565 -66.475 -37.235 ;
        RECT -66.805 -38.925 -66.475 -38.595 ;
        RECT -66.805 -40.285 -66.475 -39.955 ;
        RECT -66.805 -41.645 -66.475 -41.315 ;
        RECT -66.805 -43.005 -66.475 -42.675 ;
        RECT -66.805 -44.365 -66.475 -44.035 ;
        RECT -66.805 -45.725 -66.475 -45.395 ;
        RECT -66.805 -47.085 -66.475 -46.755 ;
        RECT -66.805 -48.445 -66.475 -48.115 ;
        RECT -66.805 -49.805 -66.475 -49.475 ;
        RECT -66.805 -51.165 -66.475 -50.835 ;
        RECT -66.805 -52.525 -66.475 -52.195 ;
        RECT -66.805 -53.885 -66.475 -53.555 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 205.875 129.8 206.205 130.93 ;
        RECT 205.875 127.675 206.205 128.005 ;
        RECT 205.875 126.315 206.205 126.645 ;
        RECT 205.875 124.955 206.205 125.285 ;
        RECT 205.875 123.595 206.205 123.925 ;
        RECT 205.875 122.215 206.205 122.545 ;
        RECT 205.875 120.165 206.205 120.495 ;
        RECT 205.875 118.235 206.205 118.565 ;
        RECT 205.875 116.395 206.205 116.725 ;
        RECT 205.875 114.905 206.205 115.235 ;
        RECT 205.875 113.235 206.205 113.565 ;
        RECT 205.875 111.745 206.205 112.075 ;
        RECT 205.875 110.075 206.205 110.405 ;
        RECT 205.875 108.585 206.205 108.915 ;
        RECT 205.875 106.915 206.205 107.245 ;
        RECT 205.875 105.425 206.205 105.755 ;
        RECT 205.875 104.015 206.205 104.345 ;
        RECT 205.875 102.175 206.205 102.505 ;
        RECT 205.875 100.685 206.205 101.015 ;
        RECT 205.875 99.015 206.205 99.345 ;
        RECT 205.875 97.525 206.205 97.855 ;
        RECT 205.875 95.855 206.205 96.185 ;
        RECT 205.875 94.365 206.205 94.695 ;
        RECT 205.875 92.695 206.205 93.025 ;
        RECT 205.875 91.205 206.205 91.535 ;
        RECT 205.875 89.795 206.205 90.125 ;
        RECT 205.875 87.955 206.205 88.285 ;
        RECT 205.875 86.465 206.205 86.795 ;
        RECT 205.875 84.795 206.205 85.125 ;
        RECT 205.875 83.305 206.205 83.635 ;
        RECT 205.875 81.635 206.205 81.965 ;
        RECT 205.875 80.145 206.205 80.475 ;
        RECT 205.875 78.475 206.205 78.805 ;
        RECT 205.875 76.985 206.205 77.315 ;
        RECT 205.875 75.575 206.205 75.905 ;
        RECT 205.875 73.735 206.205 74.065 ;
        RECT 205.875 72.245 206.205 72.575 ;
        RECT 205.875 70.575 206.205 70.905 ;
        RECT 205.875 69.085 206.205 69.415 ;
        RECT 205.875 67.415 206.205 67.745 ;
        RECT 205.875 65.925 206.205 66.255 ;
        RECT 205.875 64.255 206.205 64.585 ;
        RECT 205.875 62.765 206.205 63.095 ;
        RECT 205.875 61.355 206.205 61.685 ;
        RECT 205.875 59.515 206.205 59.845 ;
        RECT 205.875 58.025 206.205 58.355 ;
        RECT 205.875 56.355 206.205 56.685 ;
        RECT 205.875 54.865 206.205 55.195 ;
        RECT 205.875 53.195 206.205 53.525 ;
        RECT 205.875 51.705 206.205 52.035 ;
        RECT 205.875 50.035 206.205 50.365 ;
        RECT 205.875 48.545 206.205 48.875 ;
        RECT 205.875 47.135 206.205 47.465 ;
        RECT 205.875 45.295 206.205 45.625 ;
        RECT 205.875 43.805 206.205 44.135 ;
        RECT 205.875 42.135 206.205 42.465 ;
        RECT 205.875 40.645 206.205 40.975 ;
        RECT 205.875 38.975 206.205 39.305 ;
        RECT 205.875 37.485 206.205 37.815 ;
        RECT 205.875 35.815 206.205 36.145 ;
        RECT 205.875 34.325 206.205 34.655 ;
        RECT 205.875 32.915 206.205 33.245 ;
        RECT 205.875 31.075 206.205 31.405 ;
        RECT 205.875 29.585 206.205 29.915 ;
        RECT 205.875 27.915 206.205 28.245 ;
        RECT 205.875 26.425 206.205 26.755 ;
        RECT 205.875 24.755 206.205 25.085 ;
        RECT 205.875 23.265 206.205 23.595 ;
        RECT 205.875 21.595 206.205 21.925 ;
        RECT 205.875 20.105 206.205 20.435 ;
        RECT 205.875 18.695 206.205 19.025 ;
        RECT 205.875 16.855 206.205 17.185 ;
        RECT 205.875 15.365 206.205 15.695 ;
        RECT 205.875 13.695 206.205 14.025 ;
        RECT 205.875 12.205 206.205 12.535 ;
        RECT 205.875 10.535 206.205 10.865 ;
        RECT 205.875 9.045 206.205 9.375 ;
        RECT 205.875 7.375 206.205 7.705 ;
        RECT 205.875 5.885 206.205 6.215 ;
        RECT 205.875 4.475 206.205 4.805 ;
        RECT 205.875 2.115 206.205 2.445 ;
        RECT 205.875 0.06 206.205 0.39 ;
        RECT 205.875 -1.525 206.205 -1.195 ;
        RECT 205.875 -2.885 206.205 -2.555 ;
        RECT 205.875 -4.245 206.205 -3.915 ;
        RECT 205.875 -5.605 206.205 -5.275 ;
        RECT 205.875 -6.965 206.205 -6.635 ;
        RECT 205.875 -8.325 206.205 -7.995 ;
        RECT 205.875 -9.685 206.205 -9.355 ;
        RECT 205.875 -11.045 206.205 -10.715 ;
        RECT 205.875 -12.405 206.205 -12.075 ;
        RECT 205.875 -13.765 206.205 -13.435 ;
        RECT 205.875 -15.125 206.205 -14.795 ;
        RECT 205.875 -16.485 206.205 -16.155 ;
        RECT 205.875 -17.845 206.205 -17.515 ;
        RECT 205.875 -19.205 206.205 -18.875 ;
        RECT 205.875 -20.565 206.205 -20.235 ;
        RECT 205.875 -21.925 206.205 -21.595 ;
        RECT 205.875 -23.285 206.205 -22.955 ;
        RECT 205.875 -24.645 206.205 -24.315 ;
        RECT 205.875 -26.005 206.205 -25.675 ;
        RECT 205.875 -27.365 206.205 -27.035 ;
        RECT 205.875 -28.725 206.205 -28.395 ;
        RECT 205.875 -30.085 206.205 -29.755 ;
        RECT 205.875 -31.445 206.205 -31.115 ;
        RECT 205.875 -32.805 206.205 -32.475 ;
        RECT 205.875 -34.165 206.205 -33.835 ;
        RECT 205.875 -35.525 206.205 -35.195 ;
        RECT 205.875 -36.885 206.205 -36.555 ;
        RECT 205.875 -38.245 206.205 -37.915 ;
        RECT 205.875 -39.605 206.205 -39.275 ;
        RECT 205.875 -40.965 206.205 -40.635 ;
        RECT 205.875 -42.325 206.205 -41.995 ;
        RECT 205.875 -43.685 206.205 -43.355 ;
        RECT 205.875 -45.045 206.205 -44.715 ;
        RECT 205.875 -46.405 206.205 -46.075 ;
        RECT 205.875 -47.765 206.205 -47.435 ;
        RECT 205.875 -49.125 206.205 -48.795 ;
        RECT 205.875 -50.485 206.205 -50.155 ;
        RECT 205.875 -51.845 206.205 -51.515 ;
        RECT 205.875 -53.205 206.205 -52.875 ;
        RECT 205.875 -54.565 206.205 -54.235 ;
        RECT 205.875 -55.925 206.205 -55.595 ;
        RECT 205.875 -57.285 206.205 -56.955 ;
        RECT 205.875 -58.645 206.205 -58.315 ;
        RECT 205.875 -60.005 206.205 -59.675 ;
        RECT 205.875 -61.365 206.205 -61.035 ;
        RECT 205.875 -62.725 206.205 -62.395 ;
        RECT 205.875 -64.085 206.205 -63.755 ;
        RECT 205.875 -65.445 206.205 -65.115 ;
        RECT 205.875 -66.805 206.205 -66.475 ;
        RECT 205.875 -68.165 206.205 -67.835 ;
        RECT 205.875 -69.525 206.205 -69.195 ;
        RECT 205.875 -70.885 206.205 -70.555 ;
        RECT 205.875 -72.245 206.205 -71.915 ;
        RECT 205.875 -73.605 206.205 -73.275 ;
        RECT 205.875 -74.965 206.205 -74.635 ;
        RECT 205.875 -76.325 206.205 -75.995 ;
        RECT 205.875 -77.685 206.205 -77.355 ;
        RECT 205.875 -79.045 206.205 -78.715 ;
        RECT 205.875 -80.405 206.205 -80.075 ;
        RECT 205.875 -81.765 206.205 -81.435 ;
        RECT 205.875 -83.125 206.205 -82.795 ;
        RECT 205.875 -84.485 206.205 -84.155 ;
        RECT 205.875 -85.845 206.205 -85.515 ;
        RECT 205.875 -87.205 206.205 -86.875 ;
        RECT 205.875 -88.565 206.205 -88.235 ;
        RECT 205.875 -89.925 206.205 -89.595 ;
        RECT 205.875 -91.285 206.205 -90.955 ;
        RECT 205.875 -92.645 206.205 -92.315 ;
        RECT 205.875 -94.005 206.205 -93.675 ;
        RECT 205.875 -95.365 206.205 -95.035 ;
        RECT 205.875 -96.725 206.205 -96.395 ;
        RECT 205.875 -98.085 206.205 -97.755 ;
        RECT 205.875 -99.445 206.205 -99.115 ;
        RECT 205.875 -100.805 206.205 -100.475 ;
        RECT 205.875 -102.165 206.205 -101.835 ;
        RECT 205.875 -103.525 206.205 -103.195 ;
        RECT 205.875 -104.885 206.205 -104.555 ;
        RECT 205.875 -106.245 206.205 -105.915 ;
        RECT 205.875 -107.605 206.205 -107.275 ;
        RECT 205.875 -108.965 206.205 -108.635 ;
        RECT 205.875 -110.325 206.205 -109.995 ;
        RECT 205.875 -111.685 206.205 -111.355 ;
        RECT 205.875 -113.045 206.205 -112.715 ;
        RECT 205.875 -114.405 206.205 -114.075 ;
        RECT 205.875 -115.765 206.205 -115.435 ;
        RECT 205.875 -117.125 206.205 -116.795 ;
        RECT 205.875 -118.485 206.205 -118.155 ;
        RECT 205.875 -119.845 206.205 -119.515 ;
        RECT 205.875 -121.205 206.205 -120.875 ;
        RECT 205.875 -122.565 206.205 -122.235 ;
        RECT 205.875 -123.925 206.205 -123.595 ;
        RECT 205.875 -125.285 206.205 -124.955 ;
        RECT 205.875 -126.645 206.205 -126.315 ;
        RECT 205.875 -128.005 206.205 -127.675 ;
        RECT 205.875 -129.365 206.205 -129.035 ;
        RECT 205.875 -130.725 206.205 -130.395 ;
        RECT 205.875 -132.085 206.205 -131.755 ;
        RECT 205.875 -133.445 206.205 -133.115 ;
        RECT 205.875 -134.805 206.205 -134.475 ;
        RECT 205.875 -136.165 206.205 -135.835 ;
        RECT 205.875 -137.525 206.205 -137.195 ;
        RECT 205.875 -138.885 206.205 -138.555 ;
        RECT 205.875 -140.245 206.205 -139.915 ;
        RECT 205.875 -141.605 206.205 -141.275 ;
        RECT 205.875 -142.965 206.205 -142.635 ;
        RECT 205.875 -144.325 206.205 -143.995 ;
        RECT 205.875 -145.685 206.205 -145.355 ;
        RECT 205.875 -147.045 206.205 -146.715 ;
        RECT 205.875 -148.405 206.205 -148.075 ;
        RECT 205.875 -149.765 206.205 -149.435 ;
        RECT 205.875 -151.125 206.205 -150.795 ;
        RECT 205.875 -152.485 206.205 -152.155 ;
        RECT 205.875 -153.845 206.205 -153.515 ;
        RECT 205.875 -155.205 206.205 -154.875 ;
        RECT 205.875 -156.565 206.205 -156.235 ;
        RECT 205.875 -157.925 206.205 -157.595 ;
        RECT 205.875 -159.285 206.205 -158.955 ;
        RECT 205.875 -160.645 206.205 -160.315 ;
        RECT 205.875 -162.005 206.205 -161.675 ;
        RECT 205.875 -163.365 206.205 -163.035 ;
        RECT 205.875 -164.725 206.205 -164.395 ;
        RECT 205.875 -166.085 206.205 -165.755 ;
        RECT 205.875 -167.445 206.205 -167.115 ;
        RECT 205.875 -168.805 206.205 -168.475 ;
        RECT 205.875 -170.165 206.205 -169.835 ;
        RECT 205.875 -171.525 206.205 -171.195 ;
        RECT 205.875 -172.885 206.205 -172.555 ;
        RECT 205.875 -174.245 206.205 -173.915 ;
        RECT 205.875 -175.605 206.205 -175.275 ;
        RECT 205.875 -176.965 206.205 -176.635 ;
        RECT 205.875 -178.325 206.205 -177.995 ;
        RECT 205.875 -179.685 206.205 -179.355 ;
        RECT 205.875 -181.045 206.205 -180.715 ;
        RECT 205.875 -182.405 206.205 -182.075 ;
        RECT 205.875 -183.765 206.205 -183.435 ;
        RECT 205.875 -185.125 206.205 -184.795 ;
        RECT 205.875 -186.485 206.205 -186.155 ;
        RECT 205.875 -187.845 206.205 -187.515 ;
        RECT 205.875 -189.205 206.205 -188.875 ;
        RECT 205.875 -190.565 206.205 -190.235 ;
        RECT 205.875 -191.925 206.205 -191.595 ;
        RECT 205.875 -193.285 206.205 -192.955 ;
        RECT 205.875 -194.645 206.205 -194.315 ;
        RECT 205.875 -196.005 206.205 -195.675 ;
        RECT 205.875 -197.365 206.205 -197.035 ;
        RECT 205.875 -198.725 206.205 -198.395 ;
        RECT 205.875 -200.085 206.205 -199.755 ;
        RECT 205.875 -201.445 206.205 -201.115 ;
        RECT 205.875 -202.805 206.205 -202.475 ;
        RECT 205.875 -204.165 206.205 -203.835 ;
        RECT 205.875 -205.525 206.205 -205.195 ;
        RECT 205.875 -206.885 206.205 -206.555 ;
        RECT 205.875 -208.245 206.205 -207.915 ;
        RECT 205.875 -209.605 206.205 -209.275 ;
        RECT 205.875 -210.965 206.205 -210.635 ;
        RECT 205.875 -212.325 206.205 -211.995 ;
        RECT 205.875 -213.685 206.205 -213.355 ;
        RECT 205.875 -215.045 206.205 -214.715 ;
        RECT 205.875 -216.405 206.205 -216.075 ;
        RECT 205.875 -217.765 206.205 -217.435 ;
        RECT 205.875 -219.125 206.205 -218.795 ;
        RECT 205.875 -221.37 206.205 -220.24 ;
        RECT 205.88 -221.485 206.2 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.235 129.8 207.565 130.93 ;
        RECT 207.235 127.675 207.565 128.005 ;
        RECT 207.235 126.315 207.565 126.645 ;
        RECT 207.235 124.955 207.565 125.285 ;
        RECT 207.235 123.595 207.565 123.925 ;
        RECT 207.235 -1.525 207.565 -1.195 ;
        RECT 207.235 -2.885 207.565 -2.555 ;
        RECT 207.235 -4.245 207.565 -3.915 ;
        RECT 207.235 -5.605 207.565 -5.275 ;
        RECT 207.235 -6.965 207.565 -6.635 ;
        RECT 207.235 -8.325 207.565 -7.995 ;
        RECT 207.235 -9.685 207.565 -9.355 ;
        RECT 207.235 -11.045 207.565 -10.715 ;
        RECT 207.235 -12.405 207.565 -12.075 ;
        RECT 207.235 -13.765 207.565 -13.435 ;
        RECT 207.235 -15.125 207.565 -14.795 ;
        RECT 207.235 -16.485 207.565 -16.155 ;
        RECT 207.235 -17.845 207.565 -17.515 ;
        RECT 207.235 -19.205 207.565 -18.875 ;
        RECT 207.235 -20.565 207.565 -20.235 ;
        RECT 207.235 -21.925 207.565 -21.595 ;
        RECT 207.235 -23.285 207.565 -22.955 ;
        RECT 207.235 -24.645 207.565 -24.315 ;
        RECT 207.235 -26.005 207.565 -25.675 ;
        RECT 207.235 -27.365 207.565 -27.035 ;
        RECT 207.235 -28.725 207.565 -28.395 ;
        RECT 207.235 -30.085 207.565 -29.755 ;
        RECT 207.235 -31.445 207.565 -31.115 ;
        RECT 207.235 -32.805 207.565 -32.475 ;
        RECT 207.235 -34.165 207.565 -33.835 ;
        RECT 207.235 -35.525 207.565 -35.195 ;
        RECT 207.235 -36.885 207.565 -36.555 ;
        RECT 207.235 -38.245 207.565 -37.915 ;
        RECT 207.235 -39.605 207.565 -39.275 ;
        RECT 207.235 -40.965 207.565 -40.635 ;
        RECT 207.235 -42.325 207.565 -41.995 ;
        RECT 207.235 -43.685 207.565 -43.355 ;
        RECT 207.235 -45.045 207.565 -44.715 ;
        RECT 207.235 -46.405 207.565 -46.075 ;
        RECT 207.235 -47.765 207.565 -47.435 ;
        RECT 207.235 -49.125 207.565 -48.795 ;
        RECT 207.235 -50.485 207.565 -50.155 ;
        RECT 207.235 -51.845 207.565 -51.515 ;
        RECT 207.235 -53.205 207.565 -52.875 ;
        RECT 207.235 -54.565 207.565 -54.235 ;
        RECT 207.235 -55.925 207.565 -55.595 ;
        RECT 207.235 -57.285 207.565 -56.955 ;
        RECT 207.235 -58.645 207.565 -58.315 ;
        RECT 207.235 -60.005 207.565 -59.675 ;
        RECT 207.235 -61.365 207.565 -61.035 ;
        RECT 207.235 -62.725 207.565 -62.395 ;
        RECT 207.235 -64.085 207.565 -63.755 ;
        RECT 207.235 -65.445 207.565 -65.115 ;
        RECT 207.235 -66.805 207.565 -66.475 ;
        RECT 207.235 -68.165 207.565 -67.835 ;
        RECT 207.235 -69.525 207.565 -69.195 ;
        RECT 207.235 -70.885 207.565 -70.555 ;
        RECT 207.235 -72.245 207.565 -71.915 ;
        RECT 207.235 -73.605 207.565 -73.275 ;
        RECT 207.235 -74.965 207.565 -74.635 ;
        RECT 207.235 -76.325 207.565 -75.995 ;
        RECT 207.235 -77.685 207.565 -77.355 ;
        RECT 207.235 -79.045 207.565 -78.715 ;
        RECT 207.235 -80.405 207.565 -80.075 ;
        RECT 207.235 -81.765 207.565 -81.435 ;
        RECT 207.235 -83.125 207.565 -82.795 ;
        RECT 207.235 -84.485 207.565 -84.155 ;
        RECT 207.235 -85.845 207.565 -85.515 ;
        RECT 207.235 -87.205 207.565 -86.875 ;
        RECT 207.235 -88.565 207.565 -88.235 ;
        RECT 207.235 -89.925 207.565 -89.595 ;
        RECT 207.235 -91.285 207.565 -90.955 ;
        RECT 207.235 -92.645 207.565 -92.315 ;
        RECT 207.235 -94.005 207.565 -93.675 ;
        RECT 207.235 -95.365 207.565 -95.035 ;
        RECT 207.235 -96.725 207.565 -96.395 ;
        RECT 207.235 -98.085 207.565 -97.755 ;
        RECT 207.235 -99.445 207.565 -99.115 ;
        RECT 207.235 -100.805 207.565 -100.475 ;
        RECT 207.235 -102.165 207.565 -101.835 ;
        RECT 207.235 -103.525 207.565 -103.195 ;
        RECT 207.235 -104.885 207.565 -104.555 ;
        RECT 207.235 -106.245 207.565 -105.915 ;
        RECT 207.235 -107.605 207.565 -107.275 ;
        RECT 207.235 -108.965 207.565 -108.635 ;
        RECT 207.235 -110.325 207.565 -109.995 ;
        RECT 207.235 -111.685 207.565 -111.355 ;
        RECT 207.235 -113.045 207.565 -112.715 ;
        RECT 207.235 -114.405 207.565 -114.075 ;
        RECT 207.235 -115.765 207.565 -115.435 ;
        RECT 207.235 -117.125 207.565 -116.795 ;
        RECT 207.235 -118.485 207.565 -118.155 ;
        RECT 207.235 -119.845 207.565 -119.515 ;
        RECT 207.235 -121.205 207.565 -120.875 ;
        RECT 207.235 -122.565 207.565 -122.235 ;
        RECT 207.235 -123.925 207.565 -123.595 ;
        RECT 207.235 -125.285 207.565 -124.955 ;
        RECT 207.235 -126.645 207.565 -126.315 ;
        RECT 207.235 -128.005 207.565 -127.675 ;
        RECT 207.235 -129.365 207.565 -129.035 ;
        RECT 207.235 -130.725 207.565 -130.395 ;
        RECT 207.235 -132.085 207.565 -131.755 ;
        RECT 207.235 -133.445 207.565 -133.115 ;
        RECT 207.235 -134.805 207.565 -134.475 ;
        RECT 207.235 -136.165 207.565 -135.835 ;
        RECT 207.235 -137.525 207.565 -137.195 ;
        RECT 207.235 -138.885 207.565 -138.555 ;
        RECT 207.235 -140.245 207.565 -139.915 ;
        RECT 207.235 -141.605 207.565 -141.275 ;
        RECT 207.235 -142.965 207.565 -142.635 ;
        RECT 207.235 -144.325 207.565 -143.995 ;
        RECT 207.235 -145.685 207.565 -145.355 ;
        RECT 207.235 -147.045 207.565 -146.715 ;
        RECT 207.235 -148.405 207.565 -148.075 ;
        RECT 207.235 -149.765 207.565 -149.435 ;
        RECT 207.235 -151.125 207.565 -150.795 ;
        RECT 207.235 -152.485 207.565 -152.155 ;
        RECT 207.235 -153.845 207.565 -153.515 ;
        RECT 207.235 -155.205 207.565 -154.875 ;
        RECT 207.235 -156.565 207.565 -156.235 ;
        RECT 207.235 -157.925 207.565 -157.595 ;
        RECT 207.235 -159.285 207.565 -158.955 ;
        RECT 207.235 -160.645 207.565 -160.315 ;
        RECT 207.235 -162.005 207.565 -161.675 ;
        RECT 207.235 -163.365 207.565 -163.035 ;
        RECT 207.235 -164.725 207.565 -164.395 ;
        RECT 207.235 -166.085 207.565 -165.755 ;
        RECT 207.235 -167.445 207.565 -167.115 ;
        RECT 207.235 -168.805 207.565 -168.475 ;
        RECT 207.235 -170.165 207.565 -169.835 ;
        RECT 207.235 -171.525 207.565 -171.195 ;
        RECT 207.235 -172.885 207.565 -172.555 ;
        RECT 207.235 -174.245 207.565 -173.915 ;
        RECT 207.235 -175.605 207.565 -175.275 ;
        RECT 207.235 -176.965 207.565 -176.635 ;
        RECT 207.235 -178.325 207.565 -177.995 ;
        RECT 207.235 -179.685 207.565 -179.355 ;
        RECT 207.235 -181.045 207.565 -180.715 ;
        RECT 207.235 -182.405 207.565 -182.075 ;
        RECT 207.235 -183.765 207.565 -183.435 ;
        RECT 207.235 -185.125 207.565 -184.795 ;
        RECT 207.235 -186.485 207.565 -186.155 ;
        RECT 207.235 -187.845 207.565 -187.515 ;
        RECT 207.235 -189.205 207.565 -188.875 ;
        RECT 207.235 -190.565 207.565 -190.235 ;
        RECT 207.235 -191.925 207.565 -191.595 ;
        RECT 207.235 -193.285 207.565 -192.955 ;
        RECT 207.235 -194.645 207.565 -194.315 ;
        RECT 207.235 -196.005 207.565 -195.675 ;
        RECT 207.235 -197.365 207.565 -197.035 ;
        RECT 207.235 -198.725 207.565 -198.395 ;
        RECT 207.235 -200.085 207.565 -199.755 ;
        RECT 207.235 -201.445 207.565 -201.115 ;
        RECT 207.235 -202.805 207.565 -202.475 ;
        RECT 207.235 -204.165 207.565 -203.835 ;
        RECT 207.235 -205.525 207.565 -205.195 ;
        RECT 207.235 -206.885 207.565 -206.555 ;
        RECT 207.235 -208.245 207.565 -207.915 ;
        RECT 207.235 -209.605 207.565 -209.275 ;
        RECT 207.235 -210.965 207.565 -210.635 ;
        RECT 207.235 -212.325 207.565 -211.995 ;
        RECT 207.235 -213.685 207.565 -213.355 ;
        RECT 207.235 -215.045 207.565 -214.715 ;
        RECT 207.235 -216.405 207.565 -216.075 ;
        RECT 207.235 -217.765 207.565 -217.435 ;
        RECT 207.235 -219.125 207.565 -218.795 ;
        RECT 207.235 -221.37 207.565 -220.24 ;
        RECT 207.24 -221.485 207.56 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 208.595 129.8 208.925 130.93 ;
        RECT 208.595 127.675 208.925 128.005 ;
        RECT 208.595 126.315 208.925 126.645 ;
        RECT 208.595 124.955 208.925 125.285 ;
        RECT 208.595 123.595 208.925 123.925 ;
        RECT 208.595 122.235 208.925 122.565 ;
        RECT 208.595 120.875 208.925 121.205 ;
        RECT 208.595 119.515 208.925 119.845 ;
        RECT 208.595 118.155 208.925 118.485 ;
        RECT 208.595 116.795 208.925 117.125 ;
        RECT 208.595 115.435 208.925 115.765 ;
        RECT 208.595 114.075 208.925 114.405 ;
        RECT 208.595 112.715 208.925 113.045 ;
        RECT 208.595 111.355 208.925 111.685 ;
        RECT 208.595 109.995 208.925 110.325 ;
        RECT 208.595 108.635 208.925 108.965 ;
        RECT 208.595 107.275 208.925 107.605 ;
        RECT 208.595 105.915 208.925 106.245 ;
        RECT 208.595 104.555 208.925 104.885 ;
        RECT 208.595 103.195 208.925 103.525 ;
        RECT 208.595 101.835 208.925 102.165 ;
        RECT 208.595 100.475 208.925 100.805 ;
        RECT 208.595 99.115 208.925 99.445 ;
        RECT 208.595 97.755 208.925 98.085 ;
        RECT 208.595 96.395 208.925 96.725 ;
        RECT 208.595 95.035 208.925 95.365 ;
        RECT 208.595 93.675 208.925 94.005 ;
        RECT 208.595 92.315 208.925 92.645 ;
        RECT 208.595 90.955 208.925 91.285 ;
        RECT 208.595 89.595 208.925 89.925 ;
        RECT 208.595 88.235 208.925 88.565 ;
        RECT 208.595 86.875 208.925 87.205 ;
        RECT 208.595 85.515 208.925 85.845 ;
        RECT 208.595 84.155 208.925 84.485 ;
        RECT 208.595 82.795 208.925 83.125 ;
        RECT 208.595 81.435 208.925 81.765 ;
        RECT 208.595 80.075 208.925 80.405 ;
        RECT 208.595 78.715 208.925 79.045 ;
        RECT 208.595 77.355 208.925 77.685 ;
        RECT 208.595 75.995 208.925 76.325 ;
        RECT 208.595 74.635 208.925 74.965 ;
        RECT 208.595 73.275 208.925 73.605 ;
        RECT 208.595 71.915 208.925 72.245 ;
        RECT 208.595 70.555 208.925 70.885 ;
        RECT 208.595 69.195 208.925 69.525 ;
        RECT 208.595 67.835 208.925 68.165 ;
        RECT 208.595 66.475 208.925 66.805 ;
        RECT 208.595 65.115 208.925 65.445 ;
        RECT 208.595 63.755 208.925 64.085 ;
        RECT 208.595 62.395 208.925 62.725 ;
        RECT 208.595 61.035 208.925 61.365 ;
        RECT 208.595 59.675 208.925 60.005 ;
        RECT 208.595 58.315 208.925 58.645 ;
        RECT 208.595 56.955 208.925 57.285 ;
        RECT 208.595 55.595 208.925 55.925 ;
        RECT 208.595 54.235 208.925 54.565 ;
        RECT 208.595 52.875 208.925 53.205 ;
        RECT 208.595 51.515 208.925 51.845 ;
        RECT 208.595 50.155 208.925 50.485 ;
        RECT 208.595 48.795 208.925 49.125 ;
        RECT 208.595 47.435 208.925 47.765 ;
        RECT 208.595 46.075 208.925 46.405 ;
        RECT 208.595 44.715 208.925 45.045 ;
        RECT 208.595 43.355 208.925 43.685 ;
        RECT 208.595 41.995 208.925 42.325 ;
        RECT 208.595 40.635 208.925 40.965 ;
        RECT 208.595 39.275 208.925 39.605 ;
        RECT 208.595 37.915 208.925 38.245 ;
        RECT 208.595 36.555 208.925 36.885 ;
        RECT 208.595 35.195 208.925 35.525 ;
        RECT 208.595 33.835 208.925 34.165 ;
        RECT 208.595 32.475 208.925 32.805 ;
        RECT 208.595 31.115 208.925 31.445 ;
        RECT 208.595 29.755 208.925 30.085 ;
        RECT 208.595 28.395 208.925 28.725 ;
        RECT 208.595 27.035 208.925 27.365 ;
        RECT 208.595 25.675 208.925 26.005 ;
        RECT 208.595 24.315 208.925 24.645 ;
        RECT 208.595 22.955 208.925 23.285 ;
        RECT 208.595 21.595 208.925 21.925 ;
        RECT 208.595 20.235 208.925 20.565 ;
        RECT 208.595 18.875 208.925 19.205 ;
        RECT 208.595 17.515 208.925 17.845 ;
        RECT 208.595 16.155 208.925 16.485 ;
        RECT 208.595 14.795 208.925 15.125 ;
        RECT 208.595 13.435 208.925 13.765 ;
        RECT 208.595 12.075 208.925 12.405 ;
        RECT 208.595 10.715 208.925 11.045 ;
        RECT 208.595 9.355 208.925 9.685 ;
        RECT 208.595 7.995 208.925 8.325 ;
        RECT 208.595 6.635 208.925 6.965 ;
        RECT 208.595 5.275 208.925 5.605 ;
        RECT 208.595 3.915 208.925 4.245 ;
        RECT 208.595 2.555 208.925 2.885 ;
        RECT 208.595 1.195 208.925 1.525 ;
        RECT 208.595 -0.165 208.925 0.165 ;
        RECT 208.595 -1.525 208.925 -1.195 ;
        RECT 208.595 -2.885 208.925 -2.555 ;
        RECT 208.595 -4.245 208.925 -3.915 ;
        RECT 208.595 -5.605 208.925 -5.275 ;
        RECT 208.595 -6.965 208.925 -6.635 ;
        RECT 208.595 -8.325 208.925 -7.995 ;
        RECT 208.595 -9.685 208.925 -9.355 ;
        RECT 208.595 -11.045 208.925 -10.715 ;
        RECT 208.595 -12.405 208.925 -12.075 ;
        RECT 208.595 -13.765 208.925 -13.435 ;
        RECT 208.595 -15.125 208.925 -14.795 ;
        RECT 208.595 -16.485 208.925 -16.155 ;
        RECT 208.595 -17.845 208.925 -17.515 ;
        RECT 208.595 -19.205 208.925 -18.875 ;
        RECT 208.595 -20.565 208.925 -20.235 ;
        RECT 208.595 -21.925 208.925 -21.595 ;
        RECT 208.595 -23.285 208.925 -22.955 ;
        RECT 208.595 -24.645 208.925 -24.315 ;
        RECT 208.595 -26.005 208.925 -25.675 ;
        RECT 208.595 -27.365 208.925 -27.035 ;
        RECT 208.595 -28.725 208.925 -28.395 ;
        RECT 208.595 -30.085 208.925 -29.755 ;
        RECT 208.595 -31.445 208.925 -31.115 ;
        RECT 208.595 -32.805 208.925 -32.475 ;
        RECT 208.595 -34.165 208.925 -33.835 ;
        RECT 208.595 -35.525 208.925 -35.195 ;
        RECT 208.595 -36.885 208.925 -36.555 ;
        RECT 208.595 -38.245 208.925 -37.915 ;
        RECT 208.595 -39.605 208.925 -39.275 ;
        RECT 208.595 -40.965 208.925 -40.635 ;
        RECT 208.595 -42.325 208.925 -41.995 ;
        RECT 208.595 -43.685 208.925 -43.355 ;
        RECT 208.595 -45.045 208.925 -44.715 ;
        RECT 208.595 -46.405 208.925 -46.075 ;
        RECT 208.595 -47.765 208.925 -47.435 ;
        RECT 208.595 -49.125 208.925 -48.795 ;
        RECT 208.595 -50.485 208.925 -50.155 ;
        RECT 208.595 -51.845 208.925 -51.515 ;
        RECT 208.595 -53.205 208.925 -52.875 ;
        RECT 208.595 -54.565 208.925 -54.235 ;
        RECT 208.595 -55.925 208.925 -55.595 ;
        RECT 208.595 -57.285 208.925 -56.955 ;
        RECT 208.595 -58.645 208.925 -58.315 ;
        RECT 208.595 -60.005 208.925 -59.675 ;
        RECT 208.595 -61.365 208.925 -61.035 ;
        RECT 208.595 -62.725 208.925 -62.395 ;
        RECT 208.595 -64.085 208.925 -63.755 ;
        RECT 208.595 -65.445 208.925 -65.115 ;
        RECT 208.595 -66.805 208.925 -66.475 ;
        RECT 208.595 -68.165 208.925 -67.835 ;
        RECT 208.595 -69.525 208.925 -69.195 ;
        RECT 208.595 -70.885 208.925 -70.555 ;
        RECT 208.595 -72.245 208.925 -71.915 ;
        RECT 208.595 -73.605 208.925 -73.275 ;
        RECT 208.595 -74.965 208.925 -74.635 ;
        RECT 208.595 -76.325 208.925 -75.995 ;
        RECT 208.595 -77.685 208.925 -77.355 ;
        RECT 208.595 -79.045 208.925 -78.715 ;
        RECT 208.595 -80.405 208.925 -80.075 ;
        RECT 208.595 -81.765 208.925 -81.435 ;
        RECT 208.595 -83.125 208.925 -82.795 ;
        RECT 208.595 -84.485 208.925 -84.155 ;
        RECT 208.595 -85.845 208.925 -85.515 ;
        RECT 208.595 -87.205 208.925 -86.875 ;
        RECT 208.595 -88.565 208.925 -88.235 ;
        RECT 208.595 -89.925 208.925 -89.595 ;
        RECT 208.595 -91.285 208.925 -90.955 ;
        RECT 208.595 -92.645 208.925 -92.315 ;
        RECT 208.595 -94.005 208.925 -93.675 ;
        RECT 208.595 -95.365 208.925 -95.035 ;
        RECT 208.595 -96.725 208.925 -96.395 ;
        RECT 208.595 -98.085 208.925 -97.755 ;
        RECT 208.595 -99.445 208.925 -99.115 ;
        RECT 208.595 -100.805 208.925 -100.475 ;
        RECT 208.595 -102.165 208.925 -101.835 ;
        RECT 208.595 -103.525 208.925 -103.195 ;
        RECT 208.595 -104.885 208.925 -104.555 ;
        RECT 208.595 -106.245 208.925 -105.915 ;
        RECT 208.595 -107.605 208.925 -107.275 ;
        RECT 208.595 -108.965 208.925 -108.635 ;
        RECT 208.595 -110.325 208.925 -109.995 ;
        RECT 208.595 -111.685 208.925 -111.355 ;
        RECT 208.595 -113.045 208.925 -112.715 ;
        RECT 208.595 -114.405 208.925 -114.075 ;
        RECT 208.595 -115.765 208.925 -115.435 ;
        RECT 208.595 -117.125 208.925 -116.795 ;
        RECT 208.595 -118.485 208.925 -118.155 ;
        RECT 208.595 -119.845 208.925 -119.515 ;
        RECT 208.595 -121.205 208.925 -120.875 ;
        RECT 208.595 -122.565 208.925 -122.235 ;
        RECT 208.595 -123.925 208.925 -123.595 ;
        RECT 208.595 -125.285 208.925 -124.955 ;
        RECT 208.595 -126.645 208.925 -126.315 ;
        RECT 208.595 -128.005 208.925 -127.675 ;
        RECT 208.595 -129.365 208.925 -129.035 ;
        RECT 208.595 -130.725 208.925 -130.395 ;
        RECT 208.595 -132.085 208.925 -131.755 ;
        RECT 208.595 -133.445 208.925 -133.115 ;
        RECT 208.595 -134.805 208.925 -134.475 ;
        RECT 208.595 -136.165 208.925 -135.835 ;
        RECT 208.595 -137.525 208.925 -137.195 ;
        RECT 208.595 -138.885 208.925 -138.555 ;
        RECT 208.595 -140.245 208.925 -139.915 ;
        RECT 208.595 -141.605 208.925 -141.275 ;
        RECT 208.595 -142.965 208.925 -142.635 ;
        RECT 208.595 -144.325 208.925 -143.995 ;
        RECT 208.595 -145.685 208.925 -145.355 ;
        RECT 208.595 -147.045 208.925 -146.715 ;
        RECT 208.595 -148.405 208.925 -148.075 ;
        RECT 208.595 -149.765 208.925 -149.435 ;
        RECT 208.595 -151.125 208.925 -150.795 ;
        RECT 208.595 -152.485 208.925 -152.155 ;
        RECT 208.595 -153.845 208.925 -153.515 ;
        RECT 208.595 -155.205 208.925 -154.875 ;
        RECT 208.595 -156.565 208.925 -156.235 ;
        RECT 208.595 -157.925 208.925 -157.595 ;
        RECT 208.595 -159.285 208.925 -158.955 ;
        RECT 208.595 -160.645 208.925 -160.315 ;
        RECT 208.595 -162.005 208.925 -161.675 ;
        RECT 208.595 -163.365 208.925 -163.035 ;
        RECT 208.595 -164.725 208.925 -164.395 ;
        RECT 208.595 -166.085 208.925 -165.755 ;
        RECT 208.595 -167.445 208.925 -167.115 ;
        RECT 208.595 -168.805 208.925 -168.475 ;
        RECT 208.595 -170.165 208.925 -169.835 ;
        RECT 208.595 -171.525 208.925 -171.195 ;
        RECT 208.595 -172.885 208.925 -172.555 ;
        RECT 208.595 -174.245 208.925 -173.915 ;
        RECT 208.595 -175.605 208.925 -175.275 ;
        RECT 208.595 -176.965 208.925 -176.635 ;
        RECT 208.595 -178.325 208.925 -177.995 ;
        RECT 208.595 -179.685 208.925 -179.355 ;
        RECT 208.595 -181.045 208.925 -180.715 ;
        RECT 208.595 -182.405 208.925 -182.075 ;
        RECT 208.595 -183.765 208.925 -183.435 ;
        RECT 208.595 -185.125 208.925 -184.795 ;
        RECT 208.595 -186.485 208.925 -186.155 ;
        RECT 208.595 -187.845 208.925 -187.515 ;
        RECT 208.595 -189.205 208.925 -188.875 ;
        RECT 208.595 -190.565 208.925 -190.235 ;
        RECT 208.595 -191.925 208.925 -191.595 ;
        RECT 208.595 -193.285 208.925 -192.955 ;
        RECT 208.595 -194.645 208.925 -194.315 ;
        RECT 208.595 -196.005 208.925 -195.675 ;
        RECT 208.595 -197.365 208.925 -197.035 ;
        RECT 208.595 -198.725 208.925 -198.395 ;
        RECT 208.595 -200.085 208.925 -199.755 ;
        RECT 208.595 -201.445 208.925 -201.115 ;
        RECT 208.595 -202.805 208.925 -202.475 ;
        RECT 208.595 -204.165 208.925 -203.835 ;
        RECT 208.595 -205.525 208.925 -205.195 ;
        RECT 208.595 -206.885 208.925 -206.555 ;
        RECT 208.595 -208.245 208.925 -207.915 ;
        RECT 208.595 -209.605 208.925 -209.275 ;
        RECT 208.595 -210.965 208.925 -210.635 ;
        RECT 208.595 -212.325 208.925 -211.995 ;
        RECT 208.595 -213.685 208.925 -213.355 ;
        RECT 208.595 -215.045 208.925 -214.715 ;
        RECT 208.595 -216.405 208.925 -216.075 ;
        RECT 208.595 -217.765 208.925 -217.435 ;
        RECT 208.595 -219.125 208.925 -218.795 ;
        RECT 208.595 -221.37 208.925 -220.24 ;
        RECT 208.6 -221.485 208.92 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.955 129.8 210.285 130.93 ;
        RECT 209.955 127.675 210.285 128.005 ;
        RECT 209.955 126.315 210.285 126.645 ;
        RECT 209.955 124.955 210.285 125.285 ;
        RECT 209.955 123.595 210.285 123.925 ;
        RECT 209.955 122.235 210.285 122.565 ;
        RECT 209.955 120.875 210.285 121.205 ;
        RECT 209.955 119.515 210.285 119.845 ;
        RECT 209.955 118.155 210.285 118.485 ;
        RECT 209.955 116.795 210.285 117.125 ;
        RECT 209.955 115.435 210.285 115.765 ;
        RECT 209.955 114.075 210.285 114.405 ;
        RECT 209.955 112.715 210.285 113.045 ;
        RECT 209.955 111.355 210.285 111.685 ;
        RECT 209.955 109.995 210.285 110.325 ;
        RECT 209.955 108.635 210.285 108.965 ;
        RECT 209.955 107.275 210.285 107.605 ;
        RECT 209.955 105.915 210.285 106.245 ;
        RECT 209.955 104.555 210.285 104.885 ;
        RECT 209.955 103.195 210.285 103.525 ;
        RECT 209.955 101.835 210.285 102.165 ;
        RECT 209.955 100.475 210.285 100.805 ;
        RECT 209.955 99.115 210.285 99.445 ;
        RECT 209.955 97.755 210.285 98.085 ;
        RECT 209.955 96.395 210.285 96.725 ;
        RECT 209.955 95.035 210.285 95.365 ;
        RECT 209.955 93.675 210.285 94.005 ;
        RECT 209.955 92.315 210.285 92.645 ;
        RECT 209.955 90.955 210.285 91.285 ;
        RECT 209.955 89.595 210.285 89.925 ;
        RECT 209.955 88.235 210.285 88.565 ;
        RECT 209.955 86.875 210.285 87.205 ;
        RECT 209.955 85.515 210.285 85.845 ;
        RECT 209.955 84.155 210.285 84.485 ;
        RECT 209.955 82.795 210.285 83.125 ;
        RECT 209.955 81.435 210.285 81.765 ;
        RECT 209.955 80.075 210.285 80.405 ;
        RECT 209.955 78.715 210.285 79.045 ;
        RECT 209.955 77.355 210.285 77.685 ;
        RECT 209.955 75.995 210.285 76.325 ;
        RECT 209.955 74.635 210.285 74.965 ;
        RECT 209.955 73.275 210.285 73.605 ;
        RECT 209.955 71.915 210.285 72.245 ;
        RECT 209.955 70.555 210.285 70.885 ;
        RECT 209.955 69.195 210.285 69.525 ;
        RECT 209.955 67.835 210.285 68.165 ;
        RECT 209.955 66.475 210.285 66.805 ;
        RECT 209.955 65.115 210.285 65.445 ;
        RECT 209.955 63.755 210.285 64.085 ;
        RECT 209.955 62.395 210.285 62.725 ;
        RECT 209.955 61.035 210.285 61.365 ;
        RECT 209.955 59.675 210.285 60.005 ;
        RECT 209.955 58.315 210.285 58.645 ;
        RECT 209.955 56.955 210.285 57.285 ;
        RECT 209.955 55.595 210.285 55.925 ;
        RECT 209.955 54.235 210.285 54.565 ;
        RECT 209.955 52.875 210.285 53.205 ;
        RECT 209.955 51.515 210.285 51.845 ;
        RECT 209.955 50.155 210.285 50.485 ;
        RECT 209.955 48.795 210.285 49.125 ;
        RECT 209.955 47.435 210.285 47.765 ;
        RECT 209.955 46.075 210.285 46.405 ;
        RECT 209.955 44.715 210.285 45.045 ;
        RECT 209.955 43.355 210.285 43.685 ;
        RECT 209.955 41.995 210.285 42.325 ;
        RECT 209.955 40.635 210.285 40.965 ;
        RECT 209.955 39.275 210.285 39.605 ;
        RECT 209.955 37.915 210.285 38.245 ;
        RECT 209.955 36.555 210.285 36.885 ;
        RECT 209.955 35.195 210.285 35.525 ;
        RECT 209.955 33.835 210.285 34.165 ;
        RECT 209.955 32.475 210.285 32.805 ;
        RECT 209.955 31.115 210.285 31.445 ;
        RECT 209.955 29.755 210.285 30.085 ;
        RECT 209.955 28.395 210.285 28.725 ;
        RECT 209.955 27.035 210.285 27.365 ;
        RECT 209.955 25.675 210.285 26.005 ;
        RECT 209.955 24.315 210.285 24.645 ;
        RECT 209.955 22.955 210.285 23.285 ;
        RECT 209.955 21.595 210.285 21.925 ;
        RECT 209.955 20.235 210.285 20.565 ;
        RECT 209.955 18.875 210.285 19.205 ;
        RECT 209.955 17.515 210.285 17.845 ;
        RECT 209.955 16.155 210.285 16.485 ;
        RECT 209.955 14.795 210.285 15.125 ;
        RECT 209.955 13.435 210.285 13.765 ;
        RECT 209.955 12.075 210.285 12.405 ;
        RECT 209.955 10.715 210.285 11.045 ;
        RECT 209.955 9.355 210.285 9.685 ;
        RECT 209.955 7.995 210.285 8.325 ;
        RECT 209.955 6.635 210.285 6.965 ;
        RECT 209.955 5.275 210.285 5.605 ;
        RECT 209.955 3.915 210.285 4.245 ;
        RECT 209.955 2.555 210.285 2.885 ;
        RECT 209.955 1.195 210.285 1.525 ;
        RECT 209.955 -0.165 210.285 0.165 ;
        RECT 209.955 -1.525 210.285 -1.195 ;
        RECT 209.955 -2.885 210.285 -2.555 ;
        RECT 209.955 -4.245 210.285 -3.915 ;
        RECT 209.955 -5.605 210.285 -5.275 ;
        RECT 209.955 -6.965 210.285 -6.635 ;
        RECT 209.955 -8.325 210.285 -7.995 ;
        RECT 209.955 -9.685 210.285 -9.355 ;
        RECT 209.955 -11.045 210.285 -10.715 ;
        RECT 209.955 -12.405 210.285 -12.075 ;
        RECT 209.955 -13.765 210.285 -13.435 ;
        RECT 209.955 -15.125 210.285 -14.795 ;
        RECT 209.955 -16.485 210.285 -16.155 ;
        RECT 209.955 -17.845 210.285 -17.515 ;
        RECT 209.955 -19.205 210.285 -18.875 ;
        RECT 209.955 -20.565 210.285 -20.235 ;
        RECT 209.955 -21.925 210.285 -21.595 ;
        RECT 209.955 -23.285 210.285 -22.955 ;
        RECT 209.955 -24.645 210.285 -24.315 ;
        RECT 209.955 -26.005 210.285 -25.675 ;
        RECT 209.955 -27.365 210.285 -27.035 ;
        RECT 209.955 -28.725 210.285 -28.395 ;
        RECT 209.955 -30.085 210.285 -29.755 ;
        RECT 209.955 -31.445 210.285 -31.115 ;
        RECT 209.955 -32.805 210.285 -32.475 ;
        RECT 209.955 -34.165 210.285 -33.835 ;
        RECT 209.955 -35.525 210.285 -35.195 ;
        RECT 209.955 -36.885 210.285 -36.555 ;
        RECT 209.955 -38.245 210.285 -37.915 ;
        RECT 209.955 -39.605 210.285 -39.275 ;
        RECT 209.955 -40.965 210.285 -40.635 ;
        RECT 209.955 -42.325 210.285 -41.995 ;
        RECT 209.955 -43.685 210.285 -43.355 ;
        RECT 209.955 -45.045 210.285 -44.715 ;
        RECT 209.955 -46.405 210.285 -46.075 ;
        RECT 209.955 -47.765 210.285 -47.435 ;
        RECT 209.955 -49.125 210.285 -48.795 ;
        RECT 209.955 -50.485 210.285 -50.155 ;
        RECT 209.955 -51.845 210.285 -51.515 ;
        RECT 209.955 -53.205 210.285 -52.875 ;
        RECT 209.955 -54.565 210.285 -54.235 ;
        RECT 209.955 -55.925 210.285 -55.595 ;
        RECT 209.955 -57.285 210.285 -56.955 ;
        RECT 209.955 -58.645 210.285 -58.315 ;
        RECT 209.955 -60.005 210.285 -59.675 ;
        RECT 209.955 -61.365 210.285 -61.035 ;
        RECT 209.955 -62.725 210.285 -62.395 ;
        RECT 209.955 -64.085 210.285 -63.755 ;
        RECT 209.955 -65.445 210.285 -65.115 ;
        RECT 209.955 -66.805 210.285 -66.475 ;
        RECT 209.955 -68.165 210.285 -67.835 ;
        RECT 209.955 -69.525 210.285 -69.195 ;
        RECT 209.955 -70.885 210.285 -70.555 ;
        RECT 209.955 -72.245 210.285 -71.915 ;
        RECT 209.955 -73.605 210.285 -73.275 ;
        RECT 209.955 -74.965 210.285 -74.635 ;
        RECT 209.955 -76.325 210.285 -75.995 ;
        RECT 209.955 -77.685 210.285 -77.355 ;
        RECT 209.955 -79.045 210.285 -78.715 ;
        RECT 209.955 -80.405 210.285 -80.075 ;
        RECT 209.955 -81.765 210.285 -81.435 ;
        RECT 209.955 -83.125 210.285 -82.795 ;
        RECT 209.955 -84.485 210.285 -84.155 ;
        RECT 209.955 -85.845 210.285 -85.515 ;
        RECT 209.955 -87.205 210.285 -86.875 ;
        RECT 209.955 -88.565 210.285 -88.235 ;
        RECT 209.955 -89.925 210.285 -89.595 ;
        RECT 209.955 -91.285 210.285 -90.955 ;
        RECT 209.955 -92.645 210.285 -92.315 ;
        RECT 209.955 -94.005 210.285 -93.675 ;
        RECT 209.955 -95.365 210.285 -95.035 ;
        RECT 209.955 -96.725 210.285 -96.395 ;
        RECT 209.955 -98.085 210.285 -97.755 ;
        RECT 209.955 -99.445 210.285 -99.115 ;
        RECT 209.955 -100.805 210.285 -100.475 ;
        RECT 209.955 -102.165 210.285 -101.835 ;
        RECT 209.955 -103.525 210.285 -103.195 ;
        RECT 209.955 -104.885 210.285 -104.555 ;
        RECT 209.955 -106.245 210.285 -105.915 ;
        RECT 209.955 -107.605 210.285 -107.275 ;
        RECT 209.955 -108.965 210.285 -108.635 ;
        RECT 209.955 -110.325 210.285 -109.995 ;
        RECT 209.955 -111.685 210.285 -111.355 ;
        RECT 209.955 -113.045 210.285 -112.715 ;
        RECT 209.955 -114.405 210.285 -114.075 ;
        RECT 209.955 -115.765 210.285 -115.435 ;
        RECT 209.955 -117.125 210.285 -116.795 ;
        RECT 209.955 -118.485 210.285 -118.155 ;
        RECT 209.955 -119.845 210.285 -119.515 ;
        RECT 209.955 -121.205 210.285 -120.875 ;
        RECT 209.955 -122.565 210.285 -122.235 ;
        RECT 209.955 -123.925 210.285 -123.595 ;
        RECT 209.955 -125.285 210.285 -124.955 ;
        RECT 209.955 -126.645 210.285 -126.315 ;
        RECT 209.955 -128.005 210.285 -127.675 ;
        RECT 209.955 -129.365 210.285 -129.035 ;
        RECT 209.955 -130.725 210.285 -130.395 ;
        RECT 209.955 -132.085 210.285 -131.755 ;
        RECT 209.955 -133.445 210.285 -133.115 ;
        RECT 209.955 -134.805 210.285 -134.475 ;
        RECT 209.955 -136.165 210.285 -135.835 ;
        RECT 209.955 -137.525 210.285 -137.195 ;
        RECT 209.955 -138.885 210.285 -138.555 ;
        RECT 209.955 -140.245 210.285 -139.915 ;
        RECT 209.955 -141.605 210.285 -141.275 ;
        RECT 209.955 -142.965 210.285 -142.635 ;
        RECT 209.955 -144.325 210.285 -143.995 ;
        RECT 209.955 -145.685 210.285 -145.355 ;
        RECT 209.955 -147.045 210.285 -146.715 ;
        RECT 209.955 -148.405 210.285 -148.075 ;
        RECT 209.955 -149.765 210.285 -149.435 ;
        RECT 209.955 -151.125 210.285 -150.795 ;
        RECT 209.955 -152.485 210.285 -152.155 ;
        RECT 209.955 -153.845 210.285 -153.515 ;
        RECT 209.955 -155.205 210.285 -154.875 ;
        RECT 209.955 -156.565 210.285 -156.235 ;
        RECT 209.955 -157.925 210.285 -157.595 ;
        RECT 209.955 -159.285 210.285 -158.955 ;
        RECT 209.955 -160.645 210.285 -160.315 ;
        RECT 209.955 -162.005 210.285 -161.675 ;
        RECT 209.955 -163.365 210.285 -163.035 ;
        RECT 209.955 -164.725 210.285 -164.395 ;
        RECT 209.955 -166.085 210.285 -165.755 ;
        RECT 209.955 -167.445 210.285 -167.115 ;
        RECT 209.955 -168.805 210.285 -168.475 ;
        RECT 209.955 -170.165 210.285 -169.835 ;
        RECT 209.955 -171.525 210.285 -171.195 ;
        RECT 209.955 -172.885 210.285 -172.555 ;
        RECT 209.955 -174.245 210.285 -173.915 ;
        RECT 209.955 -175.605 210.285 -175.275 ;
        RECT 209.955 -176.965 210.285 -176.635 ;
        RECT 209.955 -178.325 210.285 -177.995 ;
        RECT 209.955 -179.685 210.285 -179.355 ;
        RECT 209.955 -181.045 210.285 -180.715 ;
        RECT 209.955 -182.405 210.285 -182.075 ;
        RECT 209.955 -183.765 210.285 -183.435 ;
        RECT 209.955 -185.125 210.285 -184.795 ;
        RECT 209.955 -186.485 210.285 -186.155 ;
        RECT 209.955 -187.845 210.285 -187.515 ;
        RECT 209.955 -189.205 210.285 -188.875 ;
        RECT 209.955 -190.565 210.285 -190.235 ;
        RECT 209.955 -191.925 210.285 -191.595 ;
        RECT 209.955 -193.285 210.285 -192.955 ;
        RECT 209.955 -194.645 210.285 -194.315 ;
        RECT 209.955 -196.005 210.285 -195.675 ;
        RECT 209.955 -197.365 210.285 -197.035 ;
        RECT 209.955 -198.725 210.285 -198.395 ;
        RECT 209.955 -200.085 210.285 -199.755 ;
        RECT 209.955 -201.445 210.285 -201.115 ;
        RECT 209.955 -202.805 210.285 -202.475 ;
        RECT 209.955 -204.165 210.285 -203.835 ;
        RECT 209.955 -205.525 210.285 -205.195 ;
        RECT 209.955 -206.885 210.285 -206.555 ;
        RECT 209.955 -208.245 210.285 -207.915 ;
        RECT 209.955 -209.605 210.285 -209.275 ;
        RECT 209.955 -210.965 210.285 -210.635 ;
        RECT 209.955 -212.325 210.285 -211.995 ;
        RECT 209.955 -213.685 210.285 -213.355 ;
        RECT 209.955 -215.045 210.285 -214.715 ;
        RECT 209.955 -216.405 210.285 -216.075 ;
        RECT 209.955 -217.765 210.285 -217.435 ;
        RECT 209.955 -219.125 210.285 -218.795 ;
        RECT 209.96 -221.485 210.28 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.275 129.8 192.605 130.93 ;
        RECT 192.275 127.675 192.605 128.005 ;
        RECT 192.275 126.315 192.605 126.645 ;
        RECT 192.275 124.955 192.605 125.285 ;
        RECT 192.275 123.595 192.605 123.925 ;
        RECT 192.28 123.595 192.6 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.275 -122.565 192.605 -122.235 ;
        RECT 192.275 -123.925 192.605 -123.595 ;
        RECT 192.275 -125.285 192.605 -124.955 ;
        RECT 192.275 -126.645 192.605 -126.315 ;
        RECT 192.275 -128.005 192.605 -127.675 ;
        RECT 192.275 -129.365 192.605 -129.035 ;
        RECT 192.275 -130.725 192.605 -130.395 ;
        RECT 192.275 -132.085 192.605 -131.755 ;
        RECT 192.275 -133.445 192.605 -133.115 ;
        RECT 192.275 -134.805 192.605 -134.475 ;
        RECT 192.275 -136.165 192.605 -135.835 ;
        RECT 192.275 -137.525 192.605 -137.195 ;
        RECT 192.275 -138.885 192.605 -138.555 ;
        RECT 192.275 -140.245 192.605 -139.915 ;
        RECT 192.275 -141.605 192.605 -141.275 ;
        RECT 192.275 -142.965 192.605 -142.635 ;
        RECT 192.275 -144.325 192.605 -143.995 ;
        RECT 192.275 -145.685 192.605 -145.355 ;
        RECT 192.275 -147.045 192.605 -146.715 ;
        RECT 192.275 -148.405 192.605 -148.075 ;
        RECT 192.275 -149.765 192.605 -149.435 ;
        RECT 192.275 -151.125 192.605 -150.795 ;
        RECT 192.275 -152.485 192.605 -152.155 ;
        RECT 192.275 -153.845 192.605 -153.515 ;
        RECT 192.275 -155.205 192.605 -154.875 ;
        RECT 192.275 -156.565 192.605 -156.235 ;
        RECT 192.275 -157.925 192.605 -157.595 ;
        RECT 192.275 -159.285 192.605 -158.955 ;
        RECT 192.275 -160.645 192.605 -160.315 ;
        RECT 192.275 -162.005 192.605 -161.675 ;
        RECT 192.275 -163.365 192.605 -163.035 ;
        RECT 192.275 -164.725 192.605 -164.395 ;
        RECT 192.275 -166.085 192.605 -165.755 ;
        RECT 192.275 -167.445 192.605 -167.115 ;
        RECT 192.275 -168.805 192.605 -168.475 ;
        RECT 192.275 -170.165 192.605 -169.835 ;
        RECT 192.275 -171.525 192.605 -171.195 ;
        RECT 192.275 -172.885 192.605 -172.555 ;
        RECT 192.275 -174.245 192.605 -173.915 ;
        RECT 192.275 -175.605 192.605 -175.275 ;
        RECT 192.275 -176.965 192.605 -176.635 ;
        RECT 192.275 -178.325 192.605 -177.995 ;
        RECT 192.275 -179.685 192.605 -179.355 ;
        RECT 192.275 -181.045 192.605 -180.715 ;
        RECT 192.275 -182.405 192.605 -182.075 ;
        RECT 192.275 -183.765 192.605 -183.435 ;
        RECT 192.275 -185.125 192.605 -184.795 ;
        RECT 192.275 -186.485 192.605 -186.155 ;
        RECT 192.275 -187.845 192.605 -187.515 ;
        RECT 192.275 -189.205 192.605 -188.875 ;
        RECT 192.275 -190.565 192.605 -190.235 ;
        RECT 192.275 -191.925 192.605 -191.595 ;
        RECT 192.275 -193.285 192.605 -192.955 ;
        RECT 192.275 -194.645 192.605 -194.315 ;
        RECT 192.275 -196.005 192.605 -195.675 ;
        RECT 192.275 -197.365 192.605 -197.035 ;
        RECT 192.275 -198.725 192.605 -198.395 ;
        RECT 192.275 -200.085 192.605 -199.755 ;
        RECT 192.275 -201.445 192.605 -201.115 ;
        RECT 192.275 -202.805 192.605 -202.475 ;
        RECT 192.275 -204.165 192.605 -203.835 ;
        RECT 192.275 -205.525 192.605 -205.195 ;
        RECT 192.275 -206.885 192.605 -206.555 ;
        RECT 192.275 -208.245 192.605 -207.915 ;
        RECT 192.275 -209.605 192.605 -209.275 ;
        RECT 192.275 -210.965 192.605 -210.635 ;
        RECT 192.275 -212.325 192.605 -211.995 ;
        RECT 192.275 -213.685 192.605 -213.355 ;
        RECT 192.275 -215.045 192.605 -214.715 ;
        RECT 192.275 -216.405 192.605 -216.075 ;
        RECT 192.275 -217.765 192.605 -217.435 ;
        RECT 192.275 -219.125 192.605 -218.795 ;
        RECT 192.275 -221.37 192.605 -220.24 ;
        RECT 192.28 -221.485 192.6 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.41 -121.535 192.74 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.635 129.8 193.965 130.93 ;
        RECT 193.635 127.675 193.965 128.005 ;
        RECT 193.635 126.315 193.965 126.645 ;
        RECT 193.635 124.955 193.965 125.285 ;
        RECT 193.635 123.595 193.965 123.925 ;
        RECT 193.64 123.595 193.96 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.635 -1.525 193.965 -1.195 ;
        RECT 193.635 -2.885 193.965 -2.555 ;
        RECT 193.64 -3.56 193.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.995 129.8 195.325 130.93 ;
        RECT 194.995 127.675 195.325 128.005 ;
        RECT 194.995 126.315 195.325 126.645 ;
        RECT 194.995 124.955 195.325 125.285 ;
        RECT 194.995 123.595 195.325 123.925 ;
        RECT 195 123.595 195.32 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.995 -1.525 195.325 -1.195 ;
        RECT 194.995 -2.885 195.325 -2.555 ;
        RECT 195 -3.56 195.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.355 129.8 196.685 130.93 ;
        RECT 196.355 127.675 196.685 128.005 ;
        RECT 196.355 126.315 196.685 126.645 ;
        RECT 196.355 124.955 196.685 125.285 ;
        RECT 196.355 123.595 196.685 123.925 ;
        RECT 196.36 123.595 196.68 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.355 -1.525 196.685 -1.195 ;
        RECT 196.355 -2.885 196.685 -2.555 ;
        RECT 196.36 -3.56 196.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.355 -118.485 196.685 -118.155 ;
        RECT 196.355 -119.845 196.685 -119.515 ;
        RECT 196.355 -121.205 196.685 -120.875 ;
        RECT 196.355 -122.565 196.685 -122.235 ;
        RECT 196.355 -123.925 196.685 -123.595 ;
        RECT 196.355 -125.285 196.685 -124.955 ;
        RECT 196.355 -126.645 196.685 -126.315 ;
        RECT 196.355 -128.005 196.685 -127.675 ;
        RECT 196.355 -129.365 196.685 -129.035 ;
        RECT 196.355 -130.725 196.685 -130.395 ;
        RECT 196.355 -132.085 196.685 -131.755 ;
        RECT 196.355 -133.445 196.685 -133.115 ;
        RECT 196.355 -134.805 196.685 -134.475 ;
        RECT 196.355 -136.165 196.685 -135.835 ;
        RECT 196.355 -137.525 196.685 -137.195 ;
        RECT 196.355 -138.885 196.685 -138.555 ;
        RECT 196.355 -140.245 196.685 -139.915 ;
        RECT 196.355 -141.605 196.685 -141.275 ;
        RECT 196.355 -142.965 196.685 -142.635 ;
        RECT 196.355 -144.325 196.685 -143.995 ;
        RECT 196.355 -145.685 196.685 -145.355 ;
        RECT 196.355 -147.045 196.685 -146.715 ;
        RECT 196.355 -148.405 196.685 -148.075 ;
        RECT 196.355 -149.765 196.685 -149.435 ;
        RECT 196.355 -151.125 196.685 -150.795 ;
        RECT 196.355 -152.485 196.685 -152.155 ;
        RECT 196.355 -153.845 196.685 -153.515 ;
        RECT 196.355 -155.205 196.685 -154.875 ;
        RECT 196.355 -156.565 196.685 -156.235 ;
        RECT 196.355 -157.925 196.685 -157.595 ;
        RECT 196.355 -159.285 196.685 -158.955 ;
        RECT 196.355 -160.645 196.685 -160.315 ;
        RECT 196.355 -162.005 196.685 -161.675 ;
        RECT 196.355 -163.365 196.685 -163.035 ;
        RECT 196.355 -164.725 196.685 -164.395 ;
        RECT 196.355 -166.085 196.685 -165.755 ;
        RECT 196.355 -167.445 196.685 -167.115 ;
        RECT 196.355 -168.805 196.685 -168.475 ;
        RECT 196.355 -170.165 196.685 -169.835 ;
        RECT 196.355 -171.525 196.685 -171.195 ;
        RECT 196.355 -172.885 196.685 -172.555 ;
        RECT 196.355 -174.245 196.685 -173.915 ;
        RECT 196.355 -175.605 196.685 -175.275 ;
        RECT 196.355 -176.965 196.685 -176.635 ;
        RECT 196.355 -178.325 196.685 -177.995 ;
        RECT 196.355 -179.685 196.685 -179.355 ;
        RECT 196.355 -181.045 196.685 -180.715 ;
        RECT 196.355 -182.405 196.685 -182.075 ;
        RECT 196.355 -183.765 196.685 -183.435 ;
        RECT 196.355 -185.125 196.685 -184.795 ;
        RECT 196.355 -186.485 196.685 -186.155 ;
        RECT 196.355 -187.845 196.685 -187.515 ;
        RECT 196.355 -189.205 196.685 -188.875 ;
        RECT 196.355 -190.565 196.685 -190.235 ;
        RECT 196.355 -191.925 196.685 -191.595 ;
        RECT 196.355 -193.285 196.685 -192.955 ;
        RECT 196.355 -194.645 196.685 -194.315 ;
        RECT 196.355 -196.005 196.685 -195.675 ;
        RECT 196.355 -197.365 196.685 -197.035 ;
        RECT 196.355 -198.725 196.685 -198.395 ;
        RECT 196.355 -200.085 196.685 -199.755 ;
        RECT 196.355 -201.445 196.685 -201.115 ;
        RECT 196.355 -202.805 196.685 -202.475 ;
        RECT 196.355 -204.165 196.685 -203.835 ;
        RECT 196.355 -205.525 196.685 -205.195 ;
        RECT 196.355 -206.885 196.685 -206.555 ;
        RECT 196.355 -208.245 196.685 -207.915 ;
        RECT 196.355 -209.605 196.685 -209.275 ;
        RECT 196.355 -210.965 196.685 -210.635 ;
        RECT 196.355 -212.325 196.685 -211.995 ;
        RECT 196.355 -213.685 196.685 -213.355 ;
        RECT 196.355 -215.045 196.685 -214.715 ;
        RECT 196.355 -216.405 196.685 -216.075 ;
        RECT 196.355 -217.765 196.685 -217.435 ;
        RECT 196.355 -219.125 196.685 -218.795 ;
        RECT 196.355 -221.37 196.685 -220.24 ;
        RECT 196.36 -221.485 196.68 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.715 129.8 198.045 130.93 ;
        RECT 197.715 127.675 198.045 128.005 ;
        RECT 197.715 126.315 198.045 126.645 ;
        RECT 197.715 124.955 198.045 125.285 ;
        RECT 197.715 123.595 198.045 123.925 ;
        RECT 197.72 123.595 198.04 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.715 -122.565 198.045 -122.235 ;
        RECT 197.715 -123.925 198.045 -123.595 ;
        RECT 197.715 -125.285 198.045 -124.955 ;
        RECT 197.715 -126.645 198.045 -126.315 ;
        RECT 197.715 -128.005 198.045 -127.675 ;
        RECT 197.715 -129.365 198.045 -129.035 ;
        RECT 197.715 -130.725 198.045 -130.395 ;
        RECT 197.715 -132.085 198.045 -131.755 ;
        RECT 197.715 -133.445 198.045 -133.115 ;
        RECT 197.715 -134.805 198.045 -134.475 ;
        RECT 197.715 -136.165 198.045 -135.835 ;
        RECT 197.715 -137.525 198.045 -137.195 ;
        RECT 197.715 -138.885 198.045 -138.555 ;
        RECT 197.715 -140.245 198.045 -139.915 ;
        RECT 197.715 -141.605 198.045 -141.275 ;
        RECT 197.715 -142.965 198.045 -142.635 ;
        RECT 197.715 -144.325 198.045 -143.995 ;
        RECT 197.715 -145.685 198.045 -145.355 ;
        RECT 197.715 -147.045 198.045 -146.715 ;
        RECT 197.715 -148.405 198.045 -148.075 ;
        RECT 197.715 -149.765 198.045 -149.435 ;
        RECT 197.715 -151.125 198.045 -150.795 ;
        RECT 197.715 -152.485 198.045 -152.155 ;
        RECT 197.715 -153.845 198.045 -153.515 ;
        RECT 197.715 -155.205 198.045 -154.875 ;
        RECT 197.715 -156.565 198.045 -156.235 ;
        RECT 197.715 -157.925 198.045 -157.595 ;
        RECT 197.715 -159.285 198.045 -158.955 ;
        RECT 197.715 -160.645 198.045 -160.315 ;
        RECT 197.715 -162.005 198.045 -161.675 ;
        RECT 197.715 -163.365 198.045 -163.035 ;
        RECT 197.715 -164.725 198.045 -164.395 ;
        RECT 197.715 -166.085 198.045 -165.755 ;
        RECT 197.715 -167.445 198.045 -167.115 ;
        RECT 197.715 -168.805 198.045 -168.475 ;
        RECT 197.715 -170.165 198.045 -169.835 ;
        RECT 197.715 -171.525 198.045 -171.195 ;
        RECT 197.715 -172.885 198.045 -172.555 ;
        RECT 197.715 -174.245 198.045 -173.915 ;
        RECT 197.715 -175.605 198.045 -175.275 ;
        RECT 197.715 -176.965 198.045 -176.635 ;
        RECT 197.715 -178.325 198.045 -177.995 ;
        RECT 197.715 -179.685 198.045 -179.355 ;
        RECT 197.715 -181.045 198.045 -180.715 ;
        RECT 197.715 -182.405 198.045 -182.075 ;
        RECT 197.715 -183.765 198.045 -183.435 ;
        RECT 197.715 -185.125 198.045 -184.795 ;
        RECT 197.715 -186.485 198.045 -186.155 ;
        RECT 197.715 -187.845 198.045 -187.515 ;
        RECT 197.715 -189.205 198.045 -188.875 ;
        RECT 197.715 -190.565 198.045 -190.235 ;
        RECT 197.715 -191.925 198.045 -191.595 ;
        RECT 197.715 -193.285 198.045 -192.955 ;
        RECT 197.715 -194.645 198.045 -194.315 ;
        RECT 197.715 -196.005 198.045 -195.675 ;
        RECT 197.715 -197.365 198.045 -197.035 ;
        RECT 197.715 -198.725 198.045 -198.395 ;
        RECT 197.715 -200.085 198.045 -199.755 ;
        RECT 197.715 -201.445 198.045 -201.115 ;
        RECT 197.715 -202.805 198.045 -202.475 ;
        RECT 197.715 -204.165 198.045 -203.835 ;
        RECT 197.715 -205.525 198.045 -205.195 ;
        RECT 197.715 -206.885 198.045 -206.555 ;
        RECT 197.715 -208.245 198.045 -207.915 ;
        RECT 197.715 -209.605 198.045 -209.275 ;
        RECT 197.715 -210.965 198.045 -210.635 ;
        RECT 197.715 -212.325 198.045 -211.995 ;
        RECT 197.715 -213.685 198.045 -213.355 ;
        RECT 197.715 -215.045 198.045 -214.715 ;
        RECT 197.715 -216.405 198.045 -216.075 ;
        RECT 197.715 -217.765 198.045 -217.435 ;
        RECT 197.715 -219.125 198.045 -218.795 ;
        RECT 197.715 -221.37 198.045 -220.24 ;
        RECT 197.72 -221.485 198.04 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.86 -121.535 198.19 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.075 129.8 199.405 130.93 ;
        RECT 199.075 127.675 199.405 128.005 ;
        RECT 199.075 126.315 199.405 126.645 ;
        RECT 199.075 124.955 199.405 125.285 ;
        RECT 199.075 123.595 199.405 123.925 ;
        RECT 199.08 123.595 199.4 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.075 -122.565 199.405 -122.235 ;
        RECT 199.075 -123.925 199.405 -123.595 ;
        RECT 199.075 -125.285 199.405 -124.955 ;
        RECT 199.075 -126.645 199.405 -126.315 ;
        RECT 199.075 -128.005 199.405 -127.675 ;
        RECT 199.075 -129.365 199.405 -129.035 ;
        RECT 199.075 -130.725 199.405 -130.395 ;
        RECT 199.075 -132.085 199.405 -131.755 ;
        RECT 199.075 -133.445 199.405 -133.115 ;
        RECT 199.075 -134.805 199.405 -134.475 ;
        RECT 199.075 -136.165 199.405 -135.835 ;
        RECT 199.075 -137.525 199.405 -137.195 ;
        RECT 199.075 -138.885 199.405 -138.555 ;
        RECT 199.075 -140.245 199.405 -139.915 ;
        RECT 199.075 -141.605 199.405 -141.275 ;
        RECT 199.075 -142.965 199.405 -142.635 ;
        RECT 199.075 -144.325 199.405 -143.995 ;
        RECT 199.075 -145.685 199.405 -145.355 ;
        RECT 199.075 -147.045 199.405 -146.715 ;
        RECT 199.075 -148.405 199.405 -148.075 ;
        RECT 199.075 -149.765 199.405 -149.435 ;
        RECT 199.075 -151.125 199.405 -150.795 ;
        RECT 199.075 -152.485 199.405 -152.155 ;
        RECT 199.075 -153.845 199.405 -153.515 ;
        RECT 199.075 -155.205 199.405 -154.875 ;
        RECT 199.075 -156.565 199.405 -156.235 ;
        RECT 199.075 -157.925 199.405 -157.595 ;
        RECT 199.075 -159.285 199.405 -158.955 ;
        RECT 199.075 -160.645 199.405 -160.315 ;
        RECT 199.075 -162.005 199.405 -161.675 ;
        RECT 199.075 -163.365 199.405 -163.035 ;
        RECT 199.075 -164.725 199.405 -164.395 ;
        RECT 199.075 -166.085 199.405 -165.755 ;
        RECT 199.075 -167.445 199.405 -167.115 ;
        RECT 199.075 -168.805 199.405 -168.475 ;
        RECT 199.075 -170.165 199.405 -169.835 ;
        RECT 199.075 -171.525 199.405 -171.195 ;
        RECT 199.075 -172.885 199.405 -172.555 ;
        RECT 199.075 -174.245 199.405 -173.915 ;
        RECT 199.075 -175.605 199.405 -175.275 ;
        RECT 199.075 -176.965 199.405 -176.635 ;
        RECT 199.075 -178.325 199.405 -177.995 ;
        RECT 199.075 -179.685 199.405 -179.355 ;
        RECT 199.075 -181.045 199.405 -180.715 ;
        RECT 199.075 -182.405 199.405 -182.075 ;
        RECT 199.075 -183.765 199.405 -183.435 ;
        RECT 199.075 -185.125 199.405 -184.795 ;
        RECT 199.075 -186.485 199.405 -186.155 ;
        RECT 199.075 -187.845 199.405 -187.515 ;
        RECT 199.075 -189.205 199.405 -188.875 ;
        RECT 199.075 -190.565 199.405 -190.235 ;
        RECT 199.075 -191.925 199.405 -191.595 ;
        RECT 199.075 -193.285 199.405 -192.955 ;
        RECT 199.075 -194.645 199.405 -194.315 ;
        RECT 199.075 -196.005 199.405 -195.675 ;
        RECT 199.075 -197.365 199.405 -197.035 ;
        RECT 199.075 -198.725 199.405 -198.395 ;
        RECT 199.075 -200.085 199.405 -199.755 ;
        RECT 199.075 -201.445 199.405 -201.115 ;
        RECT 199.075 -202.805 199.405 -202.475 ;
        RECT 199.075 -204.165 199.405 -203.835 ;
        RECT 199.075 -205.525 199.405 -205.195 ;
        RECT 199.075 -206.885 199.405 -206.555 ;
        RECT 199.075 -208.245 199.405 -207.915 ;
        RECT 199.075 -209.605 199.405 -209.275 ;
        RECT 199.075 -210.965 199.405 -210.635 ;
        RECT 199.075 -212.325 199.405 -211.995 ;
        RECT 199.075 -213.685 199.405 -213.355 ;
        RECT 199.075 -215.045 199.405 -214.715 ;
        RECT 199.075 -216.405 199.405 -216.075 ;
        RECT 199.075 -217.765 199.405 -217.435 ;
        RECT 199.075 -219.125 199.405 -218.795 ;
        RECT 199.075 -221.37 199.405 -220.24 ;
        RECT 199.08 -221.485 199.4 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.435 129.8 200.765 130.93 ;
        RECT 200.435 127.675 200.765 128.005 ;
        RECT 200.435 126.315 200.765 126.645 ;
        RECT 200.435 124.955 200.765 125.285 ;
        RECT 200.435 123.595 200.765 123.925 ;
        RECT 200.44 123.595 200.76 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.435 -1.525 200.765 -1.195 ;
        RECT 200.435 -2.885 200.765 -2.555 ;
        RECT 200.44 -3.56 200.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.435 -118.485 200.765 -118.155 ;
        RECT 200.435 -119.845 200.765 -119.515 ;
        RECT 200.435 -121.205 200.765 -120.875 ;
        RECT 200.435 -122.565 200.765 -122.235 ;
        RECT 200.435 -123.925 200.765 -123.595 ;
        RECT 200.435 -125.285 200.765 -124.955 ;
        RECT 200.435 -126.645 200.765 -126.315 ;
        RECT 200.435 -128.005 200.765 -127.675 ;
        RECT 200.435 -129.365 200.765 -129.035 ;
        RECT 200.435 -130.725 200.765 -130.395 ;
        RECT 200.435 -132.085 200.765 -131.755 ;
        RECT 200.435 -133.445 200.765 -133.115 ;
        RECT 200.435 -134.805 200.765 -134.475 ;
        RECT 200.435 -136.165 200.765 -135.835 ;
        RECT 200.435 -137.525 200.765 -137.195 ;
        RECT 200.435 -138.885 200.765 -138.555 ;
        RECT 200.435 -140.245 200.765 -139.915 ;
        RECT 200.435 -141.605 200.765 -141.275 ;
        RECT 200.435 -142.965 200.765 -142.635 ;
        RECT 200.435 -144.325 200.765 -143.995 ;
        RECT 200.435 -145.685 200.765 -145.355 ;
        RECT 200.435 -147.045 200.765 -146.715 ;
        RECT 200.435 -148.405 200.765 -148.075 ;
        RECT 200.435 -149.765 200.765 -149.435 ;
        RECT 200.435 -151.125 200.765 -150.795 ;
        RECT 200.435 -152.485 200.765 -152.155 ;
        RECT 200.435 -153.845 200.765 -153.515 ;
        RECT 200.435 -155.205 200.765 -154.875 ;
        RECT 200.435 -156.565 200.765 -156.235 ;
        RECT 200.435 -157.925 200.765 -157.595 ;
        RECT 200.435 -159.285 200.765 -158.955 ;
        RECT 200.435 -160.645 200.765 -160.315 ;
        RECT 200.435 -162.005 200.765 -161.675 ;
        RECT 200.435 -163.365 200.765 -163.035 ;
        RECT 200.435 -164.725 200.765 -164.395 ;
        RECT 200.435 -166.085 200.765 -165.755 ;
        RECT 200.435 -167.445 200.765 -167.115 ;
        RECT 200.435 -168.805 200.765 -168.475 ;
        RECT 200.435 -170.165 200.765 -169.835 ;
        RECT 200.435 -171.525 200.765 -171.195 ;
        RECT 200.435 -172.885 200.765 -172.555 ;
        RECT 200.435 -174.245 200.765 -173.915 ;
        RECT 200.435 -175.605 200.765 -175.275 ;
        RECT 200.435 -176.965 200.765 -176.635 ;
        RECT 200.435 -178.325 200.765 -177.995 ;
        RECT 200.435 -179.685 200.765 -179.355 ;
        RECT 200.435 -181.045 200.765 -180.715 ;
        RECT 200.435 -182.405 200.765 -182.075 ;
        RECT 200.435 -183.765 200.765 -183.435 ;
        RECT 200.435 -185.125 200.765 -184.795 ;
        RECT 200.435 -186.485 200.765 -186.155 ;
        RECT 200.435 -187.845 200.765 -187.515 ;
        RECT 200.435 -189.205 200.765 -188.875 ;
        RECT 200.435 -190.565 200.765 -190.235 ;
        RECT 200.435 -191.925 200.765 -191.595 ;
        RECT 200.435 -193.285 200.765 -192.955 ;
        RECT 200.435 -194.645 200.765 -194.315 ;
        RECT 200.435 -196.005 200.765 -195.675 ;
        RECT 200.435 -197.365 200.765 -197.035 ;
        RECT 200.435 -198.725 200.765 -198.395 ;
        RECT 200.435 -200.085 200.765 -199.755 ;
        RECT 200.435 -201.445 200.765 -201.115 ;
        RECT 200.435 -202.805 200.765 -202.475 ;
        RECT 200.435 -204.165 200.765 -203.835 ;
        RECT 200.435 -205.525 200.765 -205.195 ;
        RECT 200.435 -206.885 200.765 -206.555 ;
        RECT 200.435 -208.245 200.765 -207.915 ;
        RECT 200.435 -209.605 200.765 -209.275 ;
        RECT 200.435 -210.965 200.765 -210.635 ;
        RECT 200.435 -212.325 200.765 -211.995 ;
        RECT 200.435 -213.685 200.765 -213.355 ;
        RECT 200.435 -215.045 200.765 -214.715 ;
        RECT 200.435 -216.405 200.765 -216.075 ;
        RECT 200.435 -217.765 200.765 -217.435 ;
        RECT 200.435 -219.125 200.765 -218.795 ;
        RECT 200.435 -221.37 200.765 -220.24 ;
        RECT 200.44 -221.485 200.76 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.795 129.8 202.125 130.93 ;
        RECT 201.795 127.675 202.125 128.005 ;
        RECT 201.795 126.315 202.125 126.645 ;
        RECT 201.795 124.955 202.125 125.285 ;
        RECT 201.795 123.595 202.125 123.925 ;
        RECT 201.8 123.595 202.12 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.795 -1.525 202.125 -1.195 ;
        RECT 201.795 -2.885 202.125 -2.555 ;
        RECT 201.8 -3.56 202.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.795 -118.485 202.125 -118.155 ;
        RECT 201.795 -119.845 202.125 -119.515 ;
        RECT 201.795 -121.205 202.125 -120.875 ;
        RECT 201.795 -122.565 202.125 -122.235 ;
        RECT 201.795 -123.925 202.125 -123.595 ;
        RECT 201.795 -125.285 202.125 -124.955 ;
        RECT 201.795 -126.645 202.125 -126.315 ;
        RECT 201.795 -128.005 202.125 -127.675 ;
        RECT 201.795 -129.365 202.125 -129.035 ;
        RECT 201.795 -130.725 202.125 -130.395 ;
        RECT 201.795 -132.085 202.125 -131.755 ;
        RECT 201.795 -133.445 202.125 -133.115 ;
        RECT 201.795 -134.805 202.125 -134.475 ;
        RECT 201.795 -136.165 202.125 -135.835 ;
        RECT 201.795 -137.525 202.125 -137.195 ;
        RECT 201.795 -138.885 202.125 -138.555 ;
        RECT 201.795 -140.245 202.125 -139.915 ;
        RECT 201.795 -141.605 202.125 -141.275 ;
        RECT 201.795 -142.965 202.125 -142.635 ;
        RECT 201.795 -144.325 202.125 -143.995 ;
        RECT 201.795 -145.685 202.125 -145.355 ;
        RECT 201.795 -147.045 202.125 -146.715 ;
        RECT 201.795 -148.405 202.125 -148.075 ;
        RECT 201.795 -149.765 202.125 -149.435 ;
        RECT 201.795 -151.125 202.125 -150.795 ;
        RECT 201.795 -152.485 202.125 -152.155 ;
        RECT 201.795 -153.845 202.125 -153.515 ;
        RECT 201.795 -155.205 202.125 -154.875 ;
        RECT 201.795 -156.565 202.125 -156.235 ;
        RECT 201.795 -157.925 202.125 -157.595 ;
        RECT 201.795 -159.285 202.125 -158.955 ;
        RECT 201.795 -160.645 202.125 -160.315 ;
        RECT 201.795 -162.005 202.125 -161.675 ;
        RECT 201.795 -163.365 202.125 -163.035 ;
        RECT 201.795 -164.725 202.125 -164.395 ;
        RECT 201.795 -166.085 202.125 -165.755 ;
        RECT 201.795 -167.445 202.125 -167.115 ;
        RECT 201.795 -168.805 202.125 -168.475 ;
        RECT 201.795 -170.165 202.125 -169.835 ;
        RECT 201.795 -171.525 202.125 -171.195 ;
        RECT 201.795 -172.885 202.125 -172.555 ;
        RECT 201.795 -174.245 202.125 -173.915 ;
        RECT 201.795 -175.605 202.125 -175.275 ;
        RECT 201.795 -176.965 202.125 -176.635 ;
        RECT 201.795 -178.325 202.125 -177.995 ;
        RECT 201.795 -179.685 202.125 -179.355 ;
        RECT 201.795 -181.045 202.125 -180.715 ;
        RECT 201.795 -182.405 202.125 -182.075 ;
        RECT 201.795 -183.765 202.125 -183.435 ;
        RECT 201.795 -185.125 202.125 -184.795 ;
        RECT 201.795 -186.485 202.125 -186.155 ;
        RECT 201.795 -187.845 202.125 -187.515 ;
        RECT 201.795 -189.205 202.125 -188.875 ;
        RECT 201.795 -190.565 202.125 -190.235 ;
        RECT 201.795 -191.925 202.125 -191.595 ;
        RECT 201.795 -193.285 202.125 -192.955 ;
        RECT 201.795 -194.645 202.125 -194.315 ;
        RECT 201.795 -196.005 202.125 -195.675 ;
        RECT 201.795 -197.365 202.125 -197.035 ;
        RECT 201.795 -198.725 202.125 -198.395 ;
        RECT 201.795 -200.085 202.125 -199.755 ;
        RECT 201.795 -201.445 202.125 -201.115 ;
        RECT 201.795 -202.805 202.125 -202.475 ;
        RECT 201.795 -204.165 202.125 -203.835 ;
        RECT 201.795 -205.525 202.125 -205.195 ;
        RECT 201.795 -206.885 202.125 -206.555 ;
        RECT 201.795 -208.245 202.125 -207.915 ;
        RECT 201.795 -209.605 202.125 -209.275 ;
        RECT 201.795 -210.965 202.125 -210.635 ;
        RECT 201.795 -212.325 202.125 -211.995 ;
        RECT 201.795 -213.685 202.125 -213.355 ;
        RECT 201.795 -215.045 202.125 -214.715 ;
        RECT 201.795 -216.405 202.125 -216.075 ;
        RECT 201.795 -217.765 202.125 -217.435 ;
        RECT 201.795 -219.125 202.125 -218.795 ;
        RECT 201.795 -221.37 202.125 -220.24 ;
        RECT 201.8 -221.485 202.12 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.155 129.8 203.485 130.93 ;
        RECT 203.155 127.675 203.485 128.005 ;
        RECT 203.155 126.315 203.485 126.645 ;
        RECT 203.155 124.955 203.485 125.285 ;
        RECT 203.155 123.595 203.485 123.925 ;
        RECT 203.155 122.215 203.485 122.545 ;
        RECT 203.155 120.165 203.485 120.495 ;
        RECT 203.155 118.235 203.485 118.565 ;
        RECT 203.155 116.395 203.485 116.725 ;
        RECT 203.155 114.905 203.485 115.235 ;
        RECT 203.155 113.235 203.485 113.565 ;
        RECT 203.155 111.745 203.485 112.075 ;
        RECT 203.155 110.075 203.485 110.405 ;
        RECT 203.155 108.585 203.485 108.915 ;
        RECT 203.155 106.915 203.485 107.245 ;
        RECT 203.155 105.425 203.485 105.755 ;
        RECT 203.155 104.015 203.485 104.345 ;
        RECT 203.155 102.175 203.485 102.505 ;
        RECT 203.155 100.685 203.485 101.015 ;
        RECT 203.155 99.015 203.485 99.345 ;
        RECT 203.155 97.525 203.485 97.855 ;
        RECT 203.155 95.855 203.485 96.185 ;
        RECT 203.155 94.365 203.485 94.695 ;
        RECT 203.155 92.695 203.485 93.025 ;
        RECT 203.155 91.205 203.485 91.535 ;
        RECT 203.155 89.795 203.485 90.125 ;
        RECT 203.155 87.955 203.485 88.285 ;
        RECT 203.155 86.465 203.485 86.795 ;
        RECT 203.155 84.795 203.485 85.125 ;
        RECT 203.155 83.305 203.485 83.635 ;
        RECT 203.155 81.635 203.485 81.965 ;
        RECT 203.155 80.145 203.485 80.475 ;
        RECT 203.155 78.475 203.485 78.805 ;
        RECT 203.155 76.985 203.485 77.315 ;
        RECT 203.155 75.575 203.485 75.905 ;
        RECT 203.155 73.735 203.485 74.065 ;
        RECT 203.155 72.245 203.485 72.575 ;
        RECT 203.155 70.575 203.485 70.905 ;
        RECT 203.155 69.085 203.485 69.415 ;
        RECT 203.155 67.415 203.485 67.745 ;
        RECT 203.155 65.925 203.485 66.255 ;
        RECT 203.155 64.255 203.485 64.585 ;
        RECT 203.155 62.765 203.485 63.095 ;
        RECT 203.155 61.355 203.485 61.685 ;
        RECT 203.155 59.515 203.485 59.845 ;
        RECT 203.155 58.025 203.485 58.355 ;
        RECT 203.155 56.355 203.485 56.685 ;
        RECT 203.155 54.865 203.485 55.195 ;
        RECT 203.155 53.195 203.485 53.525 ;
        RECT 203.155 51.705 203.485 52.035 ;
        RECT 203.155 50.035 203.485 50.365 ;
        RECT 203.155 48.545 203.485 48.875 ;
        RECT 203.155 47.135 203.485 47.465 ;
        RECT 203.155 45.295 203.485 45.625 ;
        RECT 203.155 43.805 203.485 44.135 ;
        RECT 203.155 42.135 203.485 42.465 ;
        RECT 203.155 40.645 203.485 40.975 ;
        RECT 203.155 38.975 203.485 39.305 ;
        RECT 203.155 37.485 203.485 37.815 ;
        RECT 203.155 35.815 203.485 36.145 ;
        RECT 203.155 34.325 203.485 34.655 ;
        RECT 203.155 32.915 203.485 33.245 ;
        RECT 203.155 31.075 203.485 31.405 ;
        RECT 203.155 29.585 203.485 29.915 ;
        RECT 203.155 27.915 203.485 28.245 ;
        RECT 203.155 26.425 203.485 26.755 ;
        RECT 203.155 24.755 203.485 25.085 ;
        RECT 203.155 23.265 203.485 23.595 ;
        RECT 203.155 21.595 203.485 21.925 ;
        RECT 203.155 20.105 203.485 20.435 ;
        RECT 203.155 18.695 203.485 19.025 ;
        RECT 203.155 16.855 203.485 17.185 ;
        RECT 203.155 15.365 203.485 15.695 ;
        RECT 203.155 13.695 203.485 14.025 ;
        RECT 203.155 12.205 203.485 12.535 ;
        RECT 203.155 10.535 203.485 10.865 ;
        RECT 203.155 9.045 203.485 9.375 ;
        RECT 203.155 7.375 203.485 7.705 ;
        RECT 203.155 5.885 203.485 6.215 ;
        RECT 203.155 4.475 203.485 4.805 ;
        RECT 203.155 2.115 203.485 2.445 ;
        RECT 203.155 0.06 203.485 0.39 ;
        RECT 203.155 -1.525 203.485 -1.195 ;
        RECT 203.155 -2.885 203.485 -2.555 ;
        RECT 203.155 -4.245 203.485 -3.915 ;
        RECT 203.155 -5.605 203.485 -5.275 ;
        RECT 203.155 -6.965 203.485 -6.635 ;
        RECT 203.155 -8.325 203.485 -7.995 ;
        RECT 203.155 -9.685 203.485 -9.355 ;
        RECT 203.155 -11.045 203.485 -10.715 ;
        RECT 203.155 -12.405 203.485 -12.075 ;
        RECT 203.155 -13.765 203.485 -13.435 ;
        RECT 203.155 -15.125 203.485 -14.795 ;
        RECT 203.155 -16.485 203.485 -16.155 ;
        RECT 203.155 -17.845 203.485 -17.515 ;
        RECT 203.155 -19.205 203.485 -18.875 ;
        RECT 203.155 -20.565 203.485 -20.235 ;
        RECT 203.155 -21.925 203.485 -21.595 ;
        RECT 203.155 -23.285 203.485 -22.955 ;
        RECT 203.155 -24.645 203.485 -24.315 ;
        RECT 203.155 -26.005 203.485 -25.675 ;
        RECT 203.155 -27.365 203.485 -27.035 ;
        RECT 203.155 -28.725 203.485 -28.395 ;
        RECT 203.155 -30.085 203.485 -29.755 ;
        RECT 203.155 -31.445 203.485 -31.115 ;
        RECT 203.155 -32.805 203.485 -32.475 ;
        RECT 203.155 -34.165 203.485 -33.835 ;
        RECT 203.155 -35.525 203.485 -35.195 ;
        RECT 203.155 -36.885 203.485 -36.555 ;
        RECT 203.155 -38.245 203.485 -37.915 ;
        RECT 203.155 -39.605 203.485 -39.275 ;
        RECT 203.155 -40.965 203.485 -40.635 ;
        RECT 203.155 -42.325 203.485 -41.995 ;
        RECT 203.155 -43.685 203.485 -43.355 ;
        RECT 203.155 -45.045 203.485 -44.715 ;
        RECT 203.155 -46.405 203.485 -46.075 ;
        RECT 203.155 -47.765 203.485 -47.435 ;
        RECT 203.155 -49.125 203.485 -48.795 ;
        RECT 203.155 -50.485 203.485 -50.155 ;
        RECT 203.155 -51.845 203.485 -51.515 ;
        RECT 203.155 -53.205 203.485 -52.875 ;
        RECT 203.155 -54.565 203.485 -54.235 ;
        RECT 203.155 -55.925 203.485 -55.595 ;
        RECT 203.155 -57.285 203.485 -56.955 ;
        RECT 203.155 -58.645 203.485 -58.315 ;
        RECT 203.155 -60.005 203.485 -59.675 ;
        RECT 203.155 -61.365 203.485 -61.035 ;
        RECT 203.155 -62.725 203.485 -62.395 ;
        RECT 203.155 -64.085 203.485 -63.755 ;
        RECT 203.155 -65.445 203.485 -65.115 ;
        RECT 203.155 -66.805 203.485 -66.475 ;
        RECT 203.155 -68.165 203.485 -67.835 ;
        RECT 203.155 -69.525 203.485 -69.195 ;
        RECT 203.155 -70.885 203.485 -70.555 ;
        RECT 203.155 -72.245 203.485 -71.915 ;
        RECT 203.155 -73.605 203.485 -73.275 ;
        RECT 203.155 -74.965 203.485 -74.635 ;
        RECT 203.155 -76.325 203.485 -75.995 ;
        RECT 203.155 -77.685 203.485 -77.355 ;
        RECT 203.155 -79.045 203.485 -78.715 ;
        RECT 203.155 -80.405 203.485 -80.075 ;
        RECT 203.155 -81.765 203.485 -81.435 ;
        RECT 203.155 -83.125 203.485 -82.795 ;
        RECT 203.155 -84.485 203.485 -84.155 ;
        RECT 203.155 -85.845 203.485 -85.515 ;
        RECT 203.155 -87.205 203.485 -86.875 ;
        RECT 203.155 -88.565 203.485 -88.235 ;
        RECT 203.155 -89.925 203.485 -89.595 ;
        RECT 203.155 -91.285 203.485 -90.955 ;
        RECT 203.155 -92.645 203.485 -92.315 ;
        RECT 203.155 -94.005 203.485 -93.675 ;
        RECT 203.155 -95.365 203.485 -95.035 ;
        RECT 203.155 -96.725 203.485 -96.395 ;
        RECT 203.155 -98.085 203.485 -97.755 ;
        RECT 203.155 -99.445 203.485 -99.115 ;
        RECT 203.155 -100.805 203.485 -100.475 ;
        RECT 203.155 -102.165 203.485 -101.835 ;
        RECT 203.155 -103.525 203.485 -103.195 ;
        RECT 203.155 -104.885 203.485 -104.555 ;
        RECT 203.155 -106.245 203.485 -105.915 ;
        RECT 203.155 -107.605 203.485 -107.275 ;
        RECT 203.155 -108.965 203.485 -108.635 ;
        RECT 203.155 -110.325 203.485 -109.995 ;
        RECT 203.155 -111.685 203.485 -111.355 ;
        RECT 203.155 -113.045 203.485 -112.715 ;
        RECT 203.155 -114.405 203.485 -114.075 ;
        RECT 203.155 -115.765 203.485 -115.435 ;
        RECT 203.155 -117.125 203.485 -116.795 ;
        RECT 203.155 -118.485 203.485 -118.155 ;
        RECT 203.155 -119.845 203.485 -119.515 ;
        RECT 203.155 -121.205 203.485 -120.875 ;
        RECT 203.155 -122.565 203.485 -122.235 ;
        RECT 203.155 -123.925 203.485 -123.595 ;
        RECT 203.155 -125.285 203.485 -124.955 ;
        RECT 203.155 -126.645 203.485 -126.315 ;
        RECT 203.155 -128.005 203.485 -127.675 ;
        RECT 203.155 -129.365 203.485 -129.035 ;
        RECT 203.155 -130.725 203.485 -130.395 ;
        RECT 203.155 -132.085 203.485 -131.755 ;
        RECT 203.155 -133.445 203.485 -133.115 ;
        RECT 203.155 -134.805 203.485 -134.475 ;
        RECT 203.155 -136.165 203.485 -135.835 ;
        RECT 203.155 -137.525 203.485 -137.195 ;
        RECT 203.155 -138.885 203.485 -138.555 ;
        RECT 203.155 -140.245 203.485 -139.915 ;
        RECT 203.155 -141.605 203.485 -141.275 ;
        RECT 203.155 -142.965 203.485 -142.635 ;
        RECT 203.155 -144.325 203.485 -143.995 ;
        RECT 203.155 -145.685 203.485 -145.355 ;
        RECT 203.155 -147.045 203.485 -146.715 ;
        RECT 203.155 -148.405 203.485 -148.075 ;
        RECT 203.155 -149.765 203.485 -149.435 ;
        RECT 203.155 -151.125 203.485 -150.795 ;
        RECT 203.155 -152.485 203.485 -152.155 ;
        RECT 203.155 -153.845 203.485 -153.515 ;
        RECT 203.155 -155.205 203.485 -154.875 ;
        RECT 203.155 -156.565 203.485 -156.235 ;
        RECT 203.155 -157.925 203.485 -157.595 ;
        RECT 203.155 -159.285 203.485 -158.955 ;
        RECT 203.155 -160.645 203.485 -160.315 ;
        RECT 203.155 -162.005 203.485 -161.675 ;
        RECT 203.155 -163.365 203.485 -163.035 ;
        RECT 203.155 -164.725 203.485 -164.395 ;
        RECT 203.155 -166.085 203.485 -165.755 ;
        RECT 203.155 -167.445 203.485 -167.115 ;
        RECT 203.155 -168.805 203.485 -168.475 ;
        RECT 203.155 -170.165 203.485 -169.835 ;
        RECT 203.155 -171.525 203.485 -171.195 ;
        RECT 203.155 -172.885 203.485 -172.555 ;
        RECT 203.155 -174.245 203.485 -173.915 ;
        RECT 203.155 -175.605 203.485 -175.275 ;
        RECT 203.155 -176.965 203.485 -176.635 ;
        RECT 203.155 -178.325 203.485 -177.995 ;
        RECT 203.155 -179.685 203.485 -179.355 ;
        RECT 203.155 -181.045 203.485 -180.715 ;
        RECT 203.155 -182.405 203.485 -182.075 ;
        RECT 203.155 -183.765 203.485 -183.435 ;
        RECT 203.155 -185.125 203.485 -184.795 ;
        RECT 203.155 -186.485 203.485 -186.155 ;
        RECT 203.155 -187.845 203.485 -187.515 ;
        RECT 203.155 -189.205 203.485 -188.875 ;
        RECT 203.155 -190.565 203.485 -190.235 ;
        RECT 203.155 -191.925 203.485 -191.595 ;
        RECT 203.155 -193.285 203.485 -192.955 ;
        RECT 203.155 -194.645 203.485 -194.315 ;
        RECT 203.155 -196.005 203.485 -195.675 ;
        RECT 203.155 -197.365 203.485 -197.035 ;
        RECT 203.155 -198.725 203.485 -198.395 ;
        RECT 203.155 -200.085 203.485 -199.755 ;
        RECT 203.155 -201.445 203.485 -201.115 ;
        RECT 203.155 -202.805 203.485 -202.475 ;
        RECT 203.155 -204.165 203.485 -203.835 ;
        RECT 203.155 -205.525 203.485 -205.195 ;
        RECT 203.155 -206.885 203.485 -206.555 ;
        RECT 203.155 -208.245 203.485 -207.915 ;
        RECT 203.155 -209.605 203.485 -209.275 ;
        RECT 203.155 -210.965 203.485 -210.635 ;
        RECT 203.155 -212.325 203.485 -211.995 ;
        RECT 203.155 -213.685 203.485 -213.355 ;
        RECT 203.155 -215.045 203.485 -214.715 ;
        RECT 203.155 -216.405 203.485 -216.075 ;
        RECT 203.155 -217.765 203.485 -217.435 ;
        RECT 203.155 -219.125 203.485 -218.795 ;
        RECT 203.155 -221.37 203.485 -220.24 ;
        RECT 203.16 -221.485 203.48 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.515 18.695 204.845 19.025 ;
        RECT 204.515 16.855 204.845 17.185 ;
        RECT 204.515 15.365 204.845 15.695 ;
        RECT 204.515 13.695 204.845 14.025 ;
        RECT 204.515 12.205 204.845 12.535 ;
        RECT 204.515 10.535 204.845 10.865 ;
        RECT 204.515 9.045 204.845 9.375 ;
        RECT 204.515 7.375 204.845 7.705 ;
        RECT 204.515 5.885 204.845 6.215 ;
        RECT 204.515 4.475 204.845 4.805 ;
        RECT 204.515 2.115 204.845 2.445 ;
        RECT 204.515 0.06 204.845 0.39 ;
        RECT 204.515 -1.525 204.845 -1.195 ;
        RECT 204.515 -2.885 204.845 -2.555 ;
        RECT 204.515 -4.245 204.845 -3.915 ;
        RECT 204.515 -5.605 204.845 -5.275 ;
        RECT 204.515 -6.965 204.845 -6.635 ;
        RECT 204.515 -8.325 204.845 -7.995 ;
        RECT 204.515 -9.685 204.845 -9.355 ;
        RECT 204.515 -11.045 204.845 -10.715 ;
        RECT 204.515 -12.405 204.845 -12.075 ;
        RECT 204.515 -13.765 204.845 -13.435 ;
        RECT 204.515 -15.125 204.845 -14.795 ;
        RECT 204.515 -16.485 204.845 -16.155 ;
        RECT 204.515 -17.845 204.845 -17.515 ;
        RECT 204.515 -19.205 204.845 -18.875 ;
        RECT 204.515 -20.565 204.845 -20.235 ;
        RECT 204.515 -21.925 204.845 -21.595 ;
        RECT 204.515 -23.285 204.845 -22.955 ;
        RECT 204.515 -24.645 204.845 -24.315 ;
        RECT 204.515 -26.005 204.845 -25.675 ;
        RECT 204.515 -27.365 204.845 -27.035 ;
        RECT 204.515 -28.725 204.845 -28.395 ;
        RECT 204.515 -30.085 204.845 -29.755 ;
        RECT 204.515 -31.445 204.845 -31.115 ;
        RECT 204.515 -32.805 204.845 -32.475 ;
        RECT 204.515 -34.165 204.845 -33.835 ;
        RECT 204.515 -35.525 204.845 -35.195 ;
        RECT 204.515 -36.885 204.845 -36.555 ;
        RECT 204.515 -38.245 204.845 -37.915 ;
        RECT 204.515 -39.605 204.845 -39.275 ;
        RECT 204.515 -40.965 204.845 -40.635 ;
        RECT 204.515 -42.325 204.845 -41.995 ;
        RECT 204.515 -43.685 204.845 -43.355 ;
        RECT 204.515 -45.045 204.845 -44.715 ;
        RECT 204.515 -46.405 204.845 -46.075 ;
        RECT 204.515 -47.765 204.845 -47.435 ;
        RECT 204.515 -49.125 204.845 -48.795 ;
        RECT 204.515 -50.485 204.845 -50.155 ;
        RECT 204.515 -51.845 204.845 -51.515 ;
        RECT 204.515 -53.205 204.845 -52.875 ;
        RECT 204.515 -54.565 204.845 -54.235 ;
        RECT 204.515 -55.925 204.845 -55.595 ;
        RECT 204.515 -57.285 204.845 -56.955 ;
        RECT 204.515 -58.645 204.845 -58.315 ;
        RECT 204.515 -60.005 204.845 -59.675 ;
        RECT 204.515 -61.365 204.845 -61.035 ;
        RECT 204.515 -62.725 204.845 -62.395 ;
        RECT 204.515 -64.085 204.845 -63.755 ;
        RECT 204.515 -65.445 204.845 -65.115 ;
        RECT 204.515 -66.805 204.845 -66.475 ;
        RECT 204.515 -68.165 204.845 -67.835 ;
        RECT 204.515 -69.525 204.845 -69.195 ;
        RECT 204.515 -70.885 204.845 -70.555 ;
        RECT 204.515 -72.245 204.845 -71.915 ;
        RECT 204.515 -73.605 204.845 -73.275 ;
        RECT 204.515 -74.965 204.845 -74.635 ;
        RECT 204.515 -76.325 204.845 -75.995 ;
        RECT 204.515 -77.685 204.845 -77.355 ;
        RECT 204.515 -79.045 204.845 -78.715 ;
        RECT 204.515 -80.405 204.845 -80.075 ;
        RECT 204.515 -81.765 204.845 -81.435 ;
        RECT 204.515 -83.125 204.845 -82.795 ;
        RECT 204.515 -84.485 204.845 -84.155 ;
        RECT 204.515 -85.845 204.845 -85.515 ;
        RECT 204.515 -87.205 204.845 -86.875 ;
        RECT 204.515 -88.565 204.845 -88.235 ;
        RECT 204.515 -89.925 204.845 -89.595 ;
        RECT 204.515 -91.285 204.845 -90.955 ;
        RECT 204.515 -92.645 204.845 -92.315 ;
        RECT 204.515 -94.005 204.845 -93.675 ;
        RECT 204.515 -95.365 204.845 -95.035 ;
        RECT 204.515 -96.725 204.845 -96.395 ;
        RECT 204.515 -98.085 204.845 -97.755 ;
        RECT 204.515 -99.445 204.845 -99.115 ;
        RECT 204.515 -100.805 204.845 -100.475 ;
        RECT 204.515 -102.165 204.845 -101.835 ;
        RECT 204.515 -103.525 204.845 -103.195 ;
        RECT 204.515 -104.885 204.845 -104.555 ;
        RECT 204.515 -106.245 204.845 -105.915 ;
        RECT 204.515 -107.605 204.845 -107.275 ;
        RECT 204.515 -108.965 204.845 -108.635 ;
        RECT 204.515 -110.325 204.845 -109.995 ;
        RECT 204.515 -111.685 204.845 -111.355 ;
        RECT 204.515 -113.045 204.845 -112.715 ;
        RECT 204.515 -114.405 204.845 -114.075 ;
        RECT 204.515 -115.765 204.845 -115.435 ;
        RECT 204.515 -117.125 204.845 -116.795 ;
        RECT 204.515 -118.485 204.845 -118.155 ;
        RECT 204.515 -119.845 204.845 -119.515 ;
        RECT 204.515 -121.205 204.845 -120.875 ;
        RECT 204.515 -122.565 204.845 -122.235 ;
        RECT 204.515 -123.925 204.845 -123.595 ;
        RECT 204.515 -125.285 204.845 -124.955 ;
        RECT 204.515 -126.645 204.845 -126.315 ;
        RECT 204.515 -128.005 204.845 -127.675 ;
        RECT 204.515 -129.365 204.845 -129.035 ;
        RECT 204.515 -130.725 204.845 -130.395 ;
        RECT 204.515 -132.085 204.845 -131.755 ;
        RECT 204.515 -133.445 204.845 -133.115 ;
        RECT 204.515 -134.805 204.845 -134.475 ;
        RECT 204.515 -136.165 204.845 -135.835 ;
        RECT 204.515 -137.525 204.845 -137.195 ;
        RECT 204.515 -138.885 204.845 -138.555 ;
        RECT 204.515 -140.245 204.845 -139.915 ;
        RECT 204.515 -141.605 204.845 -141.275 ;
        RECT 204.515 -142.965 204.845 -142.635 ;
        RECT 204.515 -144.325 204.845 -143.995 ;
        RECT 204.515 -145.685 204.845 -145.355 ;
        RECT 204.515 -147.045 204.845 -146.715 ;
        RECT 204.515 -148.405 204.845 -148.075 ;
        RECT 204.515 -149.765 204.845 -149.435 ;
        RECT 204.515 -151.125 204.845 -150.795 ;
        RECT 204.515 -152.485 204.845 -152.155 ;
        RECT 204.515 -153.845 204.845 -153.515 ;
        RECT 204.515 -155.205 204.845 -154.875 ;
        RECT 204.515 -156.565 204.845 -156.235 ;
        RECT 204.515 -157.925 204.845 -157.595 ;
        RECT 204.515 -159.285 204.845 -158.955 ;
        RECT 204.515 -160.645 204.845 -160.315 ;
        RECT 204.515 -162.005 204.845 -161.675 ;
        RECT 204.515 -163.365 204.845 -163.035 ;
        RECT 204.515 -164.725 204.845 -164.395 ;
        RECT 204.515 -166.085 204.845 -165.755 ;
        RECT 204.515 -167.445 204.845 -167.115 ;
        RECT 204.515 -168.805 204.845 -168.475 ;
        RECT 204.515 -170.165 204.845 -169.835 ;
        RECT 204.515 -171.525 204.845 -171.195 ;
        RECT 204.515 -172.885 204.845 -172.555 ;
        RECT 204.515 -174.245 204.845 -173.915 ;
        RECT 204.515 -175.605 204.845 -175.275 ;
        RECT 204.515 -176.965 204.845 -176.635 ;
        RECT 204.515 -178.325 204.845 -177.995 ;
        RECT 204.515 -179.685 204.845 -179.355 ;
        RECT 204.515 -181.045 204.845 -180.715 ;
        RECT 204.515 -182.405 204.845 -182.075 ;
        RECT 204.515 -183.765 204.845 -183.435 ;
        RECT 204.515 -185.125 204.845 -184.795 ;
        RECT 204.515 -186.485 204.845 -186.155 ;
        RECT 204.515 -187.845 204.845 -187.515 ;
        RECT 204.515 -189.205 204.845 -188.875 ;
        RECT 204.515 -190.565 204.845 -190.235 ;
        RECT 204.515 -191.925 204.845 -191.595 ;
        RECT 204.515 -193.285 204.845 -192.955 ;
        RECT 204.515 -194.645 204.845 -194.315 ;
        RECT 204.515 -196.005 204.845 -195.675 ;
        RECT 204.515 -197.365 204.845 -197.035 ;
        RECT 204.515 -198.725 204.845 -198.395 ;
        RECT 204.515 -200.085 204.845 -199.755 ;
        RECT 204.515 -201.445 204.845 -201.115 ;
        RECT 204.515 -202.805 204.845 -202.475 ;
        RECT 204.515 -204.165 204.845 -203.835 ;
        RECT 204.515 -205.525 204.845 -205.195 ;
        RECT 204.515 -206.885 204.845 -206.555 ;
        RECT 204.515 -208.245 204.845 -207.915 ;
        RECT 204.515 -209.605 204.845 -209.275 ;
        RECT 204.515 -210.965 204.845 -210.635 ;
        RECT 204.515 -212.325 204.845 -211.995 ;
        RECT 204.515 -213.685 204.845 -213.355 ;
        RECT 204.515 -215.045 204.845 -214.715 ;
        RECT 204.515 -216.405 204.845 -216.075 ;
        RECT 204.515 -217.765 204.845 -217.435 ;
        RECT 204.515 -219.125 204.845 -218.795 ;
        RECT 204.515 -221.37 204.845 -220.24 ;
        RECT 204.52 -221.485 204.84 131.045 ;
        RECT 204.515 129.8 204.845 130.93 ;
        RECT 204.515 127.675 204.845 128.005 ;
        RECT 204.515 126.315 204.845 126.645 ;
        RECT 204.515 124.955 204.845 125.285 ;
        RECT 204.515 123.595 204.845 123.925 ;
        RECT 204.515 122.215 204.845 122.545 ;
        RECT 204.515 120.165 204.845 120.495 ;
        RECT 204.515 118.235 204.845 118.565 ;
        RECT 204.515 116.395 204.845 116.725 ;
        RECT 204.515 114.905 204.845 115.235 ;
        RECT 204.515 113.235 204.845 113.565 ;
        RECT 204.515 111.745 204.845 112.075 ;
        RECT 204.515 110.075 204.845 110.405 ;
        RECT 204.515 108.585 204.845 108.915 ;
        RECT 204.515 106.915 204.845 107.245 ;
        RECT 204.515 105.425 204.845 105.755 ;
        RECT 204.515 104.015 204.845 104.345 ;
        RECT 204.515 102.175 204.845 102.505 ;
        RECT 204.515 100.685 204.845 101.015 ;
        RECT 204.515 99.015 204.845 99.345 ;
        RECT 204.515 97.525 204.845 97.855 ;
        RECT 204.515 95.855 204.845 96.185 ;
        RECT 204.515 94.365 204.845 94.695 ;
        RECT 204.515 92.695 204.845 93.025 ;
        RECT 204.515 91.205 204.845 91.535 ;
        RECT 204.515 89.795 204.845 90.125 ;
        RECT 204.515 87.955 204.845 88.285 ;
        RECT 204.515 86.465 204.845 86.795 ;
        RECT 204.515 84.795 204.845 85.125 ;
        RECT 204.515 83.305 204.845 83.635 ;
        RECT 204.515 81.635 204.845 81.965 ;
        RECT 204.515 80.145 204.845 80.475 ;
        RECT 204.515 78.475 204.845 78.805 ;
        RECT 204.515 76.985 204.845 77.315 ;
        RECT 204.515 75.575 204.845 75.905 ;
        RECT 204.515 73.735 204.845 74.065 ;
        RECT 204.515 72.245 204.845 72.575 ;
        RECT 204.515 70.575 204.845 70.905 ;
        RECT 204.515 69.085 204.845 69.415 ;
        RECT 204.515 67.415 204.845 67.745 ;
        RECT 204.515 65.925 204.845 66.255 ;
        RECT 204.515 64.255 204.845 64.585 ;
        RECT 204.515 62.765 204.845 63.095 ;
        RECT 204.515 61.355 204.845 61.685 ;
        RECT 204.515 59.515 204.845 59.845 ;
        RECT 204.515 58.025 204.845 58.355 ;
        RECT 204.515 56.355 204.845 56.685 ;
        RECT 204.515 54.865 204.845 55.195 ;
        RECT 204.515 53.195 204.845 53.525 ;
        RECT 204.515 51.705 204.845 52.035 ;
        RECT 204.515 50.035 204.845 50.365 ;
        RECT 204.515 48.545 204.845 48.875 ;
        RECT 204.515 47.135 204.845 47.465 ;
        RECT 204.515 45.295 204.845 45.625 ;
        RECT 204.515 43.805 204.845 44.135 ;
        RECT 204.515 42.135 204.845 42.465 ;
        RECT 204.515 40.645 204.845 40.975 ;
        RECT 204.515 38.975 204.845 39.305 ;
        RECT 204.515 37.485 204.845 37.815 ;
        RECT 204.515 35.815 204.845 36.145 ;
        RECT 204.515 34.325 204.845 34.655 ;
        RECT 204.515 32.915 204.845 33.245 ;
        RECT 204.515 31.075 204.845 31.405 ;
        RECT 204.515 29.585 204.845 29.915 ;
        RECT 204.515 27.915 204.845 28.245 ;
        RECT 204.515 26.425 204.845 26.755 ;
        RECT 204.515 24.755 204.845 25.085 ;
        RECT 204.515 23.265 204.845 23.595 ;
        RECT 204.515 21.595 204.845 21.925 ;
        RECT 204.515 20.105 204.845 20.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.435 129.8 166.765 130.93 ;
        RECT 166.435 127.675 166.765 128.005 ;
        RECT 166.435 126.315 166.765 126.645 ;
        RECT 166.435 124.955 166.765 125.285 ;
        RECT 166.435 123.595 166.765 123.925 ;
        RECT 166.44 123.595 166.76 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.435 -1.525 166.765 -1.195 ;
        RECT 166.435 -2.885 166.765 -2.555 ;
        RECT 166.44 -3.56 166.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.435 -118.485 166.765 -118.155 ;
        RECT 166.435 -119.845 166.765 -119.515 ;
        RECT 166.435 -121.205 166.765 -120.875 ;
        RECT 166.435 -122.565 166.765 -122.235 ;
        RECT 166.435 -123.925 166.765 -123.595 ;
        RECT 166.435 -125.285 166.765 -124.955 ;
        RECT 166.435 -126.645 166.765 -126.315 ;
        RECT 166.435 -128.005 166.765 -127.675 ;
        RECT 166.435 -129.365 166.765 -129.035 ;
        RECT 166.435 -130.725 166.765 -130.395 ;
        RECT 166.435 -132.085 166.765 -131.755 ;
        RECT 166.435 -133.445 166.765 -133.115 ;
        RECT 166.435 -134.805 166.765 -134.475 ;
        RECT 166.435 -136.165 166.765 -135.835 ;
        RECT 166.435 -137.525 166.765 -137.195 ;
        RECT 166.435 -138.885 166.765 -138.555 ;
        RECT 166.435 -140.245 166.765 -139.915 ;
        RECT 166.435 -141.605 166.765 -141.275 ;
        RECT 166.435 -142.965 166.765 -142.635 ;
        RECT 166.435 -144.325 166.765 -143.995 ;
        RECT 166.435 -145.685 166.765 -145.355 ;
        RECT 166.435 -147.045 166.765 -146.715 ;
        RECT 166.435 -148.405 166.765 -148.075 ;
        RECT 166.435 -149.765 166.765 -149.435 ;
        RECT 166.435 -151.125 166.765 -150.795 ;
        RECT 166.435 -152.485 166.765 -152.155 ;
        RECT 166.435 -153.845 166.765 -153.515 ;
        RECT 166.435 -155.205 166.765 -154.875 ;
        RECT 166.435 -156.565 166.765 -156.235 ;
        RECT 166.435 -157.925 166.765 -157.595 ;
        RECT 166.435 -159.285 166.765 -158.955 ;
        RECT 166.435 -160.645 166.765 -160.315 ;
        RECT 166.435 -162.005 166.765 -161.675 ;
        RECT 166.435 -163.365 166.765 -163.035 ;
        RECT 166.435 -164.725 166.765 -164.395 ;
        RECT 166.435 -166.085 166.765 -165.755 ;
        RECT 166.435 -167.445 166.765 -167.115 ;
        RECT 166.435 -168.805 166.765 -168.475 ;
        RECT 166.435 -170.165 166.765 -169.835 ;
        RECT 166.435 -171.525 166.765 -171.195 ;
        RECT 166.435 -172.885 166.765 -172.555 ;
        RECT 166.435 -174.245 166.765 -173.915 ;
        RECT 166.435 -175.605 166.765 -175.275 ;
        RECT 166.435 -176.965 166.765 -176.635 ;
        RECT 166.435 -178.325 166.765 -177.995 ;
        RECT 166.435 -179.685 166.765 -179.355 ;
        RECT 166.435 -181.045 166.765 -180.715 ;
        RECT 166.435 -182.405 166.765 -182.075 ;
        RECT 166.435 -183.765 166.765 -183.435 ;
        RECT 166.435 -185.125 166.765 -184.795 ;
        RECT 166.435 -186.485 166.765 -186.155 ;
        RECT 166.435 -187.845 166.765 -187.515 ;
        RECT 166.435 -189.205 166.765 -188.875 ;
        RECT 166.435 -190.565 166.765 -190.235 ;
        RECT 166.435 -191.925 166.765 -191.595 ;
        RECT 166.435 -193.285 166.765 -192.955 ;
        RECT 166.435 -194.645 166.765 -194.315 ;
        RECT 166.435 -196.005 166.765 -195.675 ;
        RECT 166.435 -197.365 166.765 -197.035 ;
        RECT 166.435 -198.725 166.765 -198.395 ;
        RECT 166.435 -200.085 166.765 -199.755 ;
        RECT 166.435 -201.445 166.765 -201.115 ;
        RECT 166.435 -202.805 166.765 -202.475 ;
        RECT 166.435 -204.165 166.765 -203.835 ;
        RECT 166.435 -205.525 166.765 -205.195 ;
        RECT 166.435 -206.885 166.765 -206.555 ;
        RECT 166.435 -208.245 166.765 -207.915 ;
        RECT 166.435 -209.605 166.765 -209.275 ;
        RECT 166.435 -210.965 166.765 -210.635 ;
        RECT 166.435 -212.325 166.765 -211.995 ;
        RECT 166.435 -213.685 166.765 -213.355 ;
        RECT 166.435 -215.045 166.765 -214.715 ;
        RECT 166.435 -216.405 166.765 -216.075 ;
        RECT 166.435 -217.765 166.765 -217.435 ;
        RECT 166.435 -219.125 166.765 -218.795 ;
        RECT 166.435 -221.37 166.765 -220.24 ;
        RECT 166.44 -221.485 166.76 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.795 129.8 168.125 130.93 ;
        RECT 167.795 127.675 168.125 128.005 ;
        RECT 167.795 126.315 168.125 126.645 ;
        RECT 167.795 124.955 168.125 125.285 ;
        RECT 167.795 123.595 168.125 123.925 ;
        RECT 167.8 123.595 168.12 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.795 -122.565 168.125 -122.235 ;
        RECT 167.795 -123.925 168.125 -123.595 ;
        RECT 167.795 -125.285 168.125 -124.955 ;
        RECT 167.795 -126.645 168.125 -126.315 ;
        RECT 167.795 -128.005 168.125 -127.675 ;
        RECT 167.795 -129.365 168.125 -129.035 ;
        RECT 167.795 -130.725 168.125 -130.395 ;
        RECT 167.795 -132.085 168.125 -131.755 ;
        RECT 167.795 -133.445 168.125 -133.115 ;
        RECT 167.795 -134.805 168.125 -134.475 ;
        RECT 167.795 -136.165 168.125 -135.835 ;
        RECT 167.795 -137.525 168.125 -137.195 ;
        RECT 167.795 -138.885 168.125 -138.555 ;
        RECT 167.795 -140.245 168.125 -139.915 ;
        RECT 167.795 -141.605 168.125 -141.275 ;
        RECT 167.795 -142.965 168.125 -142.635 ;
        RECT 167.795 -144.325 168.125 -143.995 ;
        RECT 167.795 -145.685 168.125 -145.355 ;
        RECT 167.795 -147.045 168.125 -146.715 ;
        RECT 167.795 -148.405 168.125 -148.075 ;
        RECT 167.795 -149.765 168.125 -149.435 ;
        RECT 167.795 -151.125 168.125 -150.795 ;
        RECT 167.795 -152.485 168.125 -152.155 ;
        RECT 167.795 -153.845 168.125 -153.515 ;
        RECT 167.795 -155.205 168.125 -154.875 ;
        RECT 167.795 -156.565 168.125 -156.235 ;
        RECT 167.795 -157.925 168.125 -157.595 ;
        RECT 167.795 -159.285 168.125 -158.955 ;
        RECT 167.795 -160.645 168.125 -160.315 ;
        RECT 167.795 -162.005 168.125 -161.675 ;
        RECT 167.795 -163.365 168.125 -163.035 ;
        RECT 167.795 -164.725 168.125 -164.395 ;
        RECT 167.795 -166.085 168.125 -165.755 ;
        RECT 167.795 -167.445 168.125 -167.115 ;
        RECT 167.795 -168.805 168.125 -168.475 ;
        RECT 167.795 -170.165 168.125 -169.835 ;
        RECT 167.795 -171.525 168.125 -171.195 ;
        RECT 167.795 -172.885 168.125 -172.555 ;
        RECT 167.795 -174.245 168.125 -173.915 ;
        RECT 167.795 -175.605 168.125 -175.275 ;
        RECT 167.795 -176.965 168.125 -176.635 ;
        RECT 167.795 -178.325 168.125 -177.995 ;
        RECT 167.795 -179.685 168.125 -179.355 ;
        RECT 167.795 -181.045 168.125 -180.715 ;
        RECT 167.795 -182.405 168.125 -182.075 ;
        RECT 167.795 -183.765 168.125 -183.435 ;
        RECT 167.795 -185.125 168.125 -184.795 ;
        RECT 167.795 -186.485 168.125 -186.155 ;
        RECT 167.795 -187.845 168.125 -187.515 ;
        RECT 167.795 -189.205 168.125 -188.875 ;
        RECT 167.795 -190.565 168.125 -190.235 ;
        RECT 167.795 -191.925 168.125 -191.595 ;
        RECT 167.795 -193.285 168.125 -192.955 ;
        RECT 167.795 -194.645 168.125 -194.315 ;
        RECT 167.795 -196.005 168.125 -195.675 ;
        RECT 167.795 -197.365 168.125 -197.035 ;
        RECT 167.795 -198.725 168.125 -198.395 ;
        RECT 167.795 -200.085 168.125 -199.755 ;
        RECT 167.795 -201.445 168.125 -201.115 ;
        RECT 167.795 -202.805 168.125 -202.475 ;
        RECT 167.795 -204.165 168.125 -203.835 ;
        RECT 167.795 -205.525 168.125 -205.195 ;
        RECT 167.795 -206.885 168.125 -206.555 ;
        RECT 167.795 -208.245 168.125 -207.915 ;
        RECT 167.795 -209.605 168.125 -209.275 ;
        RECT 167.795 -210.965 168.125 -210.635 ;
        RECT 167.795 -212.325 168.125 -211.995 ;
        RECT 167.795 -213.685 168.125 -213.355 ;
        RECT 167.795 -215.045 168.125 -214.715 ;
        RECT 167.795 -216.405 168.125 -216.075 ;
        RECT 167.795 -217.765 168.125 -217.435 ;
        RECT 167.795 -219.125 168.125 -218.795 ;
        RECT 167.795 -221.37 168.125 -220.24 ;
        RECT 167.8 -221.485 168.12 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.01 -121.535 168.34 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.155 129.8 169.485 130.93 ;
        RECT 169.155 127.675 169.485 128.005 ;
        RECT 169.155 126.315 169.485 126.645 ;
        RECT 169.155 124.955 169.485 125.285 ;
        RECT 169.155 123.595 169.485 123.925 ;
        RECT 169.16 123.595 169.48 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.155 -1.525 169.485 -1.195 ;
        RECT 169.155 -2.885 169.485 -2.555 ;
        RECT 169.16 -3.56 169.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.515 129.8 170.845 130.93 ;
        RECT 170.515 127.675 170.845 128.005 ;
        RECT 170.515 126.315 170.845 126.645 ;
        RECT 170.515 124.955 170.845 125.285 ;
        RECT 170.515 123.595 170.845 123.925 ;
        RECT 170.52 123.595 170.84 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.515 -1.525 170.845 -1.195 ;
        RECT 170.515 -2.885 170.845 -2.555 ;
        RECT 170.52 -3.56 170.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.875 129.8 172.205 130.93 ;
        RECT 171.875 127.675 172.205 128.005 ;
        RECT 171.875 126.315 172.205 126.645 ;
        RECT 171.875 124.955 172.205 125.285 ;
        RECT 171.875 123.595 172.205 123.925 ;
        RECT 171.88 123.595 172.2 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.875 -1.525 172.205 -1.195 ;
        RECT 171.875 -2.885 172.205 -2.555 ;
        RECT 171.88 -3.56 172.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.875 -118.485 172.205 -118.155 ;
        RECT 171.875 -119.845 172.205 -119.515 ;
        RECT 171.875 -121.205 172.205 -120.875 ;
        RECT 171.875 -122.565 172.205 -122.235 ;
        RECT 171.875 -123.925 172.205 -123.595 ;
        RECT 171.875 -125.285 172.205 -124.955 ;
        RECT 171.875 -126.645 172.205 -126.315 ;
        RECT 171.875 -128.005 172.205 -127.675 ;
        RECT 171.875 -129.365 172.205 -129.035 ;
        RECT 171.875 -130.725 172.205 -130.395 ;
        RECT 171.875 -132.085 172.205 -131.755 ;
        RECT 171.875 -133.445 172.205 -133.115 ;
        RECT 171.875 -134.805 172.205 -134.475 ;
        RECT 171.875 -136.165 172.205 -135.835 ;
        RECT 171.875 -137.525 172.205 -137.195 ;
        RECT 171.875 -138.885 172.205 -138.555 ;
        RECT 171.875 -140.245 172.205 -139.915 ;
        RECT 171.875 -141.605 172.205 -141.275 ;
        RECT 171.875 -142.965 172.205 -142.635 ;
        RECT 171.875 -144.325 172.205 -143.995 ;
        RECT 171.875 -145.685 172.205 -145.355 ;
        RECT 171.875 -147.045 172.205 -146.715 ;
        RECT 171.875 -148.405 172.205 -148.075 ;
        RECT 171.875 -149.765 172.205 -149.435 ;
        RECT 171.875 -151.125 172.205 -150.795 ;
        RECT 171.875 -152.485 172.205 -152.155 ;
        RECT 171.875 -153.845 172.205 -153.515 ;
        RECT 171.875 -155.205 172.205 -154.875 ;
        RECT 171.875 -156.565 172.205 -156.235 ;
        RECT 171.875 -157.925 172.205 -157.595 ;
        RECT 171.875 -159.285 172.205 -158.955 ;
        RECT 171.875 -160.645 172.205 -160.315 ;
        RECT 171.875 -162.005 172.205 -161.675 ;
        RECT 171.875 -163.365 172.205 -163.035 ;
        RECT 171.875 -164.725 172.205 -164.395 ;
        RECT 171.875 -166.085 172.205 -165.755 ;
        RECT 171.875 -167.445 172.205 -167.115 ;
        RECT 171.875 -168.805 172.205 -168.475 ;
        RECT 171.875 -170.165 172.205 -169.835 ;
        RECT 171.875 -171.525 172.205 -171.195 ;
        RECT 171.875 -172.885 172.205 -172.555 ;
        RECT 171.875 -174.245 172.205 -173.915 ;
        RECT 171.875 -175.605 172.205 -175.275 ;
        RECT 171.875 -176.965 172.205 -176.635 ;
        RECT 171.875 -178.325 172.205 -177.995 ;
        RECT 171.875 -179.685 172.205 -179.355 ;
        RECT 171.875 -181.045 172.205 -180.715 ;
        RECT 171.875 -182.405 172.205 -182.075 ;
        RECT 171.875 -183.765 172.205 -183.435 ;
        RECT 171.875 -185.125 172.205 -184.795 ;
        RECT 171.875 -186.485 172.205 -186.155 ;
        RECT 171.875 -187.845 172.205 -187.515 ;
        RECT 171.875 -189.205 172.205 -188.875 ;
        RECT 171.875 -190.565 172.205 -190.235 ;
        RECT 171.875 -191.925 172.205 -191.595 ;
        RECT 171.875 -193.285 172.205 -192.955 ;
        RECT 171.875 -194.645 172.205 -194.315 ;
        RECT 171.875 -196.005 172.205 -195.675 ;
        RECT 171.875 -197.365 172.205 -197.035 ;
        RECT 171.875 -198.725 172.205 -198.395 ;
        RECT 171.875 -200.085 172.205 -199.755 ;
        RECT 171.875 -201.445 172.205 -201.115 ;
        RECT 171.875 -202.805 172.205 -202.475 ;
        RECT 171.875 -204.165 172.205 -203.835 ;
        RECT 171.875 -205.525 172.205 -205.195 ;
        RECT 171.875 -206.885 172.205 -206.555 ;
        RECT 171.875 -208.245 172.205 -207.915 ;
        RECT 171.875 -209.605 172.205 -209.275 ;
        RECT 171.875 -210.965 172.205 -210.635 ;
        RECT 171.875 -212.325 172.205 -211.995 ;
        RECT 171.875 -213.685 172.205 -213.355 ;
        RECT 171.875 -215.045 172.205 -214.715 ;
        RECT 171.875 -216.405 172.205 -216.075 ;
        RECT 171.875 -217.765 172.205 -217.435 ;
        RECT 171.875 -219.125 172.205 -218.795 ;
        RECT 171.875 -221.37 172.205 -220.24 ;
        RECT 171.88 -221.485 172.2 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.235 129.8 173.565 130.93 ;
        RECT 173.235 127.675 173.565 128.005 ;
        RECT 173.235 126.315 173.565 126.645 ;
        RECT 173.235 124.955 173.565 125.285 ;
        RECT 173.235 123.595 173.565 123.925 ;
        RECT 173.24 123.595 173.56 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.235 -122.565 173.565 -122.235 ;
        RECT 173.235 -123.925 173.565 -123.595 ;
        RECT 173.235 -125.285 173.565 -124.955 ;
        RECT 173.235 -126.645 173.565 -126.315 ;
        RECT 173.235 -128.005 173.565 -127.675 ;
        RECT 173.235 -129.365 173.565 -129.035 ;
        RECT 173.235 -130.725 173.565 -130.395 ;
        RECT 173.235 -132.085 173.565 -131.755 ;
        RECT 173.235 -133.445 173.565 -133.115 ;
        RECT 173.235 -134.805 173.565 -134.475 ;
        RECT 173.235 -136.165 173.565 -135.835 ;
        RECT 173.235 -137.525 173.565 -137.195 ;
        RECT 173.235 -138.885 173.565 -138.555 ;
        RECT 173.235 -140.245 173.565 -139.915 ;
        RECT 173.235 -141.605 173.565 -141.275 ;
        RECT 173.235 -142.965 173.565 -142.635 ;
        RECT 173.235 -144.325 173.565 -143.995 ;
        RECT 173.235 -145.685 173.565 -145.355 ;
        RECT 173.235 -147.045 173.565 -146.715 ;
        RECT 173.235 -148.405 173.565 -148.075 ;
        RECT 173.235 -149.765 173.565 -149.435 ;
        RECT 173.235 -151.125 173.565 -150.795 ;
        RECT 173.235 -152.485 173.565 -152.155 ;
        RECT 173.235 -153.845 173.565 -153.515 ;
        RECT 173.235 -155.205 173.565 -154.875 ;
        RECT 173.235 -156.565 173.565 -156.235 ;
        RECT 173.235 -157.925 173.565 -157.595 ;
        RECT 173.235 -159.285 173.565 -158.955 ;
        RECT 173.235 -160.645 173.565 -160.315 ;
        RECT 173.235 -162.005 173.565 -161.675 ;
        RECT 173.235 -163.365 173.565 -163.035 ;
        RECT 173.235 -164.725 173.565 -164.395 ;
        RECT 173.235 -166.085 173.565 -165.755 ;
        RECT 173.235 -167.445 173.565 -167.115 ;
        RECT 173.235 -168.805 173.565 -168.475 ;
        RECT 173.235 -170.165 173.565 -169.835 ;
        RECT 173.235 -171.525 173.565 -171.195 ;
        RECT 173.235 -172.885 173.565 -172.555 ;
        RECT 173.235 -174.245 173.565 -173.915 ;
        RECT 173.235 -175.605 173.565 -175.275 ;
        RECT 173.235 -176.965 173.565 -176.635 ;
        RECT 173.235 -178.325 173.565 -177.995 ;
        RECT 173.235 -179.685 173.565 -179.355 ;
        RECT 173.235 -181.045 173.565 -180.715 ;
        RECT 173.235 -182.405 173.565 -182.075 ;
        RECT 173.235 -183.765 173.565 -183.435 ;
        RECT 173.235 -185.125 173.565 -184.795 ;
        RECT 173.235 -186.485 173.565 -186.155 ;
        RECT 173.235 -187.845 173.565 -187.515 ;
        RECT 173.235 -189.205 173.565 -188.875 ;
        RECT 173.235 -190.565 173.565 -190.235 ;
        RECT 173.235 -191.925 173.565 -191.595 ;
        RECT 173.235 -193.285 173.565 -192.955 ;
        RECT 173.235 -194.645 173.565 -194.315 ;
        RECT 173.235 -196.005 173.565 -195.675 ;
        RECT 173.235 -197.365 173.565 -197.035 ;
        RECT 173.235 -198.725 173.565 -198.395 ;
        RECT 173.235 -200.085 173.565 -199.755 ;
        RECT 173.235 -201.445 173.565 -201.115 ;
        RECT 173.235 -202.805 173.565 -202.475 ;
        RECT 173.235 -204.165 173.565 -203.835 ;
        RECT 173.235 -205.525 173.565 -205.195 ;
        RECT 173.235 -206.885 173.565 -206.555 ;
        RECT 173.235 -208.245 173.565 -207.915 ;
        RECT 173.235 -209.605 173.565 -209.275 ;
        RECT 173.235 -210.965 173.565 -210.635 ;
        RECT 173.235 -212.325 173.565 -211.995 ;
        RECT 173.235 -213.685 173.565 -213.355 ;
        RECT 173.235 -215.045 173.565 -214.715 ;
        RECT 173.235 -216.405 173.565 -216.075 ;
        RECT 173.235 -217.765 173.565 -217.435 ;
        RECT 173.235 -219.125 173.565 -218.795 ;
        RECT 173.235 -221.37 173.565 -220.24 ;
        RECT 173.24 -221.485 173.56 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.11 -121.535 174.44 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.595 129.8 174.925 130.93 ;
        RECT 174.595 127.675 174.925 128.005 ;
        RECT 174.595 126.315 174.925 126.645 ;
        RECT 174.595 124.955 174.925 125.285 ;
        RECT 174.595 123.595 174.925 123.925 ;
        RECT 174.6 123.595 174.92 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.955 129.8 176.285 130.93 ;
        RECT 175.955 127.675 176.285 128.005 ;
        RECT 175.955 126.315 176.285 126.645 ;
        RECT 175.955 124.955 176.285 125.285 ;
        RECT 175.955 123.595 176.285 123.925 ;
        RECT 175.96 123.595 176.28 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.955 -1.525 176.285 -1.195 ;
        RECT 175.955 -2.885 176.285 -2.555 ;
        RECT 175.96 -3.56 176.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.315 129.8 177.645 130.93 ;
        RECT 177.315 127.675 177.645 128.005 ;
        RECT 177.315 126.315 177.645 126.645 ;
        RECT 177.315 124.955 177.645 125.285 ;
        RECT 177.315 123.595 177.645 123.925 ;
        RECT 177.32 123.595 177.64 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.315 -1.525 177.645 -1.195 ;
        RECT 177.315 -2.885 177.645 -2.555 ;
        RECT 177.32 -3.56 177.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.315 -118.485 177.645 -118.155 ;
        RECT 177.315 -119.845 177.645 -119.515 ;
        RECT 177.315 -121.205 177.645 -120.875 ;
        RECT 177.315 -122.565 177.645 -122.235 ;
        RECT 177.315 -123.925 177.645 -123.595 ;
        RECT 177.315 -125.285 177.645 -124.955 ;
        RECT 177.315 -126.645 177.645 -126.315 ;
        RECT 177.315 -128.005 177.645 -127.675 ;
        RECT 177.315 -129.365 177.645 -129.035 ;
        RECT 177.315 -130.725 177.645 -130.395 ;
        RECT 177.315 -132.085 177.645 -131.755 ;
        RECT 177.315 -133.445 177.645 -133.115 ;
        RECT 177.315 -134.805 177.645 -134.475 ;
        RECT 177.315 -136.165 177.645 -135.835 ;
        RECT 177.315 -137.525 177.645 -137.195 ;
        RECT 177.315 -138.885 177.645 -138.555 ;
        RECT 177.315 -140.245 177.645 -139.915 ;
        RECT 177.315 -141.605 177.645 -141.275 ;
        RECT 177.315 -142.965 177.645 -142.635 ;
        RECT 177.315 -144.325 177.645 -143.995 ;
        RECT 177.315 -145.685 177.645 -145.355 ;
        RECT 177.315 -147.045 177.645 -146.715 ;
        RECT 177.315 -148.405 177.645 -148.075 ;
        RECT 177.315 -149.765 177.645 -149.435 ;
        RECT 177.315 -151.125 177.645 -150.795 ;
        RECT 177.315 -152.485 177.645 -152.155 ;
        RECT 177.315 -153.845 177.645 -153.515 ;
        RECT 177.315 -155.205 177.645 -154.875 ;
        RECT 177.315 -156.565 177.645 -156.235 ;
        RECT 177.315 -157.925 177.645 -157.595 ;
        RECT 177.315 -159.285 177.645 -158.955 ;
        RECT 177.315 -160.645 177.645 -160.315 ;
        RECT 177.315 -162.005 177.645 -161.675 ;
        RECT 177.315 -163.365 177.645 -163.035 ;
        RECT 177.315 -164.725 177.645 -164.395 ;
        RECT 177.315 -166.085 177.645 -165.755 ;
        RECT 177.315 -167.445 177.645 -167.115 ;
        RECT 177.315 -168.805 177.645 -168.475 ;
        RECT 177.315 -170.165 177.645 -169.835 ;
        RECT 177.315 -171.525 177.645 -171.195 ;
        RECT 177.315 -172.885 177.645 -172.555 ;
        RECT 177.315 -174.245 177.645 -173.915 ;
        RECT 177.315 -175.605 177.645 -175.275 ;
        RECT 177.315 -176.965 177.645 -176.635 ;
        RECT 177.315 -178.325 177.645 -177.995 ;
        RECT 177.315 -179.685 177.645 -179.355 ;
        RECT 177.315 -181.045 177.645 -180.715 ;
        RECT 177.315 -182.405 177.645 -182.075 ;
        RECT 177.315 -183.765 177.645 -183.435 ;
        RECT 177.315 -185.125 177.645 -184.795 ;
        RECT 177.315 -186.485 177.645 -186.155 ;
        RECT 177.315 -187.845 177.645 -187.515 ;
        RECT 177.315 -189.205 177.645 -188.875 ;
        RECT 177.315 -190.565 177.645 -190.235 ;
        RECT 177.315 -191.925 177.645 -191.595 ;
        RECT 177.315 -193.285 177.645 -192.955 ;
        RECT 177.315 -194.645 177.645 -194.315 ;
        RECT 177.315 -196.005 177.645 -195.675 ;
        RECT 177.315 -197.365 177.645 -197.035 ;
        RECT 177.315 -198.725 177.645 -198.395 ;
        RECT 177.315 -200.085 177.645 -199.755 ;
        RECT 177.315 -201.445 177.645 -201.115 ;
        RECT 177.315 -202.805 177.645 -202.475 ;
        RECT 177.315 -204.165 177.645 -203.835 ;
        RECT 177.315 -205.525 177.645 -205.195 ;
        RECT 177.315 -206.885 177.645 -206.555 ;
        RECT 177.315 -208.245 177.645 -207.915 ;
        RECT 177.315 -209.605 177.645 -209.275 ;
        RECT 177.315 -210.965 177.645 -210.635 ;
        RECT 177.315 -212.325 177.645 -211.995 ;
        RECT 177.315 -213.685 177.645 -213.355 ;
        RECT 177.315 -215.045 177.645 -214.715 ;
        RECT 177.315 -216.405 177.645 -216.075 ;
        RECT 177.315 -217.765 177.645 -217.435 ;
        RECT 177.315 -219.125 177.645 -218.795 ;
        RECT 177.315 -221.37 177.645 -220.24 ;
        RECT 177.32 -221.485 177.64 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.675 129.8 179.005 130.93 ;
        RECT 178.675 127.675 179.005 128.005 ;
        RECT 178.675 126.315 179.005 126.645 ;
        RECT 178.675 124.955 179.005 125.285 ;
        RECT 178.675 123.595 179.005 123.925 ;
        RECT 178.68 123.595 179 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.675 -1.525 179.005 -1.195 ;
        RECT 178.675 -2.885 179.005 -2.555 ;
        RECT 178.68 -3.56 179 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.675 -118.485 179.005 -118.155 ;
        RECT 178.675 -119.845 179.005 -119.515 ;
        RECT 178.675 -121.205 179.005 -120.875 ;
        RECT 178.675 -122.565 179.005 -122.235 ;
        RECT 178.675 -123.925 179.005 -123.595 ;
        RECT 178.675 -125.285 179.005 -124.955 ;
        RECT 178.675 -126.645 179.005 -126.315 ;
        RECT 178.675 -128.005 179.005 -127.675 ;
        RECT 178.675 -129.365 179.005 -129.035 ;
        RECT 178.675 -130.725 179.005 -130.395 ;
        RECT 178.675 -132.085 179.005 -131.755 ;
        RECT 178.675 -133.445 179.005 -133.115 ;
        RECT 178.675 -134.805 179.005 -134.475 ;
        RECT 178.675 -136.165 179.005 -135.835 ;
        RECT 178.675 -137.525 179.005 -137.195 ;
        RECT 178.675 -138.885 179.005 -138.555 ;
        RECT 178.675 -140.245 179.005 -139.915 ;
        RECT 178.675 -141.605 179.005 -141.275 ;
        RECT 178.675 -142.965 179.005 -142.635 ;
        RECT 178.675 -144.325 179.005 -143.995 ;
        RECT 178.675 -145.685 179.005 -145.355 ;
        RECT 178.675 -147.045 179.005 -146.715 ;
        RECT 178.675 -148.405 179.005 -148.075 ;
        RECT 178.675 -149.765 179.005 -149.435 ;
        RECT 178.675 -151.125 179.005 -150.795 ;
        RECT 178.675 -152.485 179.005 -152.155 ;
        RECT 178.675 -153.845 179.005 -153.515 ;
        RECT 178.675 -155.205 179.005 -154.875 ;
        RECT 178.675 -156.565 179.005 -156.235 ;
        RECT 178.675 -157.925 179.005 -157.595 ;
        RECT 178.675 -159.285 179.005 -158.955 ;
        RECT 178.675 -160.645 179.005 -160.315 ;
        RECT 178.675 -162.005 179.005 -161.675 ;
        RECT 178.675 -163.365 179.005 -163.035 ;
        RECT 178.675 -164.725 179.005 -164.395 ;
        RECT 178.675 -166.085 179.005 -165.755 ;
        RECT 178.675 -167.445 179.005 -167.115 ;
        RECT 178.675 -168.805 179.005 -168.475 ;
        RECT 178.675 -170.165 179.005 -169.835 ;
        RECT 178.675 -171.525 179.005 -171.195 ;
        RECT 178.675 -172.885 179.005 -172.555 ;
        RECT 178.675 -174.245 179.005 -173.915 ;
        RECT 178.675 -175.605 179.005 -175.275 ;
        RECT 178.675 -176.965 179.005 -176.635 ;
        RECT 178.675 -178.325 179.005 -177.995 ;
        RECT 178.675 -179.685 179.005 -179.355 ;
        RECT 178.675 -181.045 179.005 -180.715 ;
        RECT 178.675 -182.405 179.005 -182.075 ;
        RECT 178.675 -183.765 179.005 -183.435 ;
        RECT 178.675 -185.125 179.005 -184.795 ;
        RECT 178.675 -186.485 179.005 -186.155 ;
        RECT 178.675 -187.845 179.005 -187.515 ;
        RECT 178.675 -189.205 179.005 -188.875 ;
        RECT 178.675 -190.565 179.005 -190.235 ;
        RECT 178.675 -191.925 179.005 -191.595 ;
        RECT 178.675 -193.285 179.005 -192.955 ;
        RECT 178.675 -194.645 179.005 -194.315 ;
        RECT 178.675 -196.005 179.005 -195.675 ;
        RECT 178.675 -197.365 179.005 -197.035 ;
        RECT 178.675 -198.725 179.005 -198.395 ;
        RECT 178.675 -200.085 179.005 -199.755 ;
        RECT 178.675 -201.445 179.005 -201.115 ;
        RECT 178.675 -202.805 179.005 -202.475 ;
        RECT 178.675 -204.165 179.005 -203.835 ;
        RECT 178.675 -205.525 179.005 -205.195 ;
        RECT 178.675 -206.885 179.005 -206.555 ;
        RECT 178.675 -208.245 179.005 -207.915 ;
        RECT 178.675 -209.605 179.005 -209.275 ;
        RECT 178.675 -210.965 179.005 -210.635 ;
        RECT 178.675 -212.325 179.005 -211.995 ;
        RECT 178.675 -213.685 179.005 -213.355 ;
        RECT 178.675 -215.045 179.005 -214.715 ;
        RECT 178.675 -216.405 179.005 -216.075 ;
        RECT 178.675 -217.765 179.005 -217.435 ;
        RECT 178.675 -219.125 179.005 -218.795 ;
        RECT 178.675 -221.37 179.005 -220.24 ;
        RECT 178.68 -221.485 179 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.035 129.8 180.365 130.93 ;
        RECT 180.035 127.675 180.365 128.005 ;
        RECT 180.035 126.315 180.365 126.645 ;
        RECT 180.035 124.955 180.365 125.285 ;
        RECT 180.035 123.595 180.365 123.925 ;
        RECT 180.04 123.595 180.36 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.035 -122.565 180.365 -122.235 ;
        RECT 180.035 -123.925 180.365 -123.595 ;
        RECT 180.035 -125.285 180.365 -124.955 ;
        RECT 180.035 -126.645 180.365 -126.315 ;
        RECT 180.035 -128.005 180.365 -127.675 ;
        RECT 180.035 -129.365 180.365 -129.035 ;
        RECT 180.035 -130.725 180.365 -130.395 ;
        RECT 180.035 -132.085 180.365 -131.755 ;
        RECT 180.035 -133.445 180.365 -133.115 ;
        RECT 180.035 -134.805 180.365 -134.475 ;
        RECT 180.035 -136.165 180.365 -135.835 ;
        RECT 180.035 -137.525 180.365 -137.195 ;
        RECT 180.035 -138.885 180.365 -138.555 ;
        RECT 180.035 -140.245 180.365 -139.915 ;
        RECT 180.035 -141.605 180.365 -141.275 ;
        RECT 180.035 -142.965 180.365 -142.635 ;
        RECT 180.035 -144.325 180.365 -143.995 ;
        RECT 180.035 -145.685 180.365 -145.355 ;
        RECT 180.035 -147.045 180.365 -146.715 ;
        RECT 180.035 -148.405 180.365 -148.075 ;
        RECT 180.035 -149.765 180.365 -149.435 ;
        RECT 180.035 -151.125 180.365 -150.795 ;
        RECT 180.035 -152.485 180.365 -152.155 ;
        RECT 180.035 -153.845 180.365 -153.515 ;
        RECT 180.035 -155.205 180.365 -154.875 ;
        RECT 180.035 -156.565 180.365 -156.235 ;
        RECT 180.035 -157.925 180.365 -157.595 ;
        RECT 180.035 -159.285 180.365 -158.955 ;
        RECT 180.035 -160.645 180.365 -160.315 ;
        RECT 180.035 -162.005 180.365 -161.675 ;
        RECT 180.035 -163.365 180.365 -163.035 ;
        RECT 180.035 -164.725 180.365 -164.395 ;
        RECT 180.035 -166.085 180.365 -165.755 ;
        RECT 180.035 -167.445 180.365 -167.115 ;
        RECT 180.035 -168.805 180.365 -168.475 ;
        RECT 180.035 -170.165 180.365 -169.835 ;
        RECT 180.035 -171.525 180.365 -171.195 ;
        RECT 180.035 -172.885 180.365 -172.555 ;
        RECT 180.035 -174.245 180.365 -173.915 ;
        RECT 180.035 -175.605 180.365 -175.275 ;
        RECT 180.035 -176.965 180.365 -176.635 ;
        RECT 180.035 -178.325 180.365 -177.995 ;
        RECT 180.035 -179.685 180.365 -179.355 ;
        RECT 180.035 -181.045 180.365 -180.715 ;
        RECT 180.035 -182.405 180.365 -182.075 ;
        RECT 180.035 -183.765 180.365 -183.435 ;
        RECT 180.035 -185.125 180.365 -184.795 ;
        RECT 180.035 -186.485 180.365 -186.155 ;
        RECT 180.035 -187.845 180.365 -187.515 ;
        RECT 180.035 -189.205 180.365 -188.875 ;
        RECT 180.035 -190.565 180.365 -190.235 ;
        RECT 180.035 -191.925 180.365 -191.595 ;
        RECT 180.035 -193.285 180.365 -192.955 ;
        RECT 180.035 -194.645 180.365 -194.315 ;
        RECT 180.035 -196.005 180.365 -195.675 ;
        RECT 180.035 -197.365 180.365 -197.035 ;
        RECT 180.035 -198.725 180.365 -198.395 ;
        RECT 180.035 -200.085 180.365 -199.755 ;
        RECT 180.035 -201.445 180.365 -201.115 ;
        RECT 180.035 -202.805 180.365 -202.475 ;
        RECT 180.035 -204.165 180.365 -203.835 ;
        RECT 180.035 -205.525 180.365 -205.195 ;
        RECT 180.035 -206.885 180.365 -206.555 ;
        RECT 180.035 -208.245 180.365 -207.915 ;
        RECT 180.035 -209.605 180.365 -209.275 ;
        RECT 180.035 -210.965 180.365 -210.635 ;
        RECT 180.035 -212.325 180.365 -211.995 ;
        RECT 180.035 -213.685 180.365 -213.355 ;
        RECT 180.035 -215.045 180.365 -214.715 ;
        RECT 180.035 -216.405 180.365 -216.075 ;
        RECT 180.035 -217.765 180.365 -217.435 ;
        RECT 180.035 -219.125 180.365 -218.795 ;
        RECT 180.035 -221.37 180.365 -220.24 ;
        RECT 180.04 -221.485 180.36 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.21 -121.535 180.54 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 181.395 129.8 181.725 130.93 ;
        RECT 181.395 127.675 181.725 128.005 ;
        RECT 181.395 126.315 181.725 126.645 ;
        RECT 181.395 124.955 181.725 125.285 ;
        RECT 181.395 123.595 181.725 123.925 ;
        RECT 181.4 123.595 181.72 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 181.395 -1.525 181.725 -1.195 ;
        RECT 181.395 -2.885 181.725 -2.555 ;
        RECT 181.4 -3.56 181.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.755 129.8 183.085 130.93 ;
        RECT 182.755 127.675 183.085 128.005 ;
        RECT 182.755 126.315 183.085 126.645 ;
        RECT 182.755 124.955 183.085 125.285 ;
        RECT 182.755 123.595 183.085 123.925 ;
        RECT 182.76 123.595 183.08 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.755 -1.525 183.085 -1.195 ;
        RECT 182.755 -2.885 183.085 -2.555 ;
        RECT 182.76 -3.56 183.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.115 129.8 184.445 130.93 ;
        RECT 184.115 127.675 184.445 128.005 ;
        RECT 184.115 126.315 184.445 126.645 ;
        RECT 184.115 124.955 184.445 125.285 ;
        RECT 184.115 123.595 184.445 123.925 ;
        RECT 184.12 123.595 184.44 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.115 -1.525 184.445 -1.195 ;
        RECT 184.115 -2.885 184.445 -2.555 ;
        RECT 184.12 -3.56 184.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.115 -118.485 184.445 -118.155 ;
        RECT 184.115 -119.845 184.445 -119.515 ;
        RECT 184.115 -121.205 184.445 -120.875 ;
        RECT 184.115 -122.565 184.445 -122.235 ;
        RECT 184.115 -123.925 184.445 -123.595 ;
        RECT 184.115 -125.285 184.445 -124.955 ;
        RECT 184.115 -126.645 184.445 -126.315 ;
        RECT 184.115 -128.005 184.445 -127.675 ;
        RECT 184.115 -129.365 184.445 -129.035 ;
        RECT 184.115 -130.725 184.445 -130.395 ;
        RECT 184.115 -132.085 184.445 -131.755 ;
        RECT 184.115 -133.445 184.445 -133.115 ;
        RECT 184.115 -134.805 184.445 -134.475 ;
        RECT 184.115 -136.165 184.445 -135.835 ;
        RECT 184.115 -137.525 184.445 -137.195 ;
        RECT 184.115 -138.885 184.445 -138.555 ;
        RECT 184.115 -140.245 184.445 -139.915 ;
        RECT 184.115 -141.605 184.445 -141.275 ;
        RECT 184.115 -142.965 184.445 -142.635 ;
        RECT 184.115 -144.325 184.445 -143.995 ;
        RECT 184.115 -145.685 184.445 -145.355 ;
        RECT 184.115 -147.045 184.445 -146.715 ;
        RECT 184.115 -148.405 184.445 -148.075 ;
        RECT 184.115 -149.765 184.445 -149.435 ;
        RECT 184.115 -151.125 184.445 -150.795 ;
        RECT 184.115 -152.485 184.445 -152.155 ;
        RECT 184.115 -153.845 184.445 -153.515 ;
        RECT 184.115 -155.205 184.445 -154.875 ;
        RECT 184.115 -156.565 184.445 -156.235 ;
        RECT 184.115 -157.925 184.445 -157.595 ;
        RECT 184.115 -159.285 184.445 -158.955 ;
        RECT 184.115 -160.645 184.445 -160.315 ;
        RECT 184.115 -162.005 184.445 -161.675 ;
        RECT 184.115 -163.365 184.445 -163.035 ;
        RECT 184.115 -164.725 184.445 -164.395 ;
        RECT 184.115 -166.085 184.445 -165.755 ;
        RECT 184.115 -167.445 184.445 -167.115 ;
        RECT 184.115 -168.805 184.445 -168.475 ;
        RECT 184.115 -170.165 184.445 -169.835 ;
        RECT 184.115 -171.525 184.445 -171.195 ;
        RECT 184.115 -172.885 184.445 -172.555 ;
        RECT 184.115 -174.245 184.445 -173.915 ;
        RECT 184.115 -175.605 184.445 -175.275 ;
        RECT 184.115 -176.965 184.445 -176.635 ;
        RECT 184.115 -178.325 184.445 -177.995 ;
        RECT 184.115 -179.685 184.445 -179.355 ;
        RECT 184.115 -181.045 184.445 -180.715 ;
        RECT 184.115 -182.405 184.445 -182.075 ;
        RECT 184.115 -183.765 184.445 -183.435 ;
        RECT 184.115 -185.125 184.445 -184.795 ;
        RECT 184.115 -186.485 184.445 -186.155 ;
        RECT 184.115 -187.845 184.445 -187.515 ;
        RECT 184.115 -189.205 184.445 -188.875 ;
        RECT 184.115 -190.565 184.445 -190.235 ;
        RECT 184.115 -191.925 184.445 -191.595 ;
        RECT 184.115 -193.285 184.445 -192.955 ;
        RECT 184.115 -194.645 184.445 -194.315 ;
        RECT 184.115 -196.005 184.445 -195.675 ;
        RECT 184.115 -197.365 184.445 -197.035 ;
        RECT 184.115 -198.725 184.445 -198.395 ;
        RECT 184.115 -200.085 184.445 -199.755 ;
        RECT 184.115 -201.445 184.445 -201.115 ;
        RECT 184.115 -202.805 184.445 -202.475 ;
        RECT 184.115 -204.165 184.445 -203.835 ;
        RECT 184.115 -205.525 184.445 -205.195 ;
        RECT 184.115 -206.885 184.445 -206.555 ;
        RECT 184.115 -208.245 184.445 -207.915 ;
        RECT 184.115 -209.605 184.445 -209.275 ;
        RECT 184.115 -210.965 184.445 -210.635 ;
        RECT 184.115 -212.325 184.445 -211.995 ;
        RECT 184.115 -213.685 184.445 -213.355 ;
        RECT 184.115 -215.045 184.445 -214.715 ;
        RECT 184.115 -216.405 184.445 -216.075 ;
        RECT 184.115 -217.765 184.445 -217.435 ;
        RECT 184.115 -219.125 184.445 -218.795 ;
        RECT 184.115 -221.37 184.445 -220.24 ;
        RECT 184.12 -221.485 184.44 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.475 129.8 185.805 130.93 ;
        RECT 185.475 127.675 185.805 128.005 ;
        RECT 185.475 126.315 185.805 126.645 ;
        RECT 185.475 124.955 185.805 125.285 ;
        RECT 185.475 123.595 185.805 123.925 ;
        RECT 185.48 123.595 185.8 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.475 -122.565 185.805 -122.235 ;
        RECT 185.475 -123.925 185.805 -123.595 ;
        RECT 185.475 -125.285 185.805 -124.955 ;
        RECT 185.475 -126.645 185.805 -126.315 ;
        RECT 185.475 -128.005 185.805 -127.675 ;
        RECT 185.475 -129.365 185.805 -129.035 ;
        RECT 185.475 -130.725 185.805 -130.395 ;
        RECT 185.475 -132.085 185.805 -131.755 ;
        RECT 185.475 -133.445 185.805 -133.115 ;
        RECT 185.475 -134.805 185.805 -134.475 ;
        RECT 185.475 -136.165 185.805 -135.835 ;
        RECT 185.475 -137.525 185.805 -137.195 ;
        RECT 185.475 -138.885 185.805 -138.555 ;
        RECT 185.475 -140.245 185.805 -139.915 ;
        RECT 185.475 -141.605 185.805 -141.275 ;
        RECT 185.475 -142.965 185.805 -142.635 ;
        RECT 185.475 -144.325 185.805 -143.995 ;
        RECT 185.475 -145.685 185.805 -145.355 ;
        RECT 185.475 -147.045 185.805 -146.715 ;
        RECT 185.475 -148.405 185.805 -148.075 ;
        RECT 185.475 -149.765 185.805 -149.435 ;
        RECT 185.475 -151.125 185.805 -150.795 ;
        RECT 185.475 -152.485 185.805 -152.155 ;
        RECT 185.475 -153.845 185.805 -153.515 ;
        RECT 185.475 -155.205 185.805 -154.875 ;
        RECT 185.475 -156.565 185.805 -156.235 ;
        RECT 185.475 -157.925 185.805 -157.595 ;
        RECT 185.475 -159.285 185.805 -158.955 ;
        RECT 185.475 -160.645 185.805 -160.315 ;
        RECT 185.475 -162.005 185.805 -161.675 ;
        RECT 185.475 -163.365 185.805 -163.035 ;
        RECT 185.475 -164.725 185.805 -164.395 ;
        RECT 185.475 -166.085 185.805 -165.755 ;
        RECT 185.475 -167.445 185.805 -167.115 ;
        RECT 185.475 -168.805 185.805 -168.475 ;
        RECT 185.475 -170.165 185.805 -169.835 ;
        RECT 185.475 -171.525 185.805 -171.195 ;
        RECT 185.475 -172.885 185.805 -172.555 ;
        RECT 185.475 -174.245 185.805 -173.915 ;
        RECT 185.475 -175.605 185.805 -175.275 ;
        RECT 185.475 -176.965 185.805 -176.635 ;
        RECT 185.475 -178.325 185.805 -177.995 ;
        RECT 185.475 -179.685 185.805 -179.355 ;
        RECT 185.475 -181.045 185.805 -180.715 ;
        RECT 185.475 -182.405 185.805 -182.075 ;
        RECT 185.475 -183.765 185.805 -183.435 ;
        RECT 185.475 -185.125 185.805 -184.795 ;
        RECT 185.475 -186.485 185.805 -186.155 ;
        RECT 185.475 -187.845 185.805 -187.515 ;
        RECT 185.475 -189.205 185.805 -188.875 ;
        RECT 185.475 -190.565 185.805 -190.235 ;
        RECT 185.475 -191.925 185.805 -191.595 ;
        RECT 185.475 -193.285 185.805 -192.955 ;
        RECT 185.475 -194.645 185.805 -194.315 ;
        RECT 185.475 -196.005 185.805 -195.675 ;
        RECT 185.475 -197.365 185.805 -197.035 ;
        RECT 185.475 -198.725 185.805 -198.395 ;
        RECT 185.475 -200.085 185.805 -199.755 ;
        RECT 185.475 -201.445 185.805 -201.115 ;
        RECT 185.475 -202.805 185.805 -202.475 ;
        RECT 185.475 -204.165 185.805 -203.835 ;
        RECT 185.475 -205.525 185.805 -205.195 ;
        RECT 185.475 -206.885 185.805 -206.555 ;
        RECT 185.475 -208.245 185.805 -207.915 ;
        RECT 185.475 -209.605 185.805 -209.275 ;
        RECT 185.475 -210.965 185.805 -210.635 ;
        RECT 185.475 -212.325 185.805 -211.995 ;
        RECT 185.475 -213.685 185.805 -213.355 ;
        RECT 185.475 -215.045 185.805 -214.715 ;
        RECT 185.475 -216.405 185.805 -216.075 ;
        RECT 185.475 -217.765 185.805 -217.435 ;
        RECT 185.475 -219.125 185.805 -218.795 ;
        RECT 185.475 -221.37 185.805 -220.24 ;
        RECT 185.48 -221.485 185.8 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.31 -121.535 186.64 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.835 129.8 187.165 130.93 ;
        RECT 186.835 127.675 187.165 128.005 ;
        RECT 186.835 126.315 187.165 126.645 ;
        RECT 186.835 124.955 187.165 125.285 ;
        RECT 186.835 123.595 187.165 123.925 ;
        RECT 186.84 123.595 187.16 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.195 129.8 188.525 130.93 ;
        RECT 188.195 127.675 188.525 128.005 ;
        RECT 188.195 126.315 188.525 126.645 ;
        RECT 188.195 124.955 188.525 125.285 ;
        RECT 188.195 123.595 188.525 123.925 ;
        RECT 188.2 123.595 188.52 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.195 -1.525 188.525 -1.195 ;
        RECT 188.195 -2.885 188.525 -2.555 ;
        RECT 188.2 -3.56 188.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.555 129.8 189.885 130.93 ;
        RECT 189.555 127.675 189.885 128.005 ;
        RECT 189.555 126.315 189.885 126.645 ;
        RECT 189.555 124.955 189.885 125.285 ;
        RECT 189.555 123.595 189.885 123.925 ;
        RECT 189.56 123.595 189.88 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.555 -1.525 189.885 -1.195 ;
        RECT 189.555 -2.885 189.885 -2.555 ;
        RECT 189.56 -3.56 189.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.555 -118.485 189.885 -118.155 ;
        RECT 189.555 -119.845 189.885 -119.515 ;
        RECT 189.555 -121.205 189.885 -120.875 ;
        RECT 189.555 -122.565 189.885 -122.235 ;
        RECT 189.555 -123.925 189.885 -123.595 ;
        RECT 189.555 -125.285 189.885 -124.955 ;
        RECT 189.555 -126.645 189.885 -126.315 ;
        RECT 189.555 -128.005 189.885 -127.675 ;
        RECT 189.555 -129.365 189.885 -129.035 ;
        RECT 189.555 -130.725 189.885 -130.395 ;
        RECT 189.555 -132.085 189.885 -131.755 ;
        RECT 189.555 -133.445 189.885 -133.115 ;
        RECT 189.555 -134.805 189.885 -134.475 ;
        RECT 189.555 -136.165 189.885 -135.835 ;
        RECT 189.555 -137.525 189.885 -137.195 ;
        RECT 189.555 -138.885 189.885 -138.555 ;
        RECT 189.555 -140.245 189.885 -139.915 ;
        RECT 189.555 -141.605 189.885 -141.275 ;
        RECT 189.555 -142.965 189.885 -142.635 ;
        RECT 189.555 -144.325 189.885 -143.995 ;
        RECT 189.555 -145.685 189.885 -145.355 ;
        RECT 189.555 -147.045 189.885 -146.715 ;
        RECT 189.555 -148.405 189.885 -148.075 ;
        RECT 189.555 -149.765 189.885 -149.435 ;
        RECT 189.555 -151.125 189.885 -150.795 ;
        RECT 189.555 -152.485 189.885 -152.155 ;
        RECT 189.555 -153.845 189.885 -153.515 ;
        RECT 189.555 -155.205 189.885 -154.875 ;
        RECT 189.555 -156.565 189.885 -156.235 ;
        RECT 189.555 -157.925 189.885 -157.595 ;
        RECT 189.555 -159.285 189.885 -158.955 ;
        RECT 189.555 -160.645 189.885 -160.315 ;
        RECT 189.555 -162.005 189.885 -161.675 ;
        RECT 189.555 -163.365 189.885 -163.035 ;
        RECT 189.555 -164.725 189.885 -164.395 ;
        RECT 189.555 -166.085 189.885 -165.755 ;
        RECT 189.555 -167.445 189.885 -167.115 ;
        RECT 189.555 -168.805 189.885 -168.475 ;
        RECT 189.555 -170.165 189.885 -169.835 ;
        RECT 189.555 -171.525 189.885 -171.195 ;
        RECT 189.555 -172.885 189.885 -172.555 ;
        RECT 189.555 -174.245 189.885 -173.915 ;
        RECT 189.555 -175.605 189.885 -175.275 ;
        RECT 189.555 -176.965 189.885 -176.635 ;
        RECT 189.555 -178.325 189.885 -177.995 ;
        RECT 189.555 -179.685 189.885 -179.355 ;
        RECT 189.555 -181.045 189.885 -180.715 ;
        RECT 189.555 -182.405 189.885 -182.075 ;
        RECT 189.555 -183.765 189.885 -183.435 ;
        RECT 189.555 -185.125 189.885 -184.795 ;
        RECT 189.555 -186.485 189.885 -186.155 ;
        RECT 189.555 -187.845 189.885 -187.515 ;
        RECT 189.555 -189.205 189.885 -188.875 ;
        RECT 189.555 -190.565 189.885 -190.235 ;
        RECT 189.555 -191.925 189.885 -191.595 ;
        RECT 189.555 -193.285 189.885 -192.955 ;
        RECT 189.555 -194.645 189.885 -194.315 ;
        RECT 189.555 -196.005 189.885 -195.675 ;
        RECT 189.555 -197.365 189.885 -197.035 ;
        RECT 189.555 -198.725 189.885 -198.395 ;
        RECT 189.555 -200.085 189.885 -199.755 ;
        RECT 189.555 -201.445 189.885 -201.115 ;
        RECT 189.555 -202.805 189.885 -202.475 ;
        RECT 189.555 -204.165 189.885 -203.835 ;
        RECT 189.555 -205.525 189.885 -205.195 ;
        RECT 189.555 -206.885 189.885 -206.555 ;
        RECT 189.555 -208.245 189.885 -207.915 ;
        RECT 189.555 -209.605 189.885 -209.275 ;
        RECT 189.555 -210.965 189.885 -210.635 ;
        RECT 189.555 -212.325 189.885 -211.995 ;
        RECT 189.555 -213.685 189.885 -213.355 ;
        RECT 189.555 -215.045 189.885 -214.715 ;
        RECT 189.555 -216.405 189.885 -216.075 ;
        RECT 189.555 -217.765 189.885 -217.435 ;
        RECT 189.555 -219.125 189.885 -218.795 ;
        RECT 189.555 -221.37 189.885 -220.24 ;
        RECT 189.56 -221.485 189.88 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.915 129.8 191.245 130.93 ;
        RECT 190.915 127.675 191.245 128.005 ;
        RECT 190.915 126.315 191.245 126.645 ;
        RECT 190.915 124.955 191.245 125.285 ;
        RECT 190.915 123.595 191.245 123.925 ;
        RECT 190.92 123.595 191.24 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.915 -1.525 191.245 -1.195 ;
        RECT 190.915 -2.885 191.245 -2.555 ;
        RECT 190.92 -3.56 191.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.915 -202.805 191.245 -202.475 ;
        RECT 190.915 -204.165 191.245 -203.835 ;
        RECT 190.915 -205.525 191.245 -205.195 ;
        RECT 190.915 -206.885 191.245 -206.555 ;
        RECT 190.915 -208.245 191.245 -207.915 ;
        RECT 190.915 -209.605 191.245 -209.275 ;
        RECT 190.915 -210.965 191.245 -210.635 ;
        RECT 190.915 -212.325 191.245 -211.995 ;
        RECT 190.915 -213.685 191.245 -213.355 ;
        RECT 190.915 -215.045 191.245 -214.715 ;
        RECT 190.915 -216.405 191.245 -216.075 ;
        RECT 190.915 -217.765 191.245 -217.435 ;
        RECT 190.915 -219.125 191.245 -218.795 ;
        RECT 190.915 -221.37 191.245 -220.24 ;
        RECT 190.92 -221.485 191.24 -118.155 ;
        RECT 190.915 -118.485 191.245 -118.155 ;
        RECT 190.915 -119.845 191.245 -119.515 ;
        RECT 190.915 -121.205 191.245 -120.875 ;
        RECT 190.915 -122.565 191.245 -122.235 ;
        RECT 190.915 -123.925 191.245 -123.595 ;
        RECT 190.915 -125.285 191.245 -124.955 ;
        RECT 190.915 -126.645 191.245 -126.315 ;
        RECT 190.915 -128.005 191.245 -127.675 ;
        RECT 190.915 -129.365 191.245 -129.035 ;
        RECT 190.915 -130.725 191.245 -130.395 ;
        RECT 190.915 -132.085 191.245 -131.755 ;
        RECT 190.915 -133.445 191.245 -133.115 ;
        RECT 190.915 -134.805 191.245 -134.475 ;
        RECT 190.915 -136.165 191.245 -135.835 ;
        RECT 190.915 -137.525 191.245 -137.195 ;
        RECT 190.915 -138.885 191.245 -138.555 ;
        RECT 190.915 -140.245 191.245 -139.915 ;
        RECT 190.915 -141.605 191.245 -141.275 ;
        RECT 190.915 -142.965 191.245 -142.635 ;
        RECT 190.915 -144.325 191.245 -143.995 ;
        RECT 190.915 -145.685 191.245 -145.355 ;
        RECT 190.915 -147.045 191.245 -146.715 ;
        RECT 190.915 -148.405 191.245 -148.075 ;
        RECT 190.915 -149.765 191.245 -149.435 ;
        RECT 190.915 -151.125 191.245 -150.795 ;
        RECT 190.915 -152.485 191.245 -152.155 ;
        RECT 190.915 -153.845 191.245 -153.515 ;
        RECT 190.915 -155.205 191.245 -154.875 ;
        RECT 190.915 -156.565 191.245 -156.235 ;
        RECT 190.915 -157.925 191.245 -157.595 ;
        RECT 190.915 -159.285 191.245 -158.955 ;
        RECT 190.915 -160.645 191.245 -160.315 ;
        RECT 190.915 -162.005 191.245 -161.675 ;
        RECT 190.915 -163.365 191.245 -163.035 ;
        RECT 190.915 -164.725 191.245 -164.395 ;
        RECT 190.915 -166.085 191.245 -165.755 ;
        RECT 190.915 -167.445 191.245 -167.115 ;
        RECT 190.915 -168.805 191.245 -168.475 ;
        RECT 190.915 -170.165 191.245 -169.835 ;
        RECT 190.915 -171.525 191.245 -171.195 ;
        RECT 190.915 -172.885 191.245 -172.555 ;
        RECT 190.915 -174.245 191.245 -173.915 ;
        RECT 190.915 -175.605 191.245 -175.275 ;
        RECT 190.915 -176.965 191.245 -176.635 ;
        RECT 190.915 -178.325 191.245 -177.995 ;
        RECT 190.915 -179.685 191.245 -179.355 ;
        RECT 190.915 -181.045 191.245 -180.715 ;
        RECT 190.915 -182.405 191.245 -182.075 ;
        RECT 190.915 -183.765 191.245 -183.435 ;
        RECT 190.915 -185.125 191.245 -184.795 ;
        RECT 190.915 -186.485 191.245 -186.155 ;
        RECT 190.915 -187.845 191.245 -187.515 ;
        RECT 190.915 -189.205 191.245 -188.875 ;
        RECT 190.915 -190.565 191.245 -190.235 ;
        RECT 190.915 -191.925 191.245 -191.595 ;
        RECT 190.915 -193.285 191.245 -192.955 ;
        RECT 190.915 -194.645 191.245 -194.315 ;
        RECT 190.915 -196.005 191.245 -195.675 ;
        RECT 190.915 -197.365 191.245 -197.035 ;
        RECT 190.915 -198.725 191.245 -198.395 ;
        RECT 190.915 -200.085 191.245 -199.755 ;
        RECT 190.915 -201.445 191.245 -201.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.515 129.8 136.845 130.93 ;
        RECT 136.515 127.675 136.845 128.005 ;
        RECT 136.515 126.315 136.845 126.645 ;
        RECT 136.515 124.955 136.845 125.285 ;
        RECT 136.515 123.595 136.845 123.925 ;
        RECT 136.52 123.595 136.84 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.515 -122.565 136.845 -122.235 ;
        RECT 136.515 -123.925 136.845 -123.595 ;
        RECT 136.515 -125.285 136.845 -124.955 ;
        RECT 136.515 -126.645 136.845 -126.315 ;
        RECT 136.515 -128.005 136.845 -127.675 ;
        RECT 136.515 -129.365 136.845 -129.035 ;
        RECT 136.515 -130.725 136.845 -130.395 ;
        RECT 136.515 -132.085 136.845 -131.755 ;
        RECT 136.515 -133.445 136.845 -133.115 ;
        RECT 136.515 -134.805 136.845 -134.475 ;
        RECT 136.515 -136.165 136.845 -135.835 ;
        RECT 136.515 -137.525 136.845 -137.195 ;
        RECT 136.515 -138.885 136.845 -138.555 ;
        RECT 136.515 -140.245 136.845 -139.915 ;
        RECT 136.515 -141.605 136.845 -141.275 ;
        RECT 136.515 -142.965 136.845 -142.635 ;
        RECT 136.515 -144.325 136.845 -143.995 ;
        RECT 136.515 -145.685 136.845 -145.355 ;
        RECT 136.515 -147.045 136.845 -146.715 ;
        RECT 136.515 -148.405 136.845 -148.075 ;
        RECT 136.515 -149.765 136.845 -149.435 ;
        RECT 136.515 -151.125 136.845 -150.795 ;
        RECT 136.515 -152.485 136.845 -152.155 ;
        RECT 136.515 -153.845 136.845 -153.515 ;
        RECT 136.515 -155.205 136.845 -154.875 ;
        RECT 136.515 -156.565 136.845 -156.235 ;
        RECT 136.515 -157.925 136.845 -157.595 ;
        RECT 136.515 -159.285 136.845 -158.955 ;
        RECT 136.515 -160.645 136.845 -160.315 ;
        RECT 136.515 -162.005 136.845 -161.675 ;
        RECT 136.515 -163.365 136.845 -163.035 ;
        RECT 136.515 -164.725 136.845 -164.395 ;
        RECT 136.515 -166.085 136.845 -165.755 ;
        RECT 136.515 -167.445 136.845 -167.115 ;
        RECT 136.515 -168.805 136.845 -168.475 ;
        RECT 136.515 -170.165 136.845 -169.835 ;
        RECT 136.515 -171.525 136.845 -171.195 ;
        RECT 136.515 -172.885 136.845 -172.555 ;
        RECT 136.515 -174.245 136.845 -173.915 ;
        RECT 136.515 -175.605 136.845 -175.275 ;
        RECT 136.515 -176.965 136.845 -176.635 ;
        RECT 136.515 -178.325 136.845 -177.995 ;
        RECT 136.515 -179.685 136.845 -179.355 ;
        RECT 136.515 -181.045 136.845 -180.715 ;
        RECT 136.515 -182.405 136.845 -182.075 ;
        RECT 136.515 -183.765 136.845 -183.435 ;
        RECT 136.515 -185.125 136.845 -184.795 ;
        RECT 136.515 -186.485 136.845 -186.155 ;
        RECT 136.515 -187.845 136.845 -187.515 ;
        RECT 136.515 -189.205 136.845 -188.875 ;
        RECT 136.515 -190.565 136.845 -190.235 ;
        RECT 136.515 -191.925 136.845 -191.595 ;
        RECT 136.515 -193.285 136.845 -192.955 ;
        RECT 136.515 -194.645 136.845 -194.315 ;
        RECT 136.515 -196.005 136.845 -195.675 ;
        RECT 136.515 -197.365 136.845 -197.035 ;
        RECT 136.515 -198.725 136.845 -198.395 ;
        RECT 136.515 -200.085 136.845 -199.755 ;
        RECT 136.515 -201.445 136.845 -201.115 ;
        RECT 136.515 -202.805 136.845 -202.475 ;
        RECT 136.515 -204.165 136.845 -203.835 ;
        RECT 136.515 -205.525 136.845 -205.195 ;
        RECT 136.515 -206.885 136.845 -206.555 ;
        RECT 136.515 -208.245 136.845 -207.915 ;
        RECT 136.515 -209.605 136.845 -209.275 ;
        RECT 136.515 -210.965 136.845 -210.635 ;
        RECT 136.515 -212.325 136.845 -211.995 ;
        RECT 136.515 -213.685 136.845 -213.355 ;
        RECT 136.515 -215.045 136.845 -214.715 ;
        RECT 136.515 -216.405 136.845 -216.075 ;
        RECT 136.515 -217.765 136.845 -217.435 ;
        RECT 136.515 -219.125 136.845 -218.795 ;
        RECT 136.515 -221.37 136.845 -220.24 ;
        RECT 136.52 -221.485 136.84 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.51 -121.535 137.84 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.875 129.8 138.205 130.93 ;
        RECT 137.875 127.675 138.205 128.005 ;
        RECT 137.875 126.315 138.205 126.645 ;
        RECT 137.875 124.955 138.205 125.285 ;
        RECT 137.875 123.595 138.205 123.925 ;
        RECT 137.88 123.595 138.2 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.235 129.8 139.565 130.93 ;
        RECT 139.235 127.675 139.565 128.005 ;
        RECT 139.235 126.315 139.565 126.645 ;
        RECT 139.235 124.955 139.565 125.285 ;
        RECT 139.235 123.595 139.565 123.925 ;
        RECT 139.24 123.595 139.56 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.235 -1.525 139.565 -1.195 ;
        RECT 139.235 -2.885 139.565 -2.555 ;
        RECT 139.24 -3.56 139.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.595 129.8 140.925 130.93 ;
        RECT 140.595 127.675 140.925 128.005 ;
        RECT 140.595 126.315 140.925 126.645 ;
        RECT 140.595 124.955 140.925 125.285 ;
        RECT 140.595 123.595 140.925 123.925 ;
        RECT 140.6 123.595 140.92 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.595 -1.525 140.925 -1.195 ;
        RECT 140.595 -2.885 140.925 -2.555 ;
        RECT 140.6 -3.56 140.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.595 -118.485 140.925 -118.155 ;
        RECT 140.595 -119.845 140.925 -119.515 ;
        RECT 140.595 -121.205 140.925 -120.875 ;
        RECT 140.595 -122.565 140.925 -122.235 ;
        RECT 140.595 -123.925 140.925 -123.595 ;
        RECT 140.595 -125.285 140.925 -124.955 ;
        RECT 140.595 -126.645 140.925 -126.315 ;
        RECT 140.595 -128.005 140.925 -127.675 ;
        RECT 140.595 -129.365 140.925 -129.035 ;
        RECT 140.595 -130.725 140.925 -130.395 ;
        RECT 140.595 -132.085 140.925 -131.755 ;
        RECT 140.595 -133.445 140.925 -133.115 ;
        RECT 140.595 -134.805 140.925 -134.475 ;
        RECT 140.595 -136.165 140.925 -135.835 ;
        RECT 140.595 -137.525 140.925 -137.195 ;
        RECT 140.595 -138.885 140.925 -138.555 ;
        RECT 140.595 -140.245 140.925 -139.915 ;
        RECT 140.595 -141.605 140.925 -141.275 ;
        RECT 140.595 -142.965 140.925 -142.635 ;
        RECT 140.595 -144.325 140.925 -143.995 ;
        RECT 140.595 -145.685 140.925 -145.355 ;
        RECT 140.595 -147.045 140.925 -146.715 ;
        RECT 140.595 -148.405 140.925 -148.075 ;
        RECT 140.595 -149.765 140.925 -149.435 ;
        RECT 140.595 -151.125 140.925 -150.795 ;
        RECT 140.595 -152.485 140.925 -152.155 ;
        RECT 140.595 -153.845 140.925 -153.515 ;
        RECT 140.595 -155.205 140.925 -154.875 ;
        RECT 140.595 -156.565 140.925 -156.235 ;
        RECT 140.595 -157.925 140.925 -157.595 ;
        RECT 140.595 -159.285 140.925 -158.955 ;
        RECT 140.595 -160.645 140.925 -160.315 ;
        RECT 140.595 -162.005 140.925 -161.675 ;
        RECT 140.595 -163.365 140.925 -163.035 ;
        RECT 140.595 -164.725 140.925 -164.395 ;
        RECT 140.595 -166.085 140.925 -165.755 ;
        RECT 140.595 -167.445 140.925 -167.115 ;
        RECT 140.595 -168.805 140.925 -168.475 ;
        RECT 140.595 -170.165 140.925 -169.835 ;
        RECT 140.595 -171.525 140.925 -171.195 ;
        RECT 140.595 -172.885 140.925 -172.555 ;
        RECT 140.595 -174.245 140.925 -173.915 ;
        RECT 140.595 -175.605 140.925 -175.275 ;
        RECT 140.595 -176.965 140.925 -176.635 ;
        RECT 140.595 -178.325 140.925 -177.995 ;
        RECT 140.595 -179.685 140.925 -179.355 ;
        RECT 140.595 -181.045 140.925 -180.715 ;
        RECT 140.595 -182.405 140.925 -182.075 ;
        RECT 140.595 -183.765 140.925 -183.435 ;
        RECT 140.595 -185.125 140.925 -184.795 ;
        RECT 140.595 -186.485 140.925 -186.155 ;
        RECT 140.595 -187.845 140.925 -187.515 ;
        RECT 140.595 -189.205 140.925 -188.875 ;
        RECT 140.595 -190.565 140.925 -190.235 ;
        RECT 140.595 -191.925 140.925 -191.595 ;
        RECT 140.595 -193.285 140.925 -192.955 ;
        RECT 140.595 -194.645 140.925 -194.315 ;
        RECT 140.595 -196.005 140.925 -195.675 ;
        RECT 140.595 -197.365 140.925 -197.035 ;
        RECT 140.595 -198.725 140.925 -198.395 ;
        RECT 140.595 -200.085 140.925 -199.755 ;
        RECT 140.595 -201.445 140.925 -201.115 ;
        RECT 140.595 -202.805 140.925 -202.475 ;
        RECT 140.595 -204.165 140.925 -203.835 ;
        RECT 140.595 -205.525 140.925 -205.195 ;
        RECT 140.595 -206.885 140.925 -206.555 ;
        RECT 140.595 -208.245 140.925 -207.915 ;
        RECT 140.595 -209.605 140.925 -209.275 ;
        RECT 140.595 -210.965 140.925 -210.635 ;
        RECT 140.595 -212.325 140.925 -211.995 ;
        RECT 140.595 -213.685 140.925 -213.355 ;
        RECT 140.595 -215.045 140.925 -214.715 ;
        RECT 140.595 -216.405 140.925 -216.075 ;
        RECT 140.595 -217.765 140.925 -217.435 ;
        RECT 140.595 -219.125 140.925 -218.795 ;
        RECT 140.595 -221.37 140.925 -220.24 ;
        RECT 140.6 -221.485 140.92 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.955 129.8 142.285 130.93 ;
        RECT 141.955 127.675 142.285 128.005 ;
        RECT 141.955 126.315 142.285 126.645 ;
        RECT 141.955 124.955 142.285 125.285 ;
        RECT 141.955 123.595 142.285 123.925 ;
        RECT 141.96 123.595 142.28 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.955 -1.525 142.285 -1.195 ;
        RECT 141.955 -2.885 142.285 -2.555 ;
        RECT 141.96 -3.56 142.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.955 -118.485 142.285 -118.155 ;
        RECT 141.955 -119.845 142.285 -119.515 ;
        RECT 141.955 -121.205 142.285 -120.875 ;
        RECT 141.955 -122.565 142.285 -122.235 ;
        RECT 141.955 -123.925 142.285 -123.595 ;
        RECT 141.955 -125.285 142.285 -124.955 ;
        RECT 141.955 -126.645 142.285 -126.315 ;
        RECT 141.955 -128.005 142.285 -127.675 ;
        RECT 141.955 -129.365 142.285 -129.035 ;
        RECT 141.955 -130.725 142.285 -130.395 ;
        RECT 141.955 -132.085 142.285 -131.755 ;
        RECT 141.955 -133.445 142.285 -133.115 ;
        RECT 141.955 -134.805 142.285 -134.475 ;
        RECT 141.955 -136.165 142.285 -135.835 ;
        RECT 141.955 -137.525 142.285 -137.195 ;
        RECT 141.955 -138.885 142.285 -138.555 ;
        RECT 141.955 -140.245 142.285 -139.915 ;
        RECT 141.955 -141.605 142.285 -141.275 ;
        RECT 141.955 -142.965 142.285 -142.635 ;
        RECT 141.955 -144.325 142.285 -143.995 ;
        RECT 141.955 -145.685 142.285 -145.355 ;
        RECT 141.955 -147.045 142.285 -146.715 ;
        RECT 141.955 -148.405 142.285 -148.075 ;
        RECT 141.955 -149.765 142.285 -149.435 ;
        RECT 141.955 -151.125 142.285 -150.795 ;
        RECT 141.955 -152.485 142.285 -152.155 ;
        RECT 141.955 -153.845 142.285 -153.515 ;
        RECT 141.955 -155.205 142.285 -154.875 ;
        RECT 141.955 -156.565 142.285 -156.235 ;
        RECT 141.955 -157.925 142.285 -157.595 ;
        RECT 141.955 -159.285 142.285 -158.955 ;
        RECT 141.955 -160.645 142.285 -160.315 ;
        RECT 141.955 -162.005 142.285 -161.675 ;
        RECT 141.955 -163.365 142.285 -163.035 ;
        RECT 141.955 -164.725 142.285 -164.395 ;
        RECT 141.955 -166.085 142.285 -165.755 ;
        RECT 141.955 -167.445 142.285 -167.115 ;
        RECT 141.955 -168.805 142.285 -168.475 ;
        RECT 141.955 -170.165 142.285 -169.835 ;
        RECT 141.955 -171.525 142.285 -171.195 ;
        RECT 141.955 -172.885 142.285 -172.555 ;
        RECT 141.955 -174.245 142.285 -173.915 ;
        RECT 141.955 -175.605 142.285 -175.275 ;
        RECT 141.955 -176.965 142.285 -176.635 ;
        RECT 141.955 -178.325 142.285 -177.995 ;
        RECT 141.955 -179.685 142.285 -179.355 ;
        RECT 141.955 -181.045 142.285 -180.715 ;
        RECT 141.955 -182.405 142.285 -182.075 ;
        RECT 141.955 -183.765 142.285 -183.435 ;
        RECT 141.955 -185.125 142.285 -184.795 ;
        RECT 141.955 -186.485 142.285 -186.155 ;
        RECT 141.955 -187.845 142.285 -187.515 ;
        RECT 141.955 -189.205 142.285 -188.875 ;
        RECT 141.955 -190.565 142.285 -190.235 ;
        RECT 141.955 -191.925 142.285 -191.595 ;
        RECT 141.955 -193.285 142.285 -192.955 ;
        RECT 141.955 -194.645 142.285 -194.315 ;
        RECT 141.955 -196.005 142.285 -195.675 ;
        RECT 141.955 -197.365 142.285 -197.035 ;
        RECT 141.955 -198.725 142.285 -198.395 ;
        RECT 141.955 -200.085 142.285 -199.755 ;
        RECT 141.955 -201.445 142.285 -201.115 ;
        RECT 141.955 -202.805 142.285 -202.475 ;
        RECT 141.955 -204.165 142.285 -203.835 ;
        RECT 141.955 -205.525 142.285 -205.195 ;
        RECT 141.955 -206.885 142.285 -206.555 ;
        RECT 141.955 -208.245 142.285 -207.915 ;
        RECT 141.955 -209.605 142.285 -209.275 ;
        RECT 141.955 -210.965 142.285 -210.635 ;
        RECT 141.955 -212.325 142.285 -211.995 ;
        RECT 141.955 -213.685 142.285 -213.355 ;
        RECT 141.955 -215.045 142.285 -214.715 ;
        RECT 141.955 -216.405 142.285 -216.075 ;
        RECT 141.955 -217.765 142.285 -217.435 ;
        RECT 141.955 -219.125 142.285 -218.795 ;
        RECT 141.955 -221.37 142.285 -220.24 ;
        RECT 141.96 -221.485 142.28 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.315 129.8 143.645 130.93 ;
        RECT 143.315 127.675 143.645 128.005 ;
        RECT 143.315 126.315 143.645 126.645 ;
        RECT 143.315 124.955 143.645 125.285 ;
        RECT 143.315 123.595 143.645 123.925 ;
        RECT 143.32 123.595 143.64 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.315 -122.565 143.645 -122.235 ;
        RECT 143.315 -123.925 143.645 -123.595 ;
        RECT 143.315 -125.285 143.645 -124.955 ;
        RECT 143.315 -126.645 143.645 -126.315 ;
        RECT 143.315 -128.005 143.645 -127.675 ;
        RECT 143.315 -129.365 143.645 -129.035 ;
        RECT 143.315 -130.725 143.645 -130.395 ;
        RECT 143.315 -132.085 143.645 -131.755 ;
        RECT 143.315 -133.445 143.645 -133.115 ;
        RECT 143.315 -134.805 143.645 -134.475 ;
        RECT 143.315 -136.165 143.645 -135.835 ;
        RECT 143.315 -137.525 143.645 -137.195 ;
        RECT 143.315 -138.885 143.645 -138.555 ;
        RECT 143.315 -140.245 143.645 -139.915 ;
        RECT 143.315 -141.605 143.645 -141.275 ;
        RECT 143.315 -142.965 143.645 -142.635 ;
        RECT 143.315 -144.325 143.645 -143.995 ;
        RECT 143.315 -145.685 143.645 -145.355 ;
        RECT 143.315 -147.045 143.645 -146.715 ;
        RECT 143.315 -148.405 143.645 -148.075 ;
        RECT 143.315 -149.765 143.645 -149.435 ;
        RECT 143.315 -151.125 143.645 -150.795 ;
        RECT 143.315 -152.485 143.645 -152.155 ;
        RECT 143.315 -153.845 143.645 -153.515 ;
        RECT 143.315 -155.205 143.645 -154.875 ;
        RECT 143.315 -156.565 143.645 -156.235 ;
        RECT 143.315 -157.925 143.645 -157.595 ;
        RECT 143.315 -159.285 143.645 -158.955 ;
        RECT 143.315 -160.645 143.645 -160.315 ;
        RECT 143.315 -162.005 143.645 -161.675 ;
        RECT 143.315 -163.365 143.645 -163.035 ;
        RECT 143.315 -164.725 143.645 -164.395 ;
        RECT 143.315 -166.085 143.645 -165.755 ;
        RECT 143.315 -167.445 143.645 -167.115 ;
        RECT 143.315 -168.805 143.645 -168.475 ;
        RECT 143.315 -170.165 143.645 -169.835 ;
        RECT 143.315 -171.525 143.645 -171.195 ;
        RECT 143.315 -172.885 143.645 -172.555 ;
        RECT 143.315 -174.245 143.645 -173.915 ;
        RECT 143.315 -175.605 143.645 -175.275 ;
        RECT 143.315 -176.965 143.645 -176.635 ;
        RECT 143.315 -178.325 143.645 -177.995 ;
        RECT 143.315 -179.685 143.645 -179.355 ;
        RECT 143.315 -181.045 143.645 -180.715 ;
        RECT 143.315 -182.405 143.645 -182.075 ;
        RECT 143.315 -183.765 143.645 -183.435 ;
        RECT 143.315 -185.125 143.645 -184.795 ;
        RECT 143.315 -186.485 143.645 -186.155 ;
        RECT 143.315 -187.845 143.645 -187.515 ;
        RECT 143.315 -189.205 143.645 -188.875 ;
        RECT 143.315 -190.565 143.645 -190.235 ;
        RECT 143.315 -191.925 143.645 -191.595 ;
        RECT 143.315 -193.285 143.645 -192.955 ;
        RECT 143.315 -194.645 143.645 -194.315 ;
        RECT 143.315 -196.005 143.645 -195.675 ;
        RECT 143.315 -197.365 143.645 -197.035 ;
        RECT 143.315 -198.725 143.645 -198.395 ;
        RECT 143.315 -200.085 143.645 -199.755 ;
        RECT 143.315 -201.445 143.645 -201.115 ;
        RECT 143.315 -202.805 143.645 -202.475 ;
        RECT 143.315 -204.165 143.645 -203.835 ;
        RECT 143.315 -205.525 143.645 -205.195 ;
        RECT 143.315 -206.885 143.645 -206.555 ;
        RECT 143.315 -208.245 143.645 -207.915 ;
        RECT 143.315 -209.605 143.645 -209.275 ;
        RECT 143.315 -210.965 143.645 -210.635 ;
        RECT 143.315 -212.325 143.645 -211.995 ;
        RECT 143.315 -213.685 143.645 -213.355 ;
        RECT 143.315 -215.045 143.645 -214.715 ;
        RECT 143.315 -216.405 143.645 -216.075 ;
        RECT 143.315 -217.765 143.645 -217.435 ;
        RECT 143.315 -219.125 143.645 -218.795 ;
        RECT 143.315 -221.37 143.645 -220.24 ;
        RECT 143.32 -221.485 143.64 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.61 -121.535 143.94 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.675 129.8 145.005 130.93 ;
        RECT 144.675 127.675 145.005 128.005 ;
        RECT 144.675 126.315 145.005 126.645 ;
        RECT 144.675 124.955 145.005 125.285 ;
        RECT 144.675 123.595 145.005 123.925 ;
        RECT 144.68 123.595 145 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.675 -1.525 145.005 -1.195 ;
        RECT 144.675 -2.885 145.005 -2.555 ;
        RECT 144.68 -3.56 145 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.035 129.8 146.365 130.93 ;
        RECT 146.035 127.675 146.365 128.005 ;
        RECT 146.035 126.315 146.365 126.645 ;
        RECT 146.035 124.955 146.365 125.285 ;
        RECT 146.035 123.595 146.365 123.925 ;
        RECT 146.04 123.595 146.36 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.035 -1.525 146.365 -1.195 ;
        RECT 146.035 -2.885 146.365 -2.555 ;
        RECT 146.04 -3.56 146.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.395 129.8 147.725 130.93 ;
        RECT 147.395 127.675 147.725 128.005 ;
        RECT 147.395 126.315 147.725 126.645 ;
        RECT 147.395 124.955 147.725 125.285 ;
        RECT 147.395 123.595 147.725 123.925 ;
        RECT 147.4 123.595 147.72 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.395 -1.525 147.725 -1.195 ;
        RECT 147.395 -2.885 147.725 -2.555 ;
        RECT 147.4 -3.56 147.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.395 -118.485 147.725 -118.155 ;
        RECT 147.395 -119.845 147.725 -119.515 ;
        RECT 147.395 -121.205 147.725 -120.875 ;
        RECT 147.395 -122.565 147.725 -122.235 ;
        RECT 147.395 -123.925 147.725 -123.595 ;
        RECT 147.395 -125.285 147.725 -124.955 ;
        RECT 147.395 -126.645 147.725 -126.315 ;
        RECT 147.395 -128.005 147.725 -127.675 ;
        RECT 147.395 -129.365 147.725 -129.035 ;
        RECT 147.395 -130.725 147.725 -130.395 ;
        RECT 147.395 -132.085 147.725 -131.755 ;
        RECT 147.395 -133.445 147.725 -133.115 ;
        RECT 147.395 -134.805 147.725 -134.475 ;
        RECT 147.395 -136.165 147.725 -135.835 ;
        RECT 147.395 -137.525 147.725 -137.195 ;
        RECT 147.395 -138.885 147.725 -138.555 ;
        RECT 147.395 -140.245 147.725 -139.915 ;
        RECT 147.395 -141.605 147.725 -141.275 ;
        RECT 147.395 -142.965 147.725 -142.635 ;
        RECT 147.395 -144.325 147.725 -143.995 ;
        RECT 147.395 -145.685 147.725 -145.355 ;
        RECT 147.395 -147.045 147.725 -146.715 ;
        RECT 147.395 -148.405 147.725 -148.075 ;
        RECT 147.395 -149.765 147.725 -149.435 ;
        RECT 147.395 -151.125 147.725 -150.795 ;
        RECT 147.395 -152.485 147.725 -152.155 ;
        RECT 147.395 -153.845 147.725 -153.515 ;
        RECT 147.395 -155.205 147.725 -154.875 ;
        RECT 147.395 -156.565 147.725 -156.235 ;
        RECT 147.395 -157.925 147.725 -157.595 ;
        RECT 147.395 -159.285 147.725 -158.955 ;
        RECT 147.395 -160.645 147.725 -160.315 ;
        RECT 147.395 -162.005 147.725 -161.675 ;
        RECT 147.395 -163.365 147.725 -163.035 ;
        RECT 147.395 -164.725 147.725 -164.395 ;
        RECT 147.395 -166.085 147.725 -165.755 ;
        RECT 147.395 -167.445 147.725 -167.115 ;
        RECT 147.395 -168.805 147.725 -168.475 ;
        RECT 147.395 -170.165 147.725 -169.835 ;
        RECT 147.395 -171.525 147.725 -171.195 ;
        RECT 147.395 -172.885 147.725 -172.555 ;
        RECT 147.395 -174.245 147.725 -173.915 ;
        RECT 147.395 -175.605 147.725 -175.275 ;
        RECT 147.395 -176.965 147.725 -176.635 ;
        RECT 147.395 -178.325 147.725 -177.995 ;
        RECT 147.395 -179.685 147.725 -179.355 ;
        RECT 147.395 -181.045 147.725 -180.715 ;
        RECT 147.395 -182.405 147.725 -182.075 ;
        RECT 147.395 -183.765 147.725 -183.435 ;
        RECT 147.395 -185.125 147.725 -184.795 ;
        RECT 147.395 -186.485 147.725 -186.155 ;
        RECT 147.395 -187.845 147.725 -187.515 ;
        RECT 147.395 -189.205 147.725 -188.875 ;
        RECT 147.395 -190.565 147.725 -190.235 ;
        RECT 147.395 -191.925 147.725 -191.595 ;
        RECT 147.395 -193.285 147.725 -192.955 ;
        RECT 147.395 -194.645 147.725 -194.315 ;
        RECT 147.395 -196.005 147.725 -195.675 ;
        RECT 147.395 -197.365 147.725 -197.035 ;
        RECT 147.395 -198.725 147.725 -198.395 ;
        RECT 147.395 -200.085 147.725 -199.755 ;
        RECT 147.395 -201.445 147.725 -201.115 ;
        RECT 147.395 -202.805 147.725 -202.475 ;
        RECT 147.395 -204.165 147.725 -203.835 ;
        RECT 147.395 -205.525 147.725 -205.195 ;
        RECT 147.395 -206.885 147.725 -206.555 ;
        RECT 147.395 -208.245 147.725 -207.915 ;
        RECT 147.395 -209.605 147.725 -209.275 ;
        RECT 147.395 -210.965 147.725 -210.635 ;
        RECT 147.395 -212.325 147.725 -211.995 ;
        RECT 147.395 -213.685 147.725 -213.355 ;
        RECT 147.395 -215.045 147.725 -214.715 ;
        RECT 147.395 -216.405 147.725 -216.075 ;
        RECT 147.395 -217.765 147.725 -217.435 ;
        RECT 147.395 -219.125 147.725 -218.795 ;
        RECT 147.395 -221.37 147.725 -220.24 ;
        RECT 147.4 -221.485 147.72 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.755 129.8 149.085 130.93 ;
        RECT 148.755 127.675 149.085 128.005 ;
        RECT 148.755 126.315 149.085 126.645 ;
        RECT 148.755 124.955 149.085 125.285 ;
        RECT 148.755 123.595 149.085 123.925 ;
        RECT 148.76 123.595 149.08 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.755 -122.565 149.085 -122.235 ;
        RECT 148.755 -123.925 149.085 -123.595 ;
        RECT 148.755 -125.285 149.085 -124.955 ;
        RECT 148.755 -126.645 149.085 -126.315 ;
        RECT 148.755 -128.005 149.085 -127.675 ;
        RECT 148.755 -129.365 149.085 -129.035 ;
        RECT 148.755 -130.725 149.085 -130.395 ;
        RECT 148.755 -132.085 149.085 -131.755 ;
        RECT 148.755 -133.445 149.085 -133.115 ;
        RECT 148.755 -134.805 149.085 -134.475 ;
        RECT 148.755 -136.165 149.085 -135.835 ;
        RECT 148.755 -137.525 149.085 -137.195 ;
        RECT 148.755 -138.885 149.085 -138.555 ;
        RECT 148.755 -140.245 149.085 -139.915 ;
        RECT 148.755 -141.605 149.085 -141.275 ;
        RECT 148.755 -142.965 149.085 -142.635 ;
        RECT 148.755 -144.325 149.085 -143.995 ;
        RECT 148.755 -145.685 149.085 -145.355 ;
        RECT 148.755 -147.045 149.085 -146.715 ;
        RECT 148.755 -148.405 149.085 -148.075 ;
        RECT 148.755 -149.765 149.085 -149.435 ;
        RECT 148.755 -151.125 149.085 -150.795 ;
        RECT 148.755 -152.485 149.085 -152.155 ;
        RECT 148.755 -153.845 149.085 -153.515 ;
        RECT 148.755 -155.205 149.085 -154.875 ;
        RECT 148.755 -156.565 149.085 -156.235 ;
        RECT 148.755 -157.925 149.085 -157.595 ;
        RECT 148.755 -159.285 149.085 -158.955 ;
        RECT 148.755 -160.645 149.085 -160.315 ;
        RECT 148.755 -162.005 149.085 -161.675 ;
        RECT 148.755 -163.365 149.085 -163.035 ;
        RECT 148.755 -164.725 149.085 -164.395 ;
        RECT 148.755 -166.085 149.085 -165.755 ;
        RECT 148.755 -167.445 149.085 -167.115 ;
        RECT 148.755 -168.805 149.085 -168.475 ;
        RECT 148.755 -170.165 149.085 -169.835 ;
        RECT 148.755 -171.525 149.085 -171.195 ;
        RECT 148.755 -172.885 149.085 -172.555 ;
        RECT 148.755 -174.245 149.085 -173.915 ;
        RECT 148.755 -175.605 149.085 -175.275 ;
        RECT 148.755 -176.965 149.085 -176.635 ;
        RECT 148.755 -178.325 149.085 -177.995 ;
        RECT 148.755 -179.685 149.085 -179.355 ;
        RECT 148.755 -181.045 149.085 -180.715 ;
        RECT 148.755 -182.405 149.085 -182.075 ;
        RECT 148.755 -183.765 149.085 -183.435 ;
        RECT 148.755 -185.125 149.085 -184.795 ;
        RECT 148.755 -186.485 149.085 -186.155 ;
        RECT 148.755 -187.845 149.085 -187.515 ;
        RECT 148.755 -189.205 149.085 -188.875 ;
        RECT 148.755 -190.565 149.085 -190.235 ;
        RECT 148.755 -191.925 149.085 -191.595 ;
        RECT 148.755 -193.285 149.085 -192.955 ;
        RECT 148.755 -194.645 149.085 -194.315 ;
        RECT 148.755 -196.005 149.085 -195.675 ;
        RECT 148.755 -197.365 149.085 -197.035 ;
        RECT 148.755 -198.725 149.085 -198.395 ;
        RECT 148.755 -200.085 149.085 -199.755 ;
        RECT 148.755 -201.445 149.085 -201.115 ;
        RECT 148.755 -202.805 149.085 -202.475 ;
        RECT 148.755 -204.165 149.085 -203.835 ;
        RECT 148.755 -205.525 149.085 -205.195 ;
        RECT 148.755 -206.885 149.085 -206.555 ;
        RECT 148.755 -208.245 149.085 -207.915 ;
        RECT 148.755 -209.605 149.085 -209.275 ;
        RECT 148.755 -210.965 149.085 -210.635 ;
        RECT 148.755 -212.325 149.085 -211.995 ;
        RECT 148.755 -213.685 149.085 -213.355 ;
        RECT 148.755 -215.045 149.085 -214.715 ;
        RECT 148.755 -216.405 149.085 -216.075 ;
        RECT 148.755 -217.765 149.085 -217.435 ;
        RECT 148.755 -219.125 149.085 -218.795 ;
        RECT 148.755 -221.37 149.085 -220.24 ;
        RECT 148.76 -221.485 149.08 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.71 -121.535 150.04 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.115 129.8 150.445 130.93 ;
        RECT 150.115 127.675 150.445 128.005 ;
        RECT 150.115 126.315 150.445 126.645 ;
        RECT 150.115 124.955 150.445 125.285 ;
        RECT 150.115 123.595 150.445 123.925 ;
        RECT 150.12 123.595 150.44 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.475 129.8 151.805 130.93 ;
        RECT 151.475 127.675 151.805 128.005 ;
        RECT 151.475 126.315 151.805 126.645 ;
        RECT 151.475 124.955 151.805 125.285 ;
        RECT 151.475 123.595 151.805 123.925 ;
        RECT 151.48 123.595 151.8 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.475 -1.525 151.805 -1.195 ;
        RECT 151.475 -2.885 151.805 -2.555 ;
        RECT 151.48 -3.56 151.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.835 129.8 153.165 130.93 ;
        RECT 152.835 127.675 153.165 128.005 ;
        RECT 152.835 126.315 153.165 126.645 ;
        RECT 152.835 124.955 153.165 125.285 ;
        RECT 152.835 123.595 153.165 123.925 ;
        RECT 152.84 123.595 153.16 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.835 -1.525 153.165 -1.195 ;
        RECT 152.835 -2.885 153.165 -2.555 ;
        RECT 152.84 -3.56 153.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.195 129.8 154.525 130.93 ;
        RECT 154.195 127.675 154.525 128.005 ;
        RECT 154.195 126.315 154.525 126.645 ;
        RECT 154.195 124.955 154.525 125.285 ;
        RECT 154.195 123.595 154.525 123.925 ;
        RECT 154.2 123.595 154.52 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.195 -1.525 154.525 -1.195 ;
        RECT 154.195 -2.885 154.525 -2.555 ;
        RECT 154.2 -3.56 154.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.195 -118.485 154.525 -118.155 ;
        RECT 154.195 -119.845 154.525 -119.515 ;
        RECT 154.195 -121.205 154.525 -120.875 ;
        RECT 154.195 -122.565 154.525 -122.235 ;
        RECT 154.195 -123.925 154.525 -123.595 ;
        RECT 154.195 -125.285 154.525 -124.955 ;
        RECT 154.195 -126.645 154.525 -126.315 ;
        RECT 154.195 -128.005 154.525 -127.675 ;
        RECT 154.195 -129.365 154.525 -129.035 ;
        RECT 154.195 -130.725 154.525 -130.395 ;
        RECT 154.195 -132.085 154.525 -131.755 ;
        RECT 154.195 -133.445 154.525 -133.115 ;
        RECT 154.195 -134.805 154.525 -134.475 ;
        RECT 154.195 -136.165 154.525 -135.835 ;
        RECT 154.195 -137.525 154.525 -137.195 ;
        RECT 154.195 -138.885 154.525 -138.555 ;
        RECT 154.195 -140.245 154.525 -139.915 ;
        RECT 154.195 -141.605 154.525 -141.275 ;
        RECT 154.195 -142.965 154.525 -142.635 ;
        RECT 154.195 -144.325 154.525 -143.995 ;
        RECT 154.195 -145.685 154.525 -145.355 ;
        RECT 154.195 -147.045 154.525 -146.715 ;
        RECT 154.195 -148.405 154.525 -148.075 ;
        RECT 154.195 -149.765 154.525 -149.435 ;
        RECT 154.195 -151.125 154.525 -150.795 ;
        RECT 154.195 -152.485 154.525 -152.155 ;
        RECT 154.195 -153.845 154.525 -153.515 ;
        RECT 154.195 -155.205 154.525 -154.875 ;
        RECT 154.195 -156.565 154.525 -156.235 ;
        RECT 154.195 -157.925 154.525 -157.595 ;
        RECT 154.195 -159.285 154.525 -158.955 ;
        RECT 154.195 -160.645 154.525 -160.315 ;
        RECT 154.195 -162.005 154.525 -161.675 ;
        RECT 154.195 -163.365 154.525 -163.035 ;
        RECT 154.195 -164.725 154.525 -164.395 ;
        RECT 154.195 -166.085 154.525 -165.755 ;
        RECT 154.195 -167.445 154.525 -167.115 ;
        RECT 154.195 -168.805 154.525 -168.475 ;
        RECT 154.195 -170.165 154.525 -169.835 ;
        RECT 154.195 -171.525 154.525 -171.195 ;
        RECT 154.195 -172.885 154.525 -172.555 ;
        RECT 154.195 -174.245 154.525 -173.915 ;
        RECT 154.195 -175.605 154.525 -175.275 ;
        RECT 154.195 -176.965 154.525 -176.635 ;
        RECT 154.195 -178.325 154.525 -177.995 ;
        RECT 154.195 -179.685 154.525 -179.355 ;
        RECT 154.195 -181.045 154.525 -180.715 ;
        RECT 154.195 -182.405 154.525 -182.075 ;
        RECT 154.195 -183.765 154.525 -183.435 ;
        RECT 154.195 -185.125 154.525 -184.795 ;
        RECT 154.195 -186.485 154.525 -186.155 ;
        RECT 154.195 -187.845 154.525 -187.515 ;
        RECT 154.195 -189.205 154.525 -188.875 ;
        RECT 154.195 -190.565 154.525 -190.235 ;
        RECT 154.195 -191.925 154.525 -191.595 ;
        RECT 154.195 -193.285 154.525 -192.955 ;
        RECT 154.195 -194.645 154.525 -194.315 ;
        RECT 154.195 -196.005 154.525 -195.675 ;
        RECT 154.195 -197.365 154.525 -197.035 ;
        RECT 154.195 -198.725 154.525 -198.395 ;
        RECT 154.195 -200.085 154.525 -199.755 ;
        RECT 154.195 -201.445 154.525 -201.115 ;
        RECT 154.195 -202.805 154.525 -202.475 ;
        RECT 154.195 -204.165 154.525 -203.835 ;
        RECT 154.195 -205.525 154.525 -205.195 ;
        RECT 154.195 -206.885 154.525 -206.555 ;
        RECT 154.195 -208.245 154.525 -207.915 ;
        RECT 154.195 -209.605 154.525 -209.275 ;
        RECT 154.195 -210.965 154.525 -210.635 ;
        RECT 154.195 -212.325 154.525 -211.995 ;
        RECT 154.195 -213.685 154.525 -213.355 ;
        RECT 154.195 -215.045 154.525 -214.715 ;
        RECT 154.195 -216.405 154.525 -216.075 ;
        RECT 154.195 -217.765 154.525 -217.435 ;
        RECT 154.195 -219.125 154.525 -218.795 ;
        RECT 154.195 -221.37 154.525 -220.24 ;
        RECT 154.2 -221.485 154.52 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.555 129.8 155.885 130.93 ;
        RECT 155.555 127.675 155.885 128.005 ;
        RECT 155.555 126.315 155.885 126.645 ;
        RECT 155.555 124.955 155.885 125.285 ;
        RECT 155.555 123.595 155.885 123.925 ;
        RECT 155.56 123.595 155.88 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.555 -122.565 155.885 -122.235 ;
        RECT 155.555 -123.925 155.885 -123.595 ;
        RECT 155.555 -125.285 155.885 -124.955 ;
        RECT 155.555 -126.645 155.885 -126.315 ;
        RECT 155.555 -128.005 155.885 -127.675 ;
        RECT 155.555 -129.365 155.885 -129.035 ;
        RECT 155.555 -130.725 155.885 -130.395 ;
        RECT 155.555 -132.085 155.885 -131.755 ;
        RECT 155.555 -133.445 155.885 -133.115 ;
        RECT 155.555 -134.805 155.885 -134.475 ;
        RECT 155.555 -136.165 155.885 -135.835 ;
        RECT 155.555 -137.525 155.885 -137.195 ;
        RECT 155.555 -138.885 155.885 -138.555 ;
        RECT 155.555 -140.245 155.885 -139.915 ;
        RECT 155.555 -141.605 155.885 -141.275 ;
        RECT 155.555 -142.965 155.885 -142.635 ;
        RECT 155.555 -144.325 155.885 -143.995 ;
        RECT 155.555 -145.685 155.885 -145.355 ;
        RECT 155.555 -147.045 155.885 -146.715 ;
        RECT 155.555 -148.405 155.885 -148.075 ;
        RECT 155.555 -149.765 155.885 -149.435 ;
        RECT 155.555 -151.125 155.885 -150.795 ;
        RECT 155.555 -152.485 155.885 -152.155 ;
        RECT 155.555 -153.845 155.885 -153.515 ;
        RECT 155.555 -155.205 155.885 -154.875 ;
        RECT 155.555 -156.565 155.885 -156.235 ;
        RECT 155.555 -157.925 155.885 -157.595 ;
        RECT 155.555 -159.285 155.885 -158.955 ;
        RECT 155.555 -160.645 155.885 -160.315 ;
        RECT 155.555 -162.005 155.885 -161.675 ;
        RECT 155.555 -163.365 155.885 -163.035 ;
        RECT 155.555 -164.725 155.885 -164.395 ;
        RECT 155.555 -166.085 155.885 -165.755 ;
        RECT 155.555 -167.445 155.885 -167.115 ;
        RECT 155.555 -168.805 155.885 -168.475 ;
        RECT 155.555 -170.165 155.885 -169.835 ;
        RECT 155.555 -171.525 155.885 -171.195 ;
        RECT 155.555 -172.885 155.885 -172.555 ;
        RECT 155.555 -174.245 155.885 -173.915 ;
        RECT 155.555 -175.605 155.885 -175.275 ;
        RECT 155.555 -176.965 155.885 -176.635 ;
        RECT 155.555 -178.325 155.885 -177.995 ;
        RECT 155.555 -179.685 155.885 -179.355 ;
        RECT 155.555 -181.045 155.885 -180.715 ;
        RECT 155.555 -182.405 155.885 -182.075 ;
        RECT 155.555 -183.765 155.885 -183.435 ;
        RECT 155.555 -185.125 155.885 -184.795 ;
        RECT 155.555 -186.485 155.885 -186.155 ;
        RECT 155.555 -187.845 155.885 -187.515 ;
        RECT 155.555 -189.205 155.885 -188.875 ;
        RECT 155.555 -190.565 155.885 -190.235 ;
        RECT 155.555 -191.925 155.885 -191.595 ;
        RECT 155.555 -193.285 155.885 -192.955 ;
        RECT 155.555 -194.645 155.885 -194.315 ;
        RECT 155.555 -196.005 155.885 -195.675 ;
        RECT 155.555 -197.365 155.885 -197.035 ;
        RECT 155.555 -198.725 155.885 -198.395 ;
        RECT 155.555 -200.085 155.885 -199.755 ;
        RECT 155.555 -201.445 155.885 -201.115 ;
        RECT 155.555 -202.805 155.885 -202.475 ;
        RECT 155.555 -204.165 155.885 -203.835 ;
        RECT 155.555 -205.525 155.885 -205.195 ;
        RECT 155.555 -206.885 155.885 -206.555 ;
        RECT 155.555 -208.245 155.885 -207.915 ;
        RECT 155.555 -209.605 155.885 -209.275 ;
        RECT 155.555 -210.965 155.885 -210.635 ;
        RECT 155.555 -212.325 155.885 -211.995 ;
        RECT 155.555 -213.685 155.885 -213.355 ;
        RECT 155.555 -215.045 155.885 -214.715 ;
        RECT 155.555 -216.405 155.885 -216.075 ;
        RECT 155.555 -217.765 155.885 -217.435 ;
        RECT 155.555 -219.125 155.885 -218.795 ;
        RECT 155.555 -221.37 155.885 -220.24 ;
        RECT 155.56 -221.485 155.88 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.81 -121.535 156.14 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.915 129.8 157.245 130.93 ;
        RECT 156.915 127.675 157.245 128.005 ;
        RECT 156.915 126.315 157.245 126.645 ;
        RECT 156.915 124.955 157.245 125.285 ;
        RECT 156.915 123.595 157.245 123.925 ;
        RECT 156.92 123.595 157.24 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.915 -1.525 157.245 -1.195 ;
        RECT 156.915 -2.885 157.245 -2.555 ;
        RECT 156.92 -3.56 157.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.275 129.8 158.605 130.93 ;
        RECT 158.275 127.675 158.605 128.005 ;
        RECT 158.275 126.315 158.605 126.645 ;
        RECT 158.275 124.955 158.605 125.285 ;
        RECT 158.275 123.595 158.605 123.925 ;
        RECT 158.28 123.595 158.6 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.275 -1.525 158.605 -1.195 ;
        RECT 158.275 -2.885 158.605 -2.555 ;
        RECT 158.28 -3.56 158.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.635 129.8 159.965 130.93 ;
        RECT 159.635 127.675 159.965 128.005 ;
        RECT 159.635 126.315 159.965 126.645 ;
        RECT 159.635 124.955 159.965 125.285 ;
        RECT 159.635 123.595 159.965 123.925 ;
        RECT 159.64 123.595 159.96 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.635 -1.525 159.965 -1.195 ;
        RECT 159.635 -2.885 159.965 -2.555 ;
        RECT 159.64 -3.56 159.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.635 -118.485 159.965 -118.155 ;
        RECT 159.635 -119.845 159.965 -119.515 ;
        RECT 159.635 -121.205 159.965 -120.875 ;
        RECT 159.635 -122.565 159.965 -122.235 ;
        RECT 159.635 -123.925 159.965 -123.595 ;
        RECT 159.635 -125.285 159.965 -124.955 ;
        RECT 159.635 -126.645 159.965 -126.315 ;
        RECT 159.635 -128.005 159.965 -127.675 ;
        RECT 159.635 -129.365 159.965 -129.035 ;
        RECT 159.635 -130.725 159.965 -130.395 ;
        RECT 159.635 -132.085 159.965 -131.755 ;
        RECT 159.635 -133.445 159.965 -133.115 ;
        RECT 159.635 -134.805 159.965 -134.475 ;
        RECT 159.635 -136.165 159.965 -135.835 ;
        RECT 159.635 -137.525 159.965 -137.195 ;
        RECT 159.635 -138.885 159.965 -138.555 ;
        RECT 159.635 -140.245 159.965 -139.915 ;
        RECT 159.635 -141.605 159.965 -141.275 ;
        RECT 159.635 -142.965 159.965 -142.635 ;
        RECT 159.635 -144.325 159.965 -143.995 ;
        RECT 159.635 -145.685 159.965 -145.355 ;
        RECT 159.635 -147.045 159.965 -146.715 ;
        RECT 159.635 -148.405 159.965 -148.075 ;
        RECT 159.635 -149.765 159.965 -149.435 ;
        RECT 159.635 -151.125 159.965 -150.795 ;
        RECT 159.635 -152.485 159.965 -152.155 ;
        RECT 159.635 -153.845 159.965 -153.515 ;
        RECT 159.635 -155.205 159.965 -154.875 ;
        RECT 159.635 -156.565 159.965 -156.235 ;
        RECT 159.635 -157.925 159.965 -157.595 ;
        RECT 159.635 -159.285 159.965 -158.955 ;
        RECT 159.635 -160.645 159.965 -160.315 ;
        RECT 159.635 -162.005 159.965 -161.675 ;
        RECT 159.635 -163.365 159.965 -163.035 ;
        RECT 159.635 -164.725 159.965 -164.395 ;
        RECT 159.635 -166.085 159.965 -165.755 ;
        RECT 159.635 -167.445 159.965 -167.115 ;
        RECT 159.635 -168.805 159.965 -168.475 ;
        RECT 159.635 -170.165 159.965 -169.835 ;
        RECT 159.635 -171.525 159.965 -171.195 ;
        RECT 159.635 -172.885 159.965 -172.555 ;
        RECT 159.635 -174.245 159.965 -173.915 ;
        RECT 159.635 -175.605 159.965 -175.275 ;
        RECT 159.635 -176.965 159.965 -176.635 ;
        RECT 159.635 -178.325 159.965 -177.995 ;
        RECT 159.635 -179.685 159.965 -179.355 ;
        RECT 159.635 -181.045 159.965 -180.715 ;
        RECT 159.635 -182.405 159.965 -182.075 ;
        RECT 159.635 -183.765 159.965 -183.435 ;
        RECT 159.635 -185.125 159.965 -184.795 ;
        RECT 159.635 -186.485 159.965 -186.155 ;
        RECT 159.635 -187.845 159.965 -187.515 ;
        RECT 159.635 -189.205 159.965 -188.875 ;
        RECT 159.635 -190.565 159.965 -190.235 ;
        RECT 159.635 -191.925 159.965 -191.595 ;
        RECT 159.635 -193.285 159.965 -192.955 ;
        RECT 159.635 -194.645 159.965 -194.315 ;
        RECT 159.635 -196.005 159.965 -195.675 ;
        RECT 159.635 -197.365 159.965 -197.035 ;
        RECT 159.635 -198.725 159.965 -198.395 ;
        RECT 159.635 -200.085 159.965 -199.755 ;
        RECT 159.635 -201.445 159.965 -201.115 ;
        RECT 159.635 -202.805 159.965 -202.475 ;
        RECT 159.635 -204.165 159.965 -203.835 ;
        RECT 159.635 -205.525 159.965 -205.195 ;
        RECT 159.635 -206.885 159.965 -206.555 ;
        RECT 159.635 -208.245 159.965 -207.915 ;
        RECT 159.635 -209.605 159.965 -209.275 ;
        RECT 159.635 -210.965 159.965 -210.635 ;
        RECT 159.635 -212.325 159.965 -211.995 ;
        RECT 159.635 -213.685 159.965 -213.355 ;
        RECT 159.635 -215.045 159.965 -214.715 ;
        RECT 159.635 -216.405 159.965 -216.075 ;
        RECT 159.635 -217.765 159.965 -217.435 ;
        RECT 159.635 -219.125 159.965 -218.795 ;
        RECT 159.635 -221.37 159.965 -220.24 ;
        RECT 159.64 -221.485 159.96 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.995 129.8 161.325 130.93 ;
        RECT 160.995 127.675 161.325 128.005 ;
        RECT 160.995 126.315 161.325 126.645 ;
        RECT 160.995 124.955 161.325 125.285 ;
        RECT 160.995 123.595 161.325 123.925 ;
        RECT 161 123.595 161.32 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.995 -122.565 161.325 -122.235 ;
        RECT 160.995 -123.925 161.325 -123.595 ;
        RECT 160.995 -125.285 161.325 -124.955 ;
        RECT 160.995 -126.645 161.325 -126.315 ;
        RECT 160.995 -128.005 161.325 -127.675 ;
        RECT 160.995 -129.365 161.325 -129.035 ;
        RECT 160.995 -130.725 161.325 -130.395 ;
        RECT 160.995 -132.085 161.325 -131.755 ;
        RECT 160.995 -133.445 161.325 -133.115 ;
        RECT 160.995 -134.805 161.325 -134.475 ;
        RECT 160.995 -136.165 161.325 -135.835 ;
        RECT 160.995 -137.525 161.325 -137.195 ;
        RECT 160.995 -138.885 161.325 -138.555 ;
        RECT 160.995 -140.245 161.325 -139.915 ;
        RECT 160.995 -141.605 161.325 -141.275 ;
        RECT 160.995 -142.965 161.325 -142.635 ;
        RECT 160.995 -144.325 161.325 -143.995 ;
        RECT 160.995 -145.685 161.325 -145.355 ;
        RECT 160.995 -147.045 161.325 -146.715 ;
        RECT 160.995 -148.405 161.325 -148.075 ;
        RECT 160.995 -149.765 161.325 -149.435 ;
        RECT 160.995 -151.125 161.325 -150.795 ;
        RECT 160.995 -152.485 161.325 -152.155 ;
        RECT 160.995 -153.845 161.325 -153.515 ;
        RECT 160.995 -155.205 161.325 -154.875 ;
        RECT 160.995 -156.565 161.325 -156.235 ;
        RECT 160.995 -157.925 161.325 -157.595 ;
        RECT 160.995 -159.285 161.325 -158.955 ;
        RECT 160.995 -160.645 161.325 -160.315 ;
        RECT 160.995 -162.005 161.325 -161.675 ;
        RECT 160.995 -163.365 161.325 -163.035 ;
        RECT 160.995 -164.725 161.325 -164.395 ;
        RECT 160.995 -166.085 161.325 -165.755 ;
        RECT 160.995 -167.445 161.325 -167.115 ;
        RECT 160.995 -168.805 161.325 -168.475 ;
        RECT 160.995 -170.165 161.325 -169.835 ;
        RECT 160.995 -171.525 161.325 -171.195 ;
        RECT 160.995 -172.885 161.325 -172.555 ;
        RECT 160.995 -174.245 161.325 -173.915 ;
        RECT 160.995 -175.605 161.325 -175.275 ;
        RECT 160.995 -176.965 161.325 -176.635 ;
        RECT 160.995 -178.325 161.325 -177.995 ;
        RECT 160.995 -179.685 161.325 -179.355 ;
        RECT 160.995 -181.045 161.325 -180.715 ;
        RECT 160.995 -182.405 161.325 -182.075 ;
        RECT 160.995 -183.765 161.325 -183.435 ;
        RECT 160.995 -185.125 161.325 -184.795 ;
        RECT 160.995 -186.485 161.325 -186.155 ;
        RECT 160.995 -187.845 161.325 -187.515 ;
        RECT 160.995 -189.205 161.325 -188.875 ;
        RECT 160.995 -190.565 161.325 -190.235 ;
        RECT 160.995 -191.925 161.325 -191.595 ;
        RECT 160.995 -193.285 161.325 -192.955 ;
        RECT 160.995 -194.645 161.325 -194.315 ;
        RECT 160.995 -196.005 161.325 -195.675 ;
        RECT 160.995 -197.365 161.325 -197.035 ;
        RECT 160.995 -198.725 161.325 -198.395 ;
        RECT 160.995 -200.085 161.325 -199.755 ;
        RECT 160.995 -201.445 161.325 -201.115 ;
        RECT 160.995 -202.805 161.325 -202.475 ;
        RECT 160.995 -204.165 161.325 -203.835 ;
        RECT 160.995 -205.525 161.325 -205.195 ;
        RECT 160.995 -206.885 161.325 -206.555 ;
        RECT 160.995 -208.245 161.325 -207.915 ;
        RECT 160.995 -209.605 161.325 -209.275 ;
        RECT 160.995 -210.965 161.325 -210.635 ;
        RECT 160.995 -212.325 161.325 -211.995 ;
        RECT 160.995 -213.685 161.325 -213.355 ;
        RECT 160.995 -215.045 161.325 -214.715 ;
        RECT 160.995 -216.405 161.325 -216.075 ;
        RECT 160.995 -217.765 161.325 -217.435 ;
        RECT 160.995 -219.125 161.325 -218.795 ;
        RECT 160.995 -221.37 161.325 -220.24 ;
        RECT 161 -221.485 161.32 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.91 -121.535 162.24 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 162.355 129.8 162.685 130.93 ;
        RECT 162.355 127.675 162.685 128.005 ;
        RECT 162.355 126.315 162.685 126.645 ;
        RECT 162.355 124.955 162.685 125.285 ;
        RECT 162.355 123.595 162.685 123.925 ;
        RECT 162.36 123.595 162.68 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.715 129.8 164.045 130.93 ;
        RECT 163.715 127.675 164.045 128.005 ;
        RECT 163.715 126.315 164.045 126.645 ;
        RECT 163.715 124.955 164.045 125.285 ;
        RECT 163.715 123.595 164.045 123.925 ;
        RECT 163.72 123.595 164.04 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.715 -1.525 164.045 -1.195 ;
        RECT 163.715 -2.885 164.045 -2.555 ;
        RECT 163.72 -3.56 164.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.075 129.8 165.405 130.93 ;
        RECT 165.075 127.675 165.405 128.005 ;
        RECT 165.075 126.315 165.405 126.645 ;
        RECT 165.075 124.955 165.405 125.285 ;
        RECT 165.075 123.595 165.405 123.925 ;
        RECT 165.08 123.595 165.4 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.075 -1.525 165.405 -1.195 ;
        RECT 165.075 -2.885 165.405 -2.555 ;
        RECT 165.08 -3.56 165.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.075 -213.685 165.405 -213.355 ;
        RECT 165.075 -215.045 165.405 -214.715 ;
        RECT 165.075 -216.405 165.405 -216.075 ;
        RECT 165.075 -217.765 165.405 -217.435 ;
        RECT 165.075 -219.125 165.405 -218.795 ;
        RECT 165.075 -221.37 165.405 -220.24 ;
        RECT 165.08 -221.485 165.4 -118.155 ;
        RECT 165.075 -118.485 165.405 -118.155 ;
        RECT 165.075 -119.845 165.405 -119.515 ;
        RECT 165.075 -121.205 165.405 -120.875 ;
        RECT 165.075 -122.565 165.405 -122.235 ;
        RECT 165.075 -123.925 165.405 -123.595 ;
        RECT 165.075 -125.285 165.405 -124.955 ;
        RECT 165.075 -126.645 165.405 -126.315 ;
        RECT 165.075 -128.005 165.405 -127.675 ;
        RECT 165.075 -129.365 165.405 -129.035 ;
        RECT 165.075 -130.725 165.405 -130.395 ;
        RECT 165.075 -132.085 165.405 -131.755 ;
        RECT 165.075 -133.445 165.405 -133.115 ;
        RECT 165.075 -134.805 165.405 -134.475 ;
        RECT 165.075 -136.165 165.405 -135.835 ;
        RECT 165.075 -137.525 165.405 -137.195 ;
        RECT 165.075 -138.885 165.405 -138.555 ;
        RECT 165.075 -140.245 165.405 -139.915 ;
        RECT 165.075 -141.605 165.405 -141.275 ;
        RECT 165.075 -142.965 165.405 -142.635 ;
        RECT 165.075 -144.325 165.405 -143.995 ;
        RECT 165.075 -145.685 165.405 -145.355 ;
        RECT 165.075 -147.045 165.405 -146.715 ;
        RECT 165.075 -148.405 165.405 -148.075 ;
        RECT 165.075 -149.765 165.405 -149.435 ;
        RECT 165.075 -151.125 165.405 -150.795 ;
        RECT 165.075 -152.485 165.405 -152.155 ;
        RECT 165.075 -153.845 165.405 -153.515 ;
        RECT 165.075 -155.205 165.405 -154.875 ;
        RECT 165.075 -156.565 165.405 -156.235 ;
        RECT 165.075 -157.925 165.405 -157.595 ;
        RECT 165.075 -159.285 165.405 -158.955 ;
        RECT 165.075 -160.645 165.405 -160.315 ;
        RECT 165.075 -162.005 165.405 -161.675 ;
        RECT 165.075 -163.365 165.405 -163.035 ;
        RECT 165.075 -164.725 165.405 -164.395 ;
        RECT 165.075 -166.085 165.405 -165.755 ;
        RECT 165.075 -167.445 165.405 -167.115 ;
        RECT 165.075 -168.805 165.405 -168.475 ;
        RECT 165.075 -170.165 165.405 -169.835 ;
        RECT 165.075 -171.525 165.405 -171.195 ;
        RECT 165.075 -172.885 165.405 -172.555 ;
        RECT 165.075 -174.245 165.405 -173.915 ;
        RECT 165.075 -175.605 165.405 -175.275 ;
        RECT 165.075 -176.965 165.405 -176.635 ;
        RECT 165.075 -178.325 165.405 -177.995 ;
        RECT 165.075 -179.685 165.405 -179.355 ;
        RECT 165.075 -181.045 165.405 -180.715 ;
        RECT 165.075 -182.405 165.405 -182.075 ;
        RECT 165.075 -183.765 165.405 -183.435 ;
        RECT 165.075 -185.125 165.405 -184.795 ;
        RECT 165.075 -186.485 165.405 -186.155 ;
        RECT 165.075 -187.845 165.405 -187.515 ;
        RECT 165.075 -189.205 165.405 -188.875 ;
        RECT 165.075 -190.565 165.405 -190.235 ;
        RECT 165.075 -191.925 165.405 -191.595 ;
        RECT 165.075 -193.285 165.405 -192.955 ;
        RECT 165.075 -194.645 165.405 -194.315 ;
        RECT 165.075 -196.005 165.405 -195.675 ;
        RECT 165.075 -197.365 165.405 -197.035 ;
        RECT 165.075 -198.725 165.405 -198.395 ;
        RECT 165.075 -200.085 165.405 -199.755 ;
        RECT 165.075 -201.445 165.405 -201.115 ;
        RECT 165.075 -202.805 165.405 -202.475 ;
        RECT 165.075 -204.165 165.405 -203.835 ;
        RECT 165.075 -205.525 165.405 -205.195 ;
        RECT 165.075 -206.885 165.405 -206.555 ;
        RECT 165.075 -208.245 165.405 -207.915 ;
        RECT 165.075 -209.605 165.405 -209.275 ;
        RECT 165.075 -210.965 165.405 -210.635 ;
        RECT 165.075 -212.325 165.405 -211.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.595 129.8 106.925 130.93 ;
        RECT 106.595 127.675 106.925 128.005 ;
        RECT 106.595 126.315 106.925 126.645 ;
        RECT 106.595 124.955 106.925 125.285 ;
        RECT 106.595 123.595 106.925 123.925 ;
        RECT 106.6 123.595 106.92 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.595 -122.565 106.925 -122.235 ;
        RECT 106.595 -123.925 106.925 -123.595 ;
        RECT 106.595 -125.285 106.925 -124.955 ;
        RECT 106.595 -126.645 106.925 -126.315 ;
        RECT 106.595 -128.005 106.925 -127.675 ;
        RECT 106.595 -129.365 106.925 -129.035 ;
        RECT 106.595 -130.725 106.925 -130.395 ;
        RECT 106.595 -132.085 106.925 -131.755 ;
        RECT 106.595 -133.445 106.925 -133.115 ;
        RECT 106.595 -134.805 106.925 -134.475 ;
        RECT 106.595 -136.165 106.925 -135.835 ;
        RECT 106.595 -137.525 106.925 -137.195 ;
        RECT 106.595 -138.885 106.925 -138.555 ;
        RECT 106.595 -140.245 106.925 -139.915 ;
        RECT 106.595 -141.605 106.925 -141.275 ;
        RECT 106.595 -142.965 106.925 -142.635 ;
        RECT 106.595 -144.325 106.925 -143.995 ;
        RECT 106.595 -145.685 106.925 -145.355 ;
        RECT 106.595 -147.045 106.925 -146.715 ;
        RECT 106.595 -148.405 106.925 -148.075 ;
        RECT 106.595 -149.765 106.925 -149.435 ;
        RECT 106.595 -151.125 106.925 -150.795 ;
        RECT 106.595 -152.485 106.925 -152.155 ;
        RECT 106.595 -153.845 106.925 -153.515 ;
        RECT 106.595 -155.205 106.925 -154.875 ;
        RECT 106.595 -156.565 106.925 -156.235 ;
        RECT 106.595 -157.925 106.925 -157.595 ;
        RECT 106.595 -159.285 106.925 -158.955 ;
        RECT 106.595 -160.645 106.925 -160.315 ;
        RECT 106.595 -162.005 106.925 -161.675 ;
        RECT 106.595 -163.365 106.925 -163.035 ;
        RECT 106.595 -164.725 106.925 -164.395 ;
        RECT 106.595 -166.085 106.925 -165.755 ;
        RECT 106.595 -167.445 106.925 -167.115 ;
        RECT 106.595 -168.805 106.925 -168.475 ;
        RECT 106.595 -170.165 106.925 -169.835 ;
        RECT 106.595 -171.525 106.925 -171.195 ;
        RECT 106.595 -172.885 106.925 -172.555 ;
        RECT 106.595 -174.245 106.925 -173.915 ;
        RECT 106.595 -175.605 106.925 -175.275 ;
        RECT 106.595 -176.965 106.925 -176.635 ;
        RECT 106.595 -178.325 106.925 -177.995 ;
        RECT 106.595 -179.685 106.925 -179.355 ;
        RECT 106.595 -181.045 106.925 -180.715 ;
        RECT 106.595 -182.405 106.925 -182.075 ;
        RECT 106.595 -183.765 106.925 -183.435 ;
        RECT 106.595 -185.125 106.925 -184.795 ;
        RECT 106.595 -186.485 106.925 -186.155 ;
        RECT 106.595 -187.845 106.925 -187.515 ;
        RECT 106.595 -189.205 106.925 -188.875 ;
        RECT 106.595 -190.565 106.925 -190.235 ;
        RECT 106.595 -191.925 106.925 -191.595 ;
        RECT 106.595 -193.285 106.925 -192.955 ;
        RECT 106.595 -194.645 106.925 -194.315 ;
        RECT 106.595 -196.005 106.925 -195.675 ;
        RECT 106.595 -197.365 106.925 -197.035 ;
        RECT 106.595 -198.725 106.925 -198.395 ;
        RECT 106.595 -200.085 106.925 -199.755 ;
        RECT 106.595 -201.445 106.925 -201.115 ;
        RECT 106.595 -202.805 106.925 -202.475 ;
        RECT 106.595 -204.165 106.925 -203.835 ;
        RECT 106.595 -205.525 106.925 -205.195 ;
        RECT 106.595 -206.885 106.925 -206.555 ;
        RECT 106.595 -208.245 106.925 -207.915 ;
        RECT 106.595 -209.605 106.925 -209.275 ;
        RECT 106.595 -210.965 106.925 -210.635 ;
        RECT 106.595 -212.325 106.925 -211.995 ;
        RECT 106.595 -213.685 106.925 -213.355 ;
        RECT 106.595 -215.045 106.925 -214.715 ;
        RECT 106.595 -216.405 106.925 -216.075 ;
        RECT 106.595 -217.765 106.925 -217.435 ;
        RECT 106.595 -219.125 106.925 -218.795 ;
        RECT 106.595 -221.37 106.925 -220.24 ;
        RECT 106.6 -221.485 106.92 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.01 -121.535 107.34 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.955 129.8 108.285 130.93 ;
        RECT 107.955 127.675 108.285 128.005 ;
        RECT 107.955 126.315 108.285 126.645 ;
        RECT 107.955 124.955 108.285 125.285 ;
        RECT 107.955 123.595 108.285 123.925 ;
        RECT 107.96 123.595 108.28 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.955 -1.525 108.285 -1.195 ;
        RECT 107.955 -2.885 108.285 -2.555 ;
        RECT 107.96 -3.56 108.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.315 129.8 109.645 130.93 ;
        RECT 109.315 127.675 109.645 128.005 ;
        RECT 109.315 126.315 109.645 126.645 ;
        RECT 109.315 124.955 109.645 125.285 ;
        RECT 109.315 123.595 109.645 123.925 ;
        RECT 109.32 123.595 109.64 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.315 -1.525 109.645 -1.195 ;
        RECT 109.315 -2.885 109.645 -2.555 ;
        RECT 109.32 -3.56 109.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.675 129.8 111.005 130.93 ;
        RECT 110.675 127.675 111.005 128.005 ;
        RECT 110.675 126.315 111.005 126.645 ;
        RECT 110.675 124.955 111.005 125.285 ;
        RECT 110.675 123.595 111.005 123.925 ;
        RECT 110.68 123.595 111 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.675 -1.525 111.005 -1.195 ;
        RECT 110.675 -2.885 111.005 -2.555 ;
        RECT 110.68 -3.56 111 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.675 -118.485 111.005 -118.155 ;
        RECT 110.675 -119.845 111.005 -119.515 ;
        RECT 110.675 -121.205 111.005 -120.875 ;
        RECT 110.675 -122.565 111.005 -122.235 ;
        RECT 110.675 -123.925 111.005 -123.595 ;
        RECT 110.675 -125.285 111.005 -124.955 ;
        RECT 110.675 -126.645 111.005 -126.315 ;
        RECT 110.675 -128.005 111.005 -127.675 ;
        RECT 110.675 -129.365 111.005 -129.035 ;
        RECT 110.675 -130.725 111.005 -130.395 ;
        RECT 110.675 -132.085 111.005 -131.755 ;
        RECT 110.675 -133.445 111.005 -133.115 ;
        RECT 110.675 -134.805 111.005 -134.475 ;
        RECT 110.675 -136.165 111.005 -135.835 ;
        RECT 110.675 -137.525 111.005 -137.195 ;
        RECT 110.675 -138.885 111.005 -138.555 ;
        RECT 110.675 -140.245 111.005 -139.915 ;
        RECT 110.675 -141.605 111.005 -141.275 ;
        RECT 110.675 -142.965 111.005 -142.635 ;
        RECT 110.675 -144.325 111.005 -143.995 ;
        RECT 110.675 -145.685 111.005 -145.355 ;
        RECT 110.675 -147.045 111.005 -146.715 ;
        RECT 110.675 -148.405 111.005 -148.075 ;
        RECT 110.675 -149.765 111.005 -149.435 ;
        RECT 110.675 -151.125 111.005 -150.795 ;
        RECT 110.675 -152.485 111.005 -152.155 ;
        RECT 110.675 -153.845 111.005 -153.515 ;
        RECT 110.675 -155.205 111.005 -154.875 ;
        RECT 110.675 -156.565 111.005 -156.235 ;
        RECT 110.675 -157.925 111.005 -157.595 ;
        RECT 110.675 -159.285 111.005 -158.955 ;
        RECT 110.675 -160.645 111.005 -160.315 ;
        RECT 110.675 -162.005 111.005 -161.675 ;
        RECT 110.675 -163.365 111.005 -163.035 ;
        RECT 110.675 -164.725 111.005 -164.395 ;
        RECT 110.675 -166.085 111.005 -165.755 ;
        RECT 110.675 -167.445 111.005 -167.115 ;
        RECT 110.675 -168.805 111.005 -168.475 ;
        RECT 110.675 -170.165 111.005 -169.835 ;
        RECT 110.675 -171.525 111.005 -171.195 ;
        RECT 110.675 -172.885 111.005 -172.555 ;
        RECT 110.675 -174.245 111.005 -173.915 ;
        RECT 110.675 -175.605 111.005 -175.275 ;
        RECT 110.675 -176.965 111.005 -176.635 ;
        RECT 110.675 -178.325 111.005 -177.995 ;
        RECT 110.675 -179.685 111.005 -179.355 ;
        RECT 110.675 -181.045 111.005 -180.715 ;
        RECT 110.675 -182.405 111.005 -182.075 ;
        RECT 110.675 -183.765 111.005 -183.435 ;
        RECT 110.675 -185.125 111.005 -184.795 ;
        RECT 110.675 -186.485 111.005 -186.155 ;
        RECT 110.675 -187.845 111.005 -187.515 ;
        RECT 110.675 -189.205 111.005 -188.875 ;
        RECT 110.675 -190.565 111.005 -190.235 ;
        RECT 110.675 -191.925 111.005 -191.595 ;
        RECT 110.675 -193.285 111.005 -192.955 ;
        RECT 110.675 -194.645 111.005 -194.315 ;
        RECT 110.675 -196.005 111.005 -195.675 ;
        RECT 110.675 -197.365 111.005 -197.035 ;
        RECT 110.675 -198.725 111.005 -198.395 ;
        RECT 110.675 -200.085 111.005 -199.755 ;
        RECT 110.675 -201.445 111.005 -201.115 ;
        RECT 110.675 -202.805 111.005 -202.475 ;
        RECT 110.675 -204.165 111.005 -203.835 ;
        RECT 110.675 -205.525 111.005 -205.195 ;
        RECT 110.675 -206.885 111.005 -206.555 ;
        RECT 110.675 -208.245 111.005 -207.915 ;
        RECT 110.675 -209.605 111.005 -209.275 ;
        RECT 110.675 -210.965 111.005 -210.635 ;
        RECT 110.675 -212.325 111.005 -211.995 ;
        RECT 110.675 -213.685 111.005 -213.355 ;
        RECT 110.675 -215.045 111.005 -214.715 ;
        RECT 110.675 -216.405 111.005 -216.075 ;
        RECT 110.675 -217.765 111.005 -217.435 ;
        RECT 110.675 -219.125 111.005 -218.795 ;
        RECT 110.675 -221.37 111.005 -220.24 ;
        RECT 110.68 -221.485 111 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.035 129.8 112.365 130.93 ;
        RECT 112.035 127.675 112.365 128.005 ;
        RECT 112.035 126.315 112.365 126.645 ;
        RECT 112.035 124.955 112.365 125.285 ;
        RECT 112.035 123.595 112.365 123.925 ;
        RECT 112.04 123.595 112.36 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.035 -122.565 112.365 -122.235 ;
        RECT 112.035 -123.925 112.365 -123.595 ;
        RECT 112.035 -125.285 112.365 -124.955 ;
        RECT 112.035 -126.645 112.365 -126.315 ;
        RECT 112.035 -128.005 112.365 -127.675 ;
        RECT 112.035 -129.365 112.365 -129.035 ;
        RECT 112.035 -130.725 112.365 -130.395 ;
        RECT 112.035 -132.085 112.365 -131.755 ;
        RECT 112.035 -133.445 112.365 -133.115 ;
        RECT 112.035 -134.805 112.365 -134.475 ;
        RECT 112.035 -136.165 112.365 -135.835 ;
        RECT 112.035 -137.525 112.365 -137.195 ;
        RECT 112.035 -138.885 112.365 -138.555 ;
        RECT 112.035 -140.245 112.365 -139.915 ;
        RECT 112.035 -141.605 112.365 -141.275 ;
        RECT 112.035 -142.965 112.365 -142.635 ;
        RECT 112.035 -144.325 112.365 -143.995 ;
        RECT 112.035 -145.685 112.365 -145.355 ;
        RECT 112.035 -147.045 112.365 -146.715 ;
        RECT 112.035 -148.405 112.365 -148.075 ;
        RECT 112.035 -149.765 112.365 -149.435 ;
        RECT 112.035 -151.125 112.365 -150.795 ;
        RECT 112.035 -152.485 112.365 -152.155 ;
        RECT 112.035 -153.845 112.365 -153.515 ;
        RECT 112.035 -155.205 112.365 -154.875 ;
        RECT 112.035 -156.565 112.365 -156.235 ;
        RECT 112.035 -157.925 112.365 -157.595 ;
        RECT 112.035 -159.285 112.365 -158.955 ;
        RECT 112.035 -160.645 112.365 -160.315 ;
        RECT 112.035 -162.005 112.365 -161.675 ;
        RECT 112.035 -163.365 112.365 -163.035 ;
        RECT 112.035 -164.725 112.365 -164.395 ;
        RECT 112.035 -166.085 112.365 -165.755 ;
        RECT 112.035 -167.445 112.365 -167.115 ;
        RECT 112.035 -168.805 112.365 -168.475 ;
        RECT 112.035 -170.165 112.365 -169.835 ;
        RECT 112.035 -171.525 112.365 -171.195 ;
        RECT 112.035 -172.885 112.365 -172.555 ;
        RECT 112.035 -174.245 112.365 -173.915 ;
        RECT 112.035 -175.605 112.365 -175.275 ;
        RECT 112.035 -176.965 112.365 -176.635 ;
        RECT 112.035 -178.325 112.365 -177.995 ;
        RECT 112.035 -179.685 112.365 -179.355 ;
        RECT 112.035 -181.045 112.365 -180.715 ;
        RECT 112.035 -182.405 112.365 -182.075 ;
        RECT 112.035 -183.765 112.365 -183.435 ;
        RECT 112.035 -185.125 112.365 -184.795 ;
        RECT 112.035 -186.485 112.365 -186.155 ;
        RECT 112.035 -187.845 112.365 -187.515 ;
        RECT 112.035 -189.205 112.365 -188.875 ;
        RECT 112.035 -190.565 112.365 -190.235 ;
        RECT 112.035 -191.925 112.365 -191.595 ;
        RECT 112.035 -193.285 112.365 -192.955 ;
        RECT 112.035 -194.645 112.365 -194.315 ;
        RECT 112.035 -196.005 112.365 -195.675 ;
        RECT 112.035 -197.365 112.365 -197.035 ;
        RECT 112.035 -198.725 112.365 -198.395 ;
        RECT 112.035 -200.085 112.365 -199.755 ;
        RECT 112.035 -201.445 112.365 -201.115 ;
        RECT 112.035 -202.805 112.365 -202.475 ;
        RECT 112.035 -204.165 112.365 -203.835 ;
        RECT 112.035 -205.525 112.365 -205.195 ;
        RECT 112.035 -206.885 112.365 -206.555 ;
        RECT 112.035 -208.245 112.365 -207.915 ;
        RECT 112.035 -209.605 112.365 -209.275 ;
        RECT 112.035 -210.965 112.365 -210.635 ;
        RECT 112.035 -212.325 112.365 -211.995 ;
        RECT 112.035 -213.685 112.365 -213.355 ;
        RECT 112.035 -215.045 112.365 -214.715 ;
        RECT 112.035 -216.405 112.365 -216.075 ;
        RECT 112.035 -217.765 112.365 -217.435 ;
        RECT 112.035 -219.125 112.365 -218.795 ;
        RECT 112.035 -221.37 112.365 -220.24 ;
        RECT 112.04 -221.485 112.36 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.11 -121.535 113.44 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.395 129.8 113.725 130.93 ;
        RECT 113.395 127.675 113.725 128.005 ;
        RECT 113.395 126.315 113.725 126.645 ;
        RECT 113.395 124.955 113.725 125.285 ;
        RECT 113.395 123.595 113.725 123.925 ;
        RECT 113.4 123.595 113.72 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.755 129.8 115.085 130.93 ;
        RECT 114.755 127.675 115.085 128.005 ;
        RECT 114.755 126.315 115.085 126.645 ;
        RECT 114.755 124.955 115.085 125.285 ;
        RECT 114.755 123.595 115.085 123.925 ;
        RECT 114.76 123.595 115.08 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.755 -1.525 115.085 -1.195 ;
        RECT 114.755 -2.885 115.085 -2.555 ;
        RECT 114.76 -3.56 115.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.115 129.8 116.445 130.93 ;
        RECT 116.115 127.675 116.445 128.005 ;
        RECT 116.115 126.315 116.445 126.645 ;
        RECT 116.115 124.955 116.445 125.285 ;
        RECT 116.115 123.595 116.445 123.925 ;
        RECT 116.12 123.595 116.44 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.115 -1.525 116.445 -1.195 ;
        RECT 116.115 -2.885 116.445 -2.555 ;
        RECT 116.12 -3.56 116.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.475 129.8 117.805 130.93 ;
        RECT 117.475 127.675 117.805 128.005 ;
        RECT 117.475 126.315 117.805 126.645 ;
        RECT 117.475 124.955 117.805 125.285 ;
        RECT 117.475 123.595 117.805 123.925 ;
        RECT 117.48 123.595 117.8 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.475 -1.525 117.805 -1.195 ;
        RECT 117.475 -2.885 117.805 -2.555 ;
        RECT 117.48 -3.56 117.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.475 -118.485 117.805 -118.155 ;
        RECT 117.475 -119.845 117.805 -119.515 ;
        RECT 117.475 -121.205 117.805 -120.875 ;
        RECT 117.475 -122.565 117.805 -122.235 ;
        RECT 117.475 -123.925 117.805 -123.595 ;
        RECT 117.475 -125.285 117.805 -124.955 ;
        RECT 117.475 -126.645 117.805 -126.315 ;
        RECT 117.475 -128.005 117.805 -127.675 ;
        RECT 117.475 -129.365 117.805 -129.035 ;
        RECT 117.475 -130.725 117.805 -130.395 ;
        RECT 117.475 -132.085 117.805 -131.755 ;
        RECT 117.475 -133.445 117.805 -133.115 ;
        RECT 117.475 -134.805 117.805 -134.475 ;
        RECT 117.475 -136.165 117.805 -135.835 ;
        RECT 117.475 -137.525 117.805 -137.195 ;
        RECT 117.475 -138.885 117.805 -138.555 ;
        RECT 117.475 -140.245 117.805 -139.915 ;
        RECT 117.475 -141.605 117.805 -141.275 ;
        RECT 117.475 -142.965 117.805 -142.635 ;
        RECT 117.475 -144.325 117.805 -143.995 ;
        RECT 117.475 -145.685 117.805 -145.355 ;
        RECT 117.475 -147.045 117.805 -146.715 ;
        RECT 117.475 -148.405 117.805 -148.075 ;
        RECT 117.475 -149.765 117.805 -149.435 ;
        RECT 117.475 -151.125 117.805 -150.795 ;
        RECT 117.475 -152.485 117.805 -152.155 ;
        RECT 117.475 -153.845 117.805 -153.515 ;
        RECT 117.475 -155.205 117.805 -154.875 ;
        RECT 117.475 -156.565 117.805 -156.235 ;
        RECT 117.475 -157.925 117.805 -157.595 ;
        RECT 117.475 -159.285 117.805 -158.955 ;
        RECT 117.475 -160.645 117.805 -160.315 ;
        RECT 117.475 -162.005 117.805 -161.675 ;
        RECT 117.475 -163.365 117.805 -163.035 ;
        RECT 117.475 -164.725 117.805 -164.395 ;
        RECT 117.475 -166.085 117.805 -165.755 ;
        RECT 117.475 -167.445 117.805 -167.115 ;
        RECT 117.475 -168.805 117.805 -168.475 ;
        RECT 117.475 -170.165 117.805 -169.835 ;
        RECT 117.475 -171.525 117.805 -171.195 ;
        RECT 117.475 -172.885 117.805 -172.555 ;
        RECT 117.475 -174.245 117.805 -173.915 ;
        RECT 117.475 -175.605 117.805 -175.275 ;
        RECT 117.475 -176.965 117.805 -176.635 ;
        RECT 117.475 -178.325 117.805 -177.995 ;
        RECT 117.475 -179.685 117.805 -179.355 ;
        RECT 117.475 -181.045 117.805 -180.715 ;
        RECT 117.475 -182.405 117.805 -182.075 ;
        RECT 117.475 -183.765 117.805 -183.435 ;
        RECT 117.475 -185.125 117.805 -184.795 ;
        RECT 117.475 -186.485 117.805 -186.155 ;
        RECT 117.475 -187.845 117.805 -187.515 ;
        RECT 117.475 -189.205 117.805 -188.875 ;
        RECT 117.475 -190.565 117.805 -190.235 ;
        RECT 117.475 -191.925 117.805 -191.595 ;
        RECT 117.475 -193.285 117.805 -192.955 ;
        RECT 117.475 -194.645 117.805 -194.315 ;
        RECT 117.475 -196.005 117.805 -195.675 ;
        RECT 117.475 -197.365 117.805 -197.035 ;
        RECT 117.475 -198.725 117.805 -198.395 ;
        RECT 117.475 -200.085 117.805 -199.755 ;
        RECT 117.475 -201.445 117.805 -201.115 ;
        RECT 117.475 -202.805 117.805 -202.475 ;
        RECT 117.475 -204.165 117.805 -203.835 ;
        RECT 117.475 -205.525 117.805 -205.195 ;
        RECT 117.475 -206.885 117.805 -206.555 ;
        RECT 117.475 -208.245 117.805 -207.915 ;
        RECT 117.475 -209.605 117.805 -209.275 ;
        RECT 117.475 -210.965 117.805 -210.635 ;
        RECT 117.475 -212.325 117.805 -211.995 ;
        RECT 117.475 -213.685 117.805 -213.355 ;
        RECT 117.475 -215.045 117.805 -214.715 ;
        RECT 117.475 -216.405 117.805 -216.075 ;
        RECT 117.475 -217.765 117.805 -217.435 ;
        RECT 117.475 -219.125 117.805 -218.795 ;
        RECT 117.475 -221.37 117.805 -220.24 ;
        RECT 117.48 -221.485 117.8 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.835 129.8 119.165 130.93 ;
        RECT 118.835 127.675 119.165 128.005 ;
        RECT 118.835 126.315 119.165 126.645 ;
        RECT 118.835 124.955 119.165 125.285 ;
        RECT 118.835 123.595 119.165 123.925 ;
        RECT 118.84 123.595 119.16 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.835 -122.565 119.165 -122.235 ;
        RECT 118.835 -123.925 119.165 -123.595 ;
        RECT 118.835 -125.285 119.165 -124.955 ;
        RECT 118.835 -126.645 119.165 -126.315 ;
        RECT 118.835 -128.005 119.165 -127.675 ;
        RECT 118.835 -129.365 119.165 -129.035 ;
        RECT 118.835 -130.725 119.165 -130.395 ;
        RECT 118.835 -132.085 119.165 -131.755 ;
        RECT 118.835 -133.445 119.165 -133.115 ;
        RECT 118.835 -134.805 119.165 -134.475 ;
        RECT 118.835 -136.165 119.165 -135.835 ;
        RECT 118.835 -137.525 119.165 -137.195 ;
        RECT 118.835 -138.885 119.165 -138.555 ;
        RECT 118.835 -140.245 119.165 -139.915 ;
        RECT 118.835 -141.605 119.165 -141.275 ;
        RECT 118.835 -142.965 119.165 -142.635 ;
        RECT 118.835 -144.325 119.165 -143.995 ;
        RECT 118.835 -145.685 119.165 -145.355 ;
        RECT 118.835 -147.045 119.165 -146.715 ;
        RECT 118.835 -148.405 119.165 -148.075 ;
        RECT 118.835 -149.765 119.165 -149.435 ;
        RECT 118.835 -151.125 119.165 -150.795 ;
        RECT 118.835 -152.485 119.165 -152.155 ;
        RECT 118.835 -153.845 119.165 -153.515 ;
        RECT 118.835 -155.205 119.165 -154.875 ;
        RECT 118.835 -156.565 119.165 -156.235 ;
        RECT 118.835 -157.925 119.165 -157.595 ;
        RECT 118.835 -159.285 119.165 -158.955 ;
        RECT 118.835 -160.645 119.165 -160.315 ;
        RECT 118.835 -162.005 119.165 -161.675 ;
        RECT 118.835 -163.365 119.165 -163.035 ;
        RECT 118.835 -164.725 119.165 -164.395 ;
        RECT 118.835 -166.085 119.165 -165.755 ;
        RECT 118.835 -167.445 119.165 -167.115 ;
        RECT 118.835 -168.805 119.165 -168.475 ;
        RECT 118.835 -170.165 119.165 -169.835 ;
        RECT 118.835 -171.525 119.165 -171.195 ;
        RECT 118.835 -172.885 119.165 -172.555 ;
        RECT 118.835 -174.245 119.165 -173.915 ;
        RECT 118.835 -175.605 119.165 -175.275 ;
        RECT 118.835 -176.965 119.165 -176.635 ;
        RECT 118.835 -178.325 119.165 -177.995 ;
        RECT 118.835 -179.685 119.165 -179.355 ;
        RECT 118.835 -181.045 119.165 -180.715 ;
        RECT 118.835 -182.405 119.165 -182.075 ;
        RECT 118.835 -183.765 119.165 -183.435 ;
        RECT 118.835 -185.125 119.165 -184.795 ;
        RECT 118.835 -186.485 119.165 -186.155 ;
        RECT 118.835 -187.845 119.165 -187.515 ;
        RECT 118.835 -189.205 119.165 -188.875 ;
        RECT 118.835 -190.565 119.165 -190.235 ;
        RECT 118.835 -191.925 119.165 -191.595 ;
        RECT 118.835 -193.285 119.165 -192.955 ;
        RECT 118.835 -194.645 119.165 -194.315 ;
        RECT 118.835 -196.005 119.165 -195.675 ;
        RECT 118.835 -197.365 119.165 -197.035 ;
        RECT 118.835 -198.725 119.165 -198.395 ;
        RECT 118.835 -200.085 119.165 -199.755 ;
        RECT 118.835 -201.445 119.165 -201.115 ;
        RECT 118.835 -202.805 119.165 -202.475 ;
        RECT 118.835 -204.165 119.165 -203.835 ;
        RECT 118.835 -205.525 119.165 -205.195 ;
        RECT 118.835 -206.885 119.165 -206.555 ;
        RECT 118.835 -208.245 119.165 -207.915 ;
        RECT 118.835 -209.605 119.165 -209.275 ;
        RECT 118.835 -210.965 119.165 -210.635 ;
        RECT 118.835 -212.325 119.165 -211.995 ;
        RECT 118.835 -213.685 119.165 -213.355 ;
        RECT 118.835 -215.045 119.165 -214.715 ;
        RECT 118.835 -216.405 119.165 -216.075 ;
        RECT 118.835 -217.765 119.165 -217.435 ;
        RECT 118.835 -219.125 119.165 -218.795 ;
        RECT 118.835 -221.37 119.165 -220.24 ;
        RECT 118.84 -221.485 119.16 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.21 -121.535 119.54 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.195 129.8 120.525 130.93 ;
        RECT 120.195 127.675 120.525 128.005 ;
        RECT 120.195 126.315 120.525 126.645 ;
        RECT 120.195 124.955 120.525 125.285 ;
        RECT 120.195 123.595 120.525 123.925 ;
        RECT 120.2 123.595 120.52 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.195 -1.525 120.525 -1.195 ;
        RECT 120.195 -2.885 120.525 -2.555 ;
        RECT 120.2 -3.56 120.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.555 129.8 121.885 130.93 ;
        RECT 121.555 127.675 121.885 128.005 ;
        RECT 121.555 126.315 121.885 126.645 ;
        RECT 121.555 124.955 121.885 125.285 ;
        RECT 121.555 123.595 121.885 123.925 ;
        RECT 121.56 123.595 121.88 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.555 -1.525 121.885 -1.195 ;
        RECT 121.555 -2.885 121.885 -2.555 ;
        RECT 121.56 -3.56 121.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.915 129.8 123.245 130.93 ;
        RECT 122.915 127.675 123.245 128.005 ;
        RECT 122.915 126.315 123.245 126.645 ;
        RECT 122.915 124.955 123.245 125.285 ;
        RECT 122.915 123.595 123.245 123.925 ;
        RECT 122.92 123.595 123.24 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.915 -1.525 123.245 -1.195 ;
        RECT 122.915 -2.885 123.245 -2.555 ;
        RECT 122.92 -3.56 123.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.915 -118.485 123.245 -118.155 ;
        RECT 122.915 -119.845 123.245 -119.515 ;
        RECT 122.915 -121.205 123.245 -120.875 ;
        RECT 122.915 -122.565 123.245 -122.235 ;
        RECT 122.915 -123.925 123.245 -123.595 ;
        RECT 122.915 -125.285 123.245 -124.955 ;
        RECT 122.915 -126.645 123.245 -126.315 ;
        RECT 122.915 -128.005 123.245 -127.675 ;
        RECT 122.915 -129.365 123.245 -129.035 ;
        RECT 122.915 -130.725 123.245 -130.395 ;
        RECT 122.915 -132.085 123.245 -131.755 ;
        RECT 122.915 -133.445 123.245 -133.115 ;
        RECT 122.915 -134.805 123.245 -134.475 ;
        RECT 122.915 -136.165 123.245 -135.835 ;
        RECT 122.915 -137.525 123.245 -137.195 ;
        RECT 122.915 -138.885 123.245 -138.555 ;
        RECT 122.915 -140.245 123.245 -139.915 ;
        RECT 122.915 -141.605 123.245 -141.275 ;
        RECT 122.915 -142.965 123.245 -142.635 ;
        RECT 122.915 -144.325 123.245 -143.995 ;
        RECT 122.915 -145.685 123.245 -145.355 ;
        RECT 122.915 -147.045 123.245 -146.715 ;
        RECT 122.915 -148.405 123.245 -148.075 ;
        RECT 122.915 -149.765 123.245 -149.435 ;
        RECT 122.915 -151.125 123.245 -150.795 ;
        RECT 122.915 -152.485 123.245 -152.155 ;
        RECT 122.915 -153.845 123.245 -153.515 ;
        RECT 122.915 -155.205 123.245 -154.875 ;
        RECT 122.915 -156.565 123.245 -156.235 ;
        RECT 122.915 -157.925 123.245 -157.595 ;
        RECT 122.915 -159.285 123.245 -158.955 ;
        RECT 122.915 -160.645 123.245 -160.315 ;
        RECT 122.915 -162.005 123.245 -161.675 ;
        RECT 122.915 -163.365 123.245 -163.035 ;
        RECT 122.915 -164.725 123.245 -164.395 ;
        RECT 122.915 -166.085 123.245 -165.755 ;
        RECT 122.915 -167.445 123.245 -167.115 ;
        RECT 122.915 -168.805 123.245 -168.475 ;
        RECT 122.915 -170.165 123.245 -169.835 ;
        RECT 122.915 -171.525 123.245 -171.195 ;
        RECT 122.915 -172.885 123.245 -172.555 ;
        RECT 122.915 -174.245 123.245 -173.915 ;
        RECT 122.915 -175.605 123.245 -175.275 ;
        RECT 122.915 -176.965 123.245 -176.635 ;
        RECT 122.915 -178.325 123.245 -177.995 ;
        RECT 122.915 -179.685 123.245 -179.355 ;
        RECT 122.915 -181.045 123.245 -180.715 ;
        RECT 122.915 -182.405 123.245 -182.075 ;
        RECT 122.915 -183.765 123.245 -183.435 ;
        RECT 122.915 -185.125 123.245 -184.795 ;
        RECT 122.915 -186.485 123.245 -186.155 ;
        RECT 122.915 -187.845 123.245 -187.515 ;
        RECT 122.915 -189.205 123.245 -188.875 ;
        RECT 122.915 -190.565 123.245 -190.235 ;
        RECT 122.915 -191.925 123.245 -191.595 ;
        RECT 122.915 -193.285 123.245 -192.955 ;
        RECT 122.915 -194.645 123.245 -194.315 ;
        RECT 122.915 -196.005 123.245 -195.675 ;
        RECT 122.915 -197.365 123.245 -197.035 ;
        RECT 122.915 -198.725 123.245 -198.395 ;
        RECT 122.915 -200.085 123.245 -199.755 ;
        RECT 122.915 -201.445 123.245 -201.115 ;
        RECT 122.915 -202.805 123.245 -202.475 ;
        RECT 122.915 -204.165 123.245 -203.835 ;
        RECT 122.915 -205.525 123.245 -205.195 ;
        RECT 122.915 -206.885 123.245 -206.555 ;
        RECT 122.915 -208.245 123.245 -207.915 ;
        RECT 122.915 -209.605 123.245 -209.275 ;
        RECT 122.915 -210.965 123.245 -210.635 ;
        RECT 122.915 -212.325 123.245 -211.995 ;
        RECT 122.915 -213.685 123.245 -213.355 ;
        RECT 122.915 -215.045 123.245 -214.715 ;
        RECT 122.915 -216.405 123.245 -216.075 ;
        RECT 122.915 -217.765 123.245 -217.435 ;
        RECT 122.915 -219.125 123.245 -218.795 ;
        RECT 122.915 -221.37 123.245 -220.24 ;
        RECT 122.92 -221.485 123.24 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.275 129.8 124.605 130.93 ;
        RECT 124.275 127.675 124.605 128.005 ;
        RECT 124.275 126.315 124.605 126.645 ;
        RECT 124.275 124.955 124.605 125.285 ;
        RECT 124.275 123.595 124.605 123.925 ;
        RECT 124.28 123.595 124.6 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.275 -122.565 124.605 -122.235 ;
        RECT 124.275 -123.925 124.605 -123.595 ;
        RECT 124.275 -125.285 124.605 -124.955 ;
        RECT 124.275 -126.645 124.605 -126.315 ;
        RECT 124.275 -128.005 124.605 -127.675 ;
        RECT 124.275 -129.365 124.605 -129.035 ;
        RECT 124.275 -130.725 124.605 -130.395 ;
        RECT 124.275 -132.085 124.605 -131.755 ;
        RECT 124.275 -133.445 124.605 -133.115 ;
        RECT 124.275 -134.805 124.605 -134.475 ;
        RECT 124.275 -136.165 124.605 -135.835 ;
        RECT 124.275 -137.525 124.605 -137.195 ;
        RECT 124.275 -138.885 124.605 -138.555 ;
        RECT 124.275 -140.245 124.605 -139.915 ;
        RECT 124.275 -141.605 124.605 -141.275 ;
        RECT 124.275 -142.965 124.605 -142.635 ;
        RECT 124.275 -144.325 124.605 -143.995 ;
        RECT 124.275 -145.685 124.605 -145.355 ;
        RECT 124.275 -147.045 124.605 -146.715 ;
        RECT 124.275 -148.405 124.605 -148.075 ;
        RECT 124.275 -149.765 124.605 -149.435 ;
        RECT 124.275 -151.125 124.605 -150.795 ;
        RECT 124.275 -152.485 124.605 -152.155 ;
        RECT 124.275 -153.845 124.605 -153.515 ;
        RECT 124.275 -155.205 124.605 -154.875 ;
        RECT 124.275 -156.565 124.605 -156.235 ;
        RECT 124.275 -157.925 124.605 -157.595 ;
        RECT 124.275 -159.285 124.605 -158.955 ;
        RECT 124.275 -160.645 124.605 -160.315 ;
        RECT 124.275 -162.005 124.605 -161.675 ;
        RECT 124.275 -163.365 124.605 -163.035 ;
        RECT 124.275 -164.725 124.605 -164.395 ;
        RECT 124.275 -166.085 124.605 -165.755 ;
        RECT 124.275 -167.445 124.605 -167.115 ;
        RECT 124.275 -168.805 124.605 -168.475 ;
        RECT 124.275 -170.165 124.605 -169.835 ;
        RECT 124.275 -171.525 124.605 -171.195 ;
        RECT 124.275 -172.885 124.605 -172.555 ;
        RECT 124.275 -174.245 124.605 -173.915 ;
        RECT 124.275 -175.605 124.605 -175.275 ;
        RECT 124.275 -176.965 124.605 -176.635 ;
        RECT 124.275 -178.325 124.605 -177.995 ;
        RECT 124.275 -179.685 124.605 -179.355 ;
        RECT 124.275 -181.045 124.605 -180.715 ;
        RECT 124.275 -182.405 124.605 -182.075 ;
        RECT 124.275 -183.765 124.605 -183.435 ;
        RECT 124.275 -185.125 124.605 -184.795 ;
        RECT 124.275 -186.485 124.605 -186.155 ;
        RECT 124.275 -187.845 124.605 -187.515 ;
        RECT 124.275 -189.205 124.605 -188.875 ;
        RECT 124.275 -190.565 124.605 -190.235 ;
        RECT 124.275 -191.925 124.605 -191.595 ;
        RECT 124.275 -193.285 124.605 -192.955 ;
        RECT 124.275 -194.645 124.605 -194.315 ;
        RECT 124.275 -196.005 124.605 -195.675 ;
        RECT 124.275 -197.365 124.605 -197.035 ;
        RECT 124.275 -198.725 124.605 -198.395 ;
        RECT 124.275 -200.085 124.605 -199.755 ;
        RECT 124.275 -201.445 124.605 -201.115 ;
        RECT 124.275 -202.805 124.605 -202.475 ;
        RECT 124.275 -204.165 124.605 -203.835 ;
        RECT 124.275 -205.525 124.605 -205.195 ;
        RECT 124.275 -206.885 124.605 -206.555 ;
        RECT 124.275 -208.245 124.605 -207.915 ;
        RECT 124.275 -209.605 124.605 -209.275 ;
        RECT 124.275 -210.965 124.605 -210.635 ;
        RECT 124.275 -212.325 124.605 -211.995 ;
        RECT 124.275 -213.685 124.605 -213.355 ;
        RECT 124.275 -215.045 124.605 -214.715 ;
        RECT 124.275 -216.405 124.605 -216.075 ;
        RECT 124.275 -217.765 124.605 -217.435 ;
        RECT 124.275 -219.125 124.605 -218.795 ;
        RECT 124.275 -221.37 124.605 -220.24 ;
        RECT 124.28 -221.485 124.6 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.31 -121.535 125.64 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.635 129.8 125.965 130.93 ;
        RECT 125.635 127.675 125.965 128.005 ;
        RECT 125.635 126.315 125.965 126.645 ;
        RECT 125.635 124.955 125.965 125.285 ;
        RECT 125.635 123.595 125.965 123.925 ;
        RECT 125.64 123.595 125.96 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.995 129.8 127.325 130.93 ;
        RECT 126.995 127.675 127.325 128.005 ;
        RECT 126.995 126.315 127.325 126.645 ;
        RECT 126.995 124.955 127.325 125.285 ;
        RECT 126.995 123.595 127.325 123.925 ;
        RECT 127 123.595 127.32 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.995 -1.525 127.325 -1.195 ;
        RECT 126.995 -2.885 127.325 -2.555 ;
        RECT 127 -3.56 127.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.355 129.8 128.685 130.93 ;
        RECT 128.355 127.675 128.685 128.005 ;
        RECT 128.355 126.315 128.685 126.645 ;
        RECT 128.355 124.955 128.685 125.285 ;
        RECT 128.355 123.595 128.685 123.925 ;
        RECT 128.36 123.595 128.68 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.355 -1.525 128.685 -1.195 ;
        RECT 128.355 -2.885 128.685 -2.555 ;
        RECT 128.36 -3.56 128.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.355 -118.485 128.685 -118.155 ;
        RECT 128.355 -119.845 128.685 -119.515 ;
        RECT 128.355 -121.205 128.685 -120.875 ;
        RECT 128.355 -122.565 128.685 -122.235 ;
        RECT 128.355 -123.925 128.685 -123.595 ;
        RECT 128.355 -125.285 128.685 -124.955 ;
        RECT 128.355 -126.645 128.685 -126.315 ;
        RECT 128.355 -128.005 128.685 -127.675 ;
        RECT 128.355 -129.365 128.685 -129.035 ;
        RECT 128.355 -130.725 128.685 -130.395 ;
        RECT 128.355 -132.085 128.685 -131.755 ;
        RECT 128.355 -133.445 128.685 -133.115 ;
        RECT 128.355 -134.805 128.685 -134.475 ;
        RECT 128.355 -136.165 128.685 -135.835 ;
        RECT 128.355 -137.525 128.685 -137.195 ;
        RECT 128.355 -138.885 128.685 -138.555 ;
        RECT 128.355 -140.245 128.685 -139.915 ;
        RECT 128.355 -141.605 128.685 -141.275 ;
        RECT 128.355 -142.965 128.685 -142.635 ;
        RECT 128.355 -144.325 128.685 -143.995 ;
        RECT 128.355 -145.685 128.685 -145.355 ;
        RECT 128.355 -147.045 128.685 -146.715 ;
        RECT 128.355 -148.405 128.685 -148.075 ;
        RECT 128.355 -149.765 128.685 -149.435 ;
        RECT 128.355 -151.125 128.685 -150.795 ;
        RECT 128.355 -152.485 128.685 -152.155 ;
        RECT 128.355 -153.845 128.685 -153.515 ;
        RECT 128.355 -155.205 128.685 -154.875 ;
        RECT 128.355 -156.565 128.685 -156.235 ;
        RECT 128.355 -157.925 128.685 -157.595 ;
        RECT 128.355 -159.285 128.685 -158.955 ;
        RECT 128.355 -160.645 128.685 -160.315 ;
        RECT 128.355 -162.005 128.685 -161.675 ;
        RECT 128.355 -163.365 128.685 -163.035 ;
        RECT 128.355 -164.725 128.685 -164.395 ;
        RECT 128.355 -166.085 128.685 -165.755 ;
        RECT 128.355 -167.445 128.685 -167.115 ;
        RECT 128.355 -168.805 128.685 -168.475 ;
        RECT 128.355 -170.165 128.685 -169.835 ;
        RECT 128.355 -171.525 128.685 -171.195 ;
        RECT 128.355 -172.885 128.685 -172.555 ;
        RECT 128.355 -174.245 128.685 -173.915 ;
        RECT 128.355 -175.605 128.685 -175.275 ;
        RECT 128.355 -176.965 128.685 -176.635 ;
        RECT 128.355 -178.325 128.685 -177.995 ;
        RECT 128.355 -179.685 128.685 -179.355 ;
        RECT 128.355 -181.045 128.685 -180.715 ;
        RECT 128.355 -182.405 128.685 -182.075 ;
        RECT 128.355 -183.765 128.685 -183.435 ;
        RECT 128.355 -185.125 128.685 -184.795 ;
        RECT 128.355 -186.485 128.685 -186.155 ;
        RECT 128.355 -187.845 128.685 -187.515 ;
        RECT 128.355 -189.205 128.685 -188.875 ;
        RECT 128.355 -190.565 128.685 -190.235 ;
        RECT 128.355 -191.925 128.685 -191.595 ;
        RECT 128.355 -193.285 128.685 -192.955 ;
        RECT 128.355 -194.645 128.685 -194.315 ;
        RECT 128.355 -196.005 128.685 -195.675 ;
        RECT 128.355 -197.365 128.685 -197.035 ;
        RECT 128.355 -198.725 128.685 -198.395 ;
        RECT 128.355 -200.085 128.685 -199.755 ;
        RECT 128.355 -201.445 128.685 -201.115 ;
        RECT 128.355 -202.805 128.685 -202.475 ;
        RECT 128.355 -204.165 128.685 -203.835 ;
        RECT 128.355 -205.525 128.685 -205.195 ;
        RECT 128.355 -206.885 128.685 -206.555 ;
        RECT 128.355 -208.245 128.685 -207.915 ;
        RECT 128.355 -209.605 128.685 -209.275 ;
        RECT 128.355 -210.965 128.685 -210.635 ;
        RECT 128.355 -212.325 128.685 -211.995 ;
        RECT 128.355 -213.685 128.685 -213.355 ;
        RECT 128.355 -215.045 128.685 -214.715 ;
        RECT 128.355 -216.405 128.685 -216.075 ;
        RECT 128.355 -217.765 128.685 -217.435 ;
        RECT 128.355 -219.125 128.685 -218.795 ;
        RECT 128.355 -221.37 128.685 -220.24 ;
        RECT 128.36 -221.485 128.68 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.715 129.8 130.045 130.93 ;
        RECT 129.715 127.675 130.045 128.005 ;
        RECT 129.715 126.315 130.045 126.645 ;
        RECT 129.715 124.955 130.045 125.285 ;
        RECT 129.715 123.595 130.045 123.925 ;
        RECT 129.72 123.595 130.04 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.715 -1.525 130.045 -1.195 ;
        RECT 129.715 -2.885 130.045 -2.555 ;
        RECT 129.72 -3.56 130.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.715 -118.485 130.045 -118.155 ;
        RECT 129.715 -119.845 130.045 -119.515 ;
        RECT 129.715 -121.205 130.045 -120.875 ;
        RECT 129.715 -122.565 130.045 -122.235 ;
        RECT 129.715 -123.925 130.045 -123.595 ;
        RECT 129.715 -125.285 130.045 -124.955 ;
        RECT 129.715 -126.645 130.045 -126.315 ;
        RECT 129.715 -128.005 130.045 -127.675 ;
        RECT 129.715 -129.365 130.045 -129.035 ;
        RECT 129.715 -130.725 130.045 -130.395 ;
        RECT 129.715 -132.085 130.045 -131.755 ;
        RECT 129.715 -133.445 130.045 -133.115 ;
        RECT 129.715 -134.805 130.045 -134.475 ;
        RECT 129.715 -136.165 130.045 -135.835 ;
        RECT 129.715 -137.525 130.045 -137.195 ;
        RECT 129.715 -138.885 130.045 -138.555 ;
        RECT 129.715 -140.245 130.045 -139.915 ;
        RECT 129.715 -141.605 130.045 -141.275 ;
        RECT 129.715 -142.965 130.045 -142.635 ;
        RECT 129.715 -144.325 130.045 -143.995 ;
        RECT 129.715 -145.685 130.045 -145.355 ;
        RECT 129.715 -147.045 130.045 -146.715 ;
        RECT 129.715 -148.405 130.045 -148.075 ;
        RECT 129.715 -149.765 130.045 -149.435 ;
        RECT 129.715 -151.125 130.045 -150.795 ;
        RECT 129.715 -152.485 130.045 -152.155 ;
        RECT 129.715 -153.845 130.045 -153.515 ;
        RECT 129.715 -155.205 130.045 -154.875 ;
        RECT 129.715 -156.565 130.045 -156.235 ;
        RECT 129.715 -157.925 130.045 -157.595 ;
        RECT 129.715 -159.285 130.045 -158.955 ;
        RECT 129.715 -160.645 130.045 -160.315 ;
        RECT 129.715 -162.005 130.045 -161.675 ;
        RECT 129.715 -163.365 130.045 -163.035 ;
        RECT 129.715 -164.725 130.045 -164.395 ;
        RECT 129.715 -166.085 130.045 -165.755 ;
        RECT 129.715 -167.445 130.045 -167.115 ;
        RECT 129.715 -168.805 130.045 -168.475 ;
        RECT 129.715 -170.165 130.045 -169.835 ;
        RECT 129.715 -171.525 130.045 -171.195 ;
        RECT 129.715 -172.885 130.045 -172.555 ;
        RECT 129.715 -174.245 130.045 -173.915 ;
        RECT 129.715 -175.605 130.045 -175.275 ;
        RECT 129.715 -176.965 130.045 -176.635 ;
        RECT 129.715 -178.325 130.045 -177.995 ;
        RECT 129.715 -179.685 130.045 -179.355 ;
        RECT 129.715 -181.045 130.045 -180.715 ;
        RECT 129.715 -182.405 130.045 -182.075 ;
        RECT 129.715 -183.765 130.045 -183.435 ;
        RECT 129.715 -185.125 130.045 -184.795 ;
        RECT 129.715 -186.485 130.045 -186.155 ;
        RECT 129.715 -187.845 130.045 -187.515 ;
        RECT 129.715 -189.205 130.045 -188.875 ;
        RECT 129.715 -190.565 130.045 -190.235 ;
        RECT 129.715 -191.925 130.045 -191.595 ;
        RECT 129.715 -193.285 130.045 -192.955 ;
        RECT 129.715 -194.645 130.045 -194.315 ;
        RECT 129.715 -196.005 130.045 -195.675 ;
        RECT 129.715 -197.365 130.045 -197.035 ;
        RECT 129.715 -198.725 130.045 -198.395 ;
        RECT 129.715 -200.085 130.045 -199.755 ;
        RECT 129.715 -201.445 130.045 -201.115 ;
        RECT 129.715 -202.805 130.045 -202.475 ;
        RECT 129.715 -204.165 130.045 -203.835 ;
        RECT 129.715 -205.525 130.045 -205.195 ;
        RECT 129.715 -206.885 130.045 -206.555 ;
        RECT 129.715 -208.245 130.045 -207.915 ;
        RECT 129.715 -209.605 130.045 -209.275 ;
        RECT 129.715 -210.965 130.045 -210.635 ;
        RECT 129.715 -212.325 130.045 -211.995 ;
        RECT 129.715 -213.685 130.045 -213.355 ;
        RECT 129.715 -215.045 130.045 -214.715 ;
        RECT 129.715 -216.405 130.045 -216.075 ;
        RECT 129.715 -217.765 130.045 -217.435 ;
        RECT 129.715 -219.125 130.045 -218.795 ;
        RECT 129.715 -221.37 130.045 -220.24 ;
        RECT 129.72 -221.485 130.04 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.075 129.8 131.405 130.93 ;
        RECT 131.075 127.675 131.405 128.005 ;
        RECT 131.075 126.315 131.405 126.645 ;
        RECT 131.075 124.955 131.405 125.285 ;
        RECT 131.075 123.595 131.405 123.925 ;
        RECT 131.08 123.595 131.4 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.075 -122.565 131.405 -122.235 ;
        RECT 131.075 -123.925 131.405 -123.595 ;
        RECT 131.075 -125.285 131.405 -124.955 ;
        RECT 131.075 -126.645 131.405 -126.315 ;
        RECT 131.075 -128.005 131.405 -127.675 ;
        RECT 131.075 -129.365 131.405 -129.035 ;
        RECT 131.075 -130.725 131.405 -130.395 ;
        RECT 131.075 -132.085 131.405 -131.755 ;
        RECT 131.075 -133.445 131.405 -133.115 ;
        RECT 131.075 -134.805 131.405 -134.475 ;
        RECT 131.075 -136.165 131.405 -135.835 ;
        RECT 131.075 -137.525 131.405 -137.195 ;
        RECT 131.075 -138.885 131.405 -138.555 ;
        RECT 131.075 -140.245 131.405 -139.915 ;
        RECT 131.075 -141.605 131.405 -141.275 ;
        RECT 131.075 -142.965 131.405 -142.635 ;
        RECT 131.075 -144.325 131.405 -143.995 ;
        RECT 131.075 -145.685 131.405 -145.355 ;
        RECT 131.075 -147.045 131.405 -146.715 ;
        RECT 131.075 -148.405 131.405 -148.075 ;
        RECT 131.075 -149.765 131.405 -149.435 ;
        RECT 131.075 -151.125 131.405 -150.795 ;
        RECT 131.075 -152.485 131.405 -152.155 ;
        RECT 131.075 -153.845 131.405 -153.515 ;
        RECT 131.075 -155.205 131.405 -154.875 ;
        RECT 131.075 -156.565 131.405 -156.235 ;
        RECT 131.075 -157.925 131.405 -157.595 ;
        RECT 131.075 -159.285 131.405 -158.955 ;
        RECT 131.075 -160.645 131.405 -160.315 ;
        RECT 131.075 -162.005 131.405 -161.675 ;
        RECT 131.075 -163.365 131.405 -163.035 ;
        RECT 131.075 -164.725 131.405 -164.395 ;
        RECT 131.075 -166.085 131.405 -165.755 ;
        RECT 131.075 -167.445 131.405 -167.115 ;
        RECT 131.075 -168.805 131.405 -168.475 ;
        RECT 131.075 -170.165 131.405 -169.835 ;
        RECT 131.075 -171.525 131.405 -171.195 ;
        RECT 131.075 -172.885 131.405 -172.555 ;
        RECT 131.075 -174.245 131.405 -173.915 ;
        RECT 131.075 -175.605 131.405 -175.275 ;
        RECT 131.075 -176.965 131.405 -176.635 ;
        RECT 131.075 -178.325 131.405 -177.995 ;
        RECT 131.075 -179.685 131.405 -179.355 ;
        RECT 131.075 -181.045 131.405 -180.715 ;
        RECT 131.075 -182.405 131.405 -182.075 ;
        RECT 131.075 -183.765 131.405 -183.435 ;
        RECT 131.075 -185.125 131.405 -184.795 ;
        RECT 131.075 -186.485 131.405 -186.155 ;
        RECT 131.075 -187.845 131.405 -187.515 ;
        RECT 131.075 -189.205 131.405 -188.875 ;
        RECT 131.075 -190.565 131.405 -190.235 ;
        RECT 131.075 -191.925 131.405 -191.595 ;
        RECT 131.075 -193.285 131.405 -192.955 ;
        RECT 131.075 -194.645 131.405 -194.315 ;
        RECT 131.075 -196.005 131.405 -195.675 ;
        RECT 131.075 -197.365 131.405 -197.035 ;
        RECT 131.075 -198.725 131.405 -198.395 ;
        RECT 131.075 -200.085 131.405 -199.755 ;
        RECT 131.075 -201.445 131.405 -201.115 ;
        RECT 131.075 -202.805 131.405 -202.475 ;
        RECT 131.075 -204.165 131.405 -203.835 ;
        RECT 131.075 -205.525 131.405 -205.195 ;
        RECT 131.075 -206.885 131.405 -206.555 ;
        RECT 131.075 -208.245 131.405 -207.915 ;
        RECT 131.075 -209.605 131.405 -209.275 ;
        RECT 131.075 -210.965 131.405 -210.635 ;
        RECT 131.075 -212.325 131.405 -211.995 ;
        RECT 131.075 -213.685 131.405 -213.355 ;
        RECT 131.075 -215.045 131.405 -214.715 ;
        RECT 131.075 -216.405 131.405 -216.075 ;
        RECT 131.075 -217.765 131.405 -217.435 ;
        RECT 131.075 -219.125 131.405 -218.795 ;
        RECT 131.075 -221.37 131.405 -220.24 ;
        RECT 131.08 -221.485 131.4 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.41 -121.535 131.74 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.435 129.8 132.765 130.93 ;
        RECT 132.435 127.675 132.765 128.005 ;
        RECT 132.435 126.315 132.765 126.645 ;
        RECT 132.435 124.955 132.765 125.285 ;
        RECT 132.435 123.595 132.765 123.925 ;
        RECT 132.44 123.595 132.76 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.435 -1.525 132.765 -1.195 ;
        RECT 132.435 -2.885 132.765 -2.555 ;
        RECT 132.44 -3.56 132.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.795 129.8 134.125 130.93 ;
        RECT 133.795 127.675 134.125 128.005 ;
        RECT 133.795 126.315 134.125 126.645 ;
        RECT 133.795 124.955 134.125 125.285 ;
        RECT 133.795 123.595 134.125 123.925 ;
        RECT 133.8 123.595 134.12 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.795 -1.525 134.125 -1.195 ;
        RECT 133.795 -2.885 134.125 -2.555 ;
        RECT 133.8 -3.56 134.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.155 129.8 135.485 130.93 ;
        RECT 135.155 127.675 135.485 128.005 ;
        RECT 135.155 126.315 135.485 126.645 ;
        RECT 135.155 124.955 135.485 125.285 ;
        RECT 135.155 123.595 135.485 123.925 ;
        RECT 135.16 123.595 135.48 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.155 -1.525 135.485 -1.195 ;
        RECT 135.155 -2.885 135.485 -2.555 ;
        RECT 135.16 -3.56 135.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.155 -198.725 135.485 -198.395 ;
        RECT 135.155 -200.085 135.485 -199.755 ;
        RECT 135.155 -201.445 135.485 -201.115 ;
        RECT 135.155 -202.805 135.485 -202.475 ;
        RECT 135.155 -204.165 135.485 -203.835 ;
        RECT 135.155 -205.525 135.485 -205.195 ;
        RECT 135.155 -206.885 135.485 -206.555 ;
        RECT 135.155 -208.245 135.485 -207.915 ;
        RECT 135.155 -209.605 135.485 -209.275 ;
        RECT 135.155 -210.965 135.485 -210.635 ;
        RECT 135.155 -212.325 135.485 -211.995 ;
        RECT 135.155 -213.685 135.485 -213.355 ;
        RECT 135.155 -215.045 135.485 -214.715 ;
        RECT 135.155 -216.405 135.485 -216.075 ;
        RECT 135.155 -217.765 135.485 -217.435 ;
        RECT 135.155 -219.125 135.485 -218.795 ;
        RECT 135.155 -221.37 135.485 -220.24 ;
        RECT 135.16 -221.485 135.48 -118.155 ;
        RECT 135.155 -118.485 135.485 -118.155 ;
        RECT 135.155 -119.845 135.485 -119.515 ;
        RECT 135.155 -121.205 135.485 -120.875 ;
        RECT 135.155 -122.565 135.485 -122.235 ;
        RECT 135.155 -123.925 135.485 -123.595 ;
        RECT 135.155 -125.285 135.485 -124.955 ;
        RECT 135.155 -126.645 135.485 -126.315 ;
        RECT 135.155 -128.005 135.485 -127.675 ;
        RECT 135.155 -129.365 135.485 -129.035 ;
        RECT 135.155 -130.725 135.485 -130.395 ;
        RECT 135.155 -132.085 135.485 -131.755 ;
        RECT 135.155 -133.445 135.485 -133.115 ;
        RECT 135.155 -134.805 135.485 -134.475 ;
        RECT 135.155 -136.165 135.485 -135.835 ;
        RECT 135.155 -137.525 135.485 -137.195 ;
        RECT 135.155 -138.885 135.485 -138.555 ;
        RECT 135.155 -140.245 135.485 -139.915 ;
        RECT 135.155 -141.605 135.485 -141.275 ;
        RECT 135.155 -142.965 135.485 -142.635 ;
        RECT 135.155 -144.325 135.485 -143.995 ;
        RECT 135.155 -145.685 135.485 -145.355 ;
        RECT 135.155 -147.045 135.485 -146.715 ;
        RECT 135.155 -148.405 135.485 -148.075 ;
        RECT 135.155 -149.765 135.485 -149.435 ;
        RECT 135.155 -151.125 135.485 -150.795 ;
        RECT 135.155 -152.485 135.485 -152.155 ;
        RECT 135.155 -153.845 135.485 -153.515 ;
        RECT 135.155 -155.205 135.485 -154.875 ;
        RECT 135.155 -156.565 135.485 -156.235 ;
        RECT 135.155 -157.925 135.485 -157.595 ;
        RECT 135.155 -159.285 135.485 -158.955 ;
        RECT 135.155 -160.645 135.485 -160.315 ;
        RECT 135.155 -162.005 135.485 -161.675 ;
        RECT 135.155 -163.365 135.485 -163.035 ;
        RECT 135.155 -164.725 135.485 -164.395 ;
        RECT 135.155 -166.085 135.485 -165.755 ;
        RECT 135.155 -167.445 135.485 -167.115 ;
        RECT 135.155 -168.805 135.485 -168.475 ;
        RECT 135.155 -170.165 135.485 -169.835 ;
        RECT 135.155 -171.525 135.485 -171.195 ;
        RECT 135.155 -172.885 135.485 -172.555 ;
        RECT 135.155 -174.245 135.485 -173.915 ;
        RECT 135.155 -175.605 135.485 -175.275 ;
        RECT 135.155 -176.965 135.485 -176.635 ;
        RECT 135.155 -178.325 135.485 -177.995 ;
        RECT 135.155 -179.685 135.485 -179.355 ;
        RECT 135.155 -181.045 135.485 -180.715 ;
        RECT 135.155 -182.405 135.485 -182.075 ;
        RECT 135.155 -183.765 135.485 -183.435 ;
        RECT 135.155 -185.125 135.485 -184.795 ;
        RECT 135.155 -186.485 135.485 -186.155 ;
        RECT 135.155 -187.845 135.485 -187.515 ;
        RECT 135.155 -189.205 135.485 -188.875 ;
        RECT 135.155 -190.565 135.485 -190.235 ;
        RECT 135.155 -191.925 135.485 -191.595 ;
        RECT 135.155 -193.285 135.485 -192.955 ;
        RECT 135.155 -194.645 135.485 -194.315 ;
        RECT 135.155 -196.005 135.485 -195.675 ;
        RECT 135.155 -197.365 135.485 -197.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.395 129.8 79.725 130.93 ;
        RECT 79.395 127.675 79.725 128.005 ;
        RECT 79.395 126.315 79.725 126.645 ;
        RECT 79.395 124.955 79.725 125.285 ;
        RECT 79.395 123.595 79.725 123.925 ;
        RECT 79.4 123.595 79.72 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.395 -1.525 79.725 -1.195 ;
        RECT 79.395 -2.885 79.725 -2.555 ;
        RECT 79.4 -3.56 79.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.755 129.8 81.085 130.93 ;
        RECT 80.755 127.675 81.085 128.005 ;
        RECT 80.755 126.315 81.085 126.645 ;
        RECT 80.755 124.955 81.085 125.285 ;
        RECT 80.755 123.595 81.085 123.925 ;
        RECT 80.76 123.595 81.08 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.755 -1.525 81.085 -1.195 ;
        RECT 80.755 -2.885 81.085 -2.555 ;
        RECT 80.76 -3.56 81.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.755 -118.485 81.085 -118.155 ;
        RECT 80.755 -119.845 81.085 -119.515 ;
        RECT 80.755 -121.205 81.085 -120.875 ;
        RECT 80.755 -122.565 81.085 -122.235 ;
        RECT 80.755 -123.925 81.085 -123.595 ;
        RECT 80.755 -125.285 81.085 -124.955 ;
        RECT 80.755 -126.645 81.085 -126.315 ;
        RECT 80.755 -128.005 81.085 -127.675 ;
        RECT 80.755 -129.365 81.085 -129.035 ;
        RECT 80.755 -130.725 81.085 -130.395 ;
        RECT 80.755 -132.085 81.085 -131.755 ;
        RECT 80.755 -133.445 81.085 -133.115 ;
        RECT 80.755 -134.805 81.085 -134.475 ;
        RECT 80.755 -136.165 81.085 -135.835 ;
        RECT 80.755 -137.525 81.085 -137.195 ;
        RECT 80.755 -138.885 81.085 -138.555 ;
        RECT 80.755 -140.245 81.085 -139.915 ;
        RECT 80.755 -141.605 81.085 -141.275 ;
        RECT 80.755 -142.965 81.085 -142.635 ;
        RECT 80.755 -144.325 81.085 -143.995 ;
        RECT 80.755 -145.685 81.085 -145.355 ;
        RECT 80.755 -147.045 81.085 -146.715 ;
        RECT 80.755 -148.405 81.085 -148.075 ;
        RECT 80.755 -149.765 81.085 -149.435 ;
        RECT 80.755 -151.125 81.085 -150.795 ;
        RECT 80.755 -152.485 81.085 -152.155 ;
        RECT 80.755 -153.845 81.085 -153.515 ;
        RECT 80.755 -155.205 81.085 -154.875 ;
        RECT 80.755 -156.565 81.085 -156.235 ;
        RECT 80.755 -157.925 81.085 -157.595 ;
        RECT 80.755 -159.285 81.085 -158.955 ;
        RECT 80.755 -160.645 81.085 -160.315 ;
        RECT 80.755 -162.005 81.085 -161.675 ;
        RECT 80.755 -163.365 81.085 -163.035 ;
        RECT 80.755 -164.725 81.085 -164.395 ;
        RECT 80.755 -166.085 81.085 -165.755 ;
        RECT 80.755 -167.445 81.085 -167.115 ;
        RECT 80.755 -168.805 81.085 -168.475 ;
        RECT 80.755 -170.165 81.085 -169.835 ;
        RECT 80.755 -171.525 81.085 -171.195 ;
        RECT 80.755 -172.885 81.085 -172.555 ;
        RECT 80.755 -174.245 81.085 -173.915 ;
        RECT 80.755 -175.605 81.085 -175.275 ;
        RECT 80.755 -176.965 81.085 -176.635 ;
        RECT 80.755 -178.325 81.085 -177.995 ;
        RECT 80.755 -179.685 81.085 -179.355 ;
        RECT 80.755 -181.045 81.085 -180.715 ;
        RECT 80.755 -182.405 81.085 -182.075 ;
        RECT 80.755 -183.765 81.085 -183.435 ;
        RECT 80.755 -185.125 81.085 -184.795 ;
        RECT 80.755 -186.485 81.085 -186.155 ;
        RECT 80.755 -187.845 81.085 -187.515 ;
        RECT 80.755 -189.205 81.085 -188.875 ;
        RECT 80.755 -190.565 81.085 -190.235 ;
        RECT 80.755 -191.925 81.085 -191.595 ;
        RECT 80.755 -193.285 81.085 -192.955 ;
        RECT 80.755 -194.645 81.085 -194.315 ;
        RECT 80.755 -196.005 81.085 -195.675 ;
        RECT 80.755 -197.365 81.085 -197.035 ;
        RECT 80.755 -198.725 81.085 -198.395 ;
        RECT 80.755 -200.085 81.085 -199.755 ;
        RECT 80.755 -201.445 81.085 -201.115 ;
        RECT 80.755 -202.805 81.085 -202.475 ;
        RECT 80.755 -204.165 81.085 -203.835 ;
        RECT 80.755 -205.525 81.085 -205.195 ;
        RECT 80.755 -206.885 81.085 -206.555 ;
        RECT 80.755 -208.245 81.085 -207.915 ;
        RECT 80.755 -209.605 81.085 -209.275 ;
        RECT 80.755 -210.965 81.085 -210.635 ;
        RECT 80.755 -212.325 81.085 -211.995 ;
        RECT 80.755 -213.685 81.085 -213.355 ;
        RECT 80.755 -215.045 81.085 -214.715 ;
        RECT 80.755 -216.405 81.085 -216.075 ;
        RECT 80.755 -217.765 81.085 -217.435 ;
        RECT 80.755 -219.125 81.085 -218.795 ;
        RECT 80.755 -221.37 81.085 -220.24 ;
        RECT 80.76 -221.485 81.08 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.115 129.8 82.445 130.93 ;
        RECT 82.115 127.675 82.445 128.005 ;
        RECT 82.115 126.315 82.445 126.645 ;
        RECT 82.115 124.955 82.445 125.285 ;
        RECT 82.115 123.595 82.445 123.925 ;
        RECT 82.12 123.595 82.44 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.115 -122.565 82.445 -122.235 ;
        RECT 82.115 -123.925 82.445 -123.595 ;
        RECT 82.115 -125.285 82.445 -124.955 ;
        RECT 82.115 -126.645 82.445 -126.315 ;
        RECT 82.115 -128.005 82.445 -127.675 ;
        RECT 82.115 -129.365 82.445 -129.035 ;
        RECT 82.115 -130.725 82.445 -130.395 ;
        RECT 82.115 -132.085 82.445 -131.755 ;
        RECT 82.115 -133.445 82.445 -133.115 ;
        RECT 82.115 -134.805 82.445 -134.475 ;
        RECT 82.115 -136.165 82.445 -135.835 ;
        RECT 82.115 -137.525 82.445 -137.195 ;
        RECT 82.115 -138.885 82.445 -138.555 ;
        RECT 82.115 -140.245 82.445 -139.915 ;
        RECT 82.115 -141.605 82.445 -141.275 ;
        RECT 82.115 -142.965 82.445 -142.635 ;
        RECT 82.115 -144.325 82.445 -143.995 ;
        RECT 82.115 -145.685 82.445 -145.355 ;
        RECT 82.115 -147.045 82.445 -146.715 ;
        RECT 82.115 -148.405 82.445 -148.075 ;
        RECT 82.115 -149.765 82.445 -149.435 ;
        RECT 82.115 -151.125 82.445 -150.795 ;
        RECT 82.115 -152.485 82.445 -152.155 ;
        RECT 82.115 -153.845 82.445 -153.515 ;
        RECT 82.115 -155.205 82.445 -154.875 ;
        RECT 82.115 -156.565 82.445 -156.235 ;
        RECT 82.115 -157.925 82.445 -157.595 ;
        RECT 82.115 -159.285 82.445 -158.955 ;
        RECT 82.115 -160.645 82.445 -160.315 ;
        RECT 82.115 -162.005 82.445 -161.675 ;
        RECT 82.115 -163.365 82.445 -163.035 ;
        RECT 82.115 -164.725 82.445 -164.395 ;
        RECT 82.115 -166.085 82.445 -165.755 ;
        RECT 82.115 -167.445 82.445 -167.115 ;
        RECT 82.115 -168.805 82.445 -168.475 ;
        RECT 82.115 -170.165 82.445 -169.835 ;
        RECT 82.115 -171.525 82.445 -171.195 ;
        RECT 82.115 -172.885 82.445 -172.555 ;
        RECT 82.115 -174.245 82.445 -173.915 ;
        RECT 82.115 -175.605 82.445 -175.275 ;
        RECT 82.115 -176.965 82.445 -176.635 ;
        RECT 82.115 -178.325 82.445 -177.995 ;
        RECT 82.115 -179.685 82.445 -179.355 ;
        RECT 82.115 -181.045 82.445 -180.715 ;
        RECT 82.115 -182.405 82.445 -182.075 ;
        RECT 82.115 -183.765 82.445 -183.435 ;
        RECT 82.115 -185.125 82.445 -184.795 ;
        RECT 82.115 -186.485 82.445 -186.155 ;
        RECT 82.115 -187.845 82.445 -187.515 ;
        RECT 82.115 -189.205 82.445 -188.875 ;
        RECT 82.115 -190.565 82.445 -190.235 ;
        RECT 82.115 -191.925 82.445 -191.595 ;
        RECT 82.115 -193.285 82.445 -192.955 ;
        RECT 82.115 -194.645 82.445 -194.315 ;
        RECT 82.115 -196.005 82.445 -195.675 ;
        RECT 82.115 -197.365 82.445 -197.035 ;
        RECT 82.115 -198.725 82.445 -198.395 ;
        RECT 82.115 -200.085 82.445 -199.755 ;
        RECT 82.115 -201.445 82.445 -201.115 ;
        RECT 82.115 -202.805 82.445 -202.475 ;
        RECT 82.115 -204.165 82.445 -203.835 ;
        RECT 82.115 -205.525 82.445 -205.195 ;
        RECT 82.115 -206.885 82.445 -206.555 ;
        RECT 82.115 -208.245 82.445 -207.915 ;
        RECT 82.115 -209.605 82.445 -209.275 ;
        RECT 82.115 -210.965 82.445 -210.635 ;
        RECT 82.115 -212.325 82.445 -211.995 ;
        RECT 82.115 -213.685 82.445 -213.355 ;
        RECT 82.115 -215.045 82.445 -214.715 ;
        RECT 82.115 -216.405 82.445 -216.075 ;
        RECT 82.115 -217.765 82.445 -217.435 ;
        RECT 82.115 -219.125 82.445 -218.795 ;
        RECT 82.115 -221.37 82.445 -220.24 ;
        RECT 82.12 -221.485 82.44 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.61 -121.535 82.94 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.475 129.8 83.805 130.93 ;
        RECT 83.475 127.675 83.805 128.005 ;
        RECT 83.475 126.315 83.805 126.645 ;
        RECT 83.475 124.955 83.805 125.285 ;
        RECT 83.475 123.595 83.805 123.925 ;
        RECT 83.48 123.595 83.8 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.475 -1.525 83.805 -1.195 ;
        RECT 83.475 -2.885 83.805 -2.555 ;
        RECT 83.48 -3.56 83.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.835 129.8 85.165 130.93 ;
        RECT 84.835 127.675 85.165 128.005 ;
        RECT 84.835 126.315 85.165 126.645 ;
        RECT 84.835 124.955 85.165 125.285 ;
        RECT 84.835 123.595 85.165 123.925 ;
        RECT 84.84 123.595 85.16 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.835 -1.525 85.165 -1.195 ;
        RECT 84.835 -2.885 85.165 -2.555 ;
        RECT 84.84 -3.56 85.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.195 129.8 86.525 130.93 ;
        RECT 86.195 127.675 86.525 128.005 ;
        RECT 86.195 126.315 86.525 126.645 ;
        RECT 86.195 124.955 86.525 125.285 ;
        RECT 86.195 123.595 86.525 123.925 ;
        RECT 86.2 123.595 86.52 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.195 -1.525 86.525 -1.195 ;
        RECT 86.195 -2.885 86.525 -2.555 ;
        RECT 86.2 -3.56 86.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.195 -118.485 86.525 -118.155 ;
        RECT 86.195 -119.845 86.525 -119.515 ;
        RECT 86.195 -121.205 86.525 -120.875 ;
        RECT 86.195 -122.565 86.525 -122.235 ;
        RECT 86.195 -123.925 86.525 -123.595 ;
        RECT 86.195 -125.285 86.525 -124.955 ;
        RECT 86.195 -126.645 86.525 -126.315 ;
        RECT 86.195 -128.005 86.525 -127.675 ;
        RECT 86.195 -129.365 86.525 -129.035 ;
        RECT 86.195 -130.725 86.525 -130.395 ;
        RECT 86.195 -132.085 86.525 -131.755 ;
        RECT 86.195 -133.445 86.525 -133.115 ;
        RECT 86.195 -134.805 86.525 -134.475 ;
        RECT 86.195 -136.165 86.525 -135.835 ;
        RECT 86.195 -137.525 86.525 -137.195 ;
        RECT 86.195 -138.885 86.525 -138.555 ;
        RECT 86.195 -140.245 86.525 -139.915 ;
        RECT 86.195 -141.605 86.525 -141.275 ;
        RECT 86.195 -142.965 86.525 -142.635 ;
        RECT 86.195 -144.325 86.525 -143.995 ;
        RECT 86.195 -145.685 86.525 -145.355 ;
        RECT 86.195 -147.045 86.525 -146.715 ;
        RECT 86.195 -148.405 86.525 -148.075 ;
        RECT 86.195 -149.765 86.525 -149.435 ;
        RECT 86.195 -151.125 86.525 -150.795 ;
        RECT 86.195 -152.485 86.525 -152.155 ;
        RECT 86.195 -153.845 86.525 -153.515 ;
        RECT 86.195 -155.205 86.525 -154.875 ;
        RECT 86.195 -156.565 86.525 -156.235 ;
        RECT 86.195 -157.925 86.525 -157.595 ;
        RECT 86.195 -159.285 86.525 -158.955 ;
        RECT 86.195 -160.645 86.525 -160.315 ;
        RECT 86.195 -162.005 86.525 -161.675 ;
        RECT 86.195 -163.365 86.525 -163.035 ;
        RECT 86.195 -164.725 86.525 -164.395 ;
        RECT 86.195 -166.085 86.525 -165.755 ;
        RECT 86.195 -167.445 86.525 -167.115 ;
        RECT 86.195 -168.805 86.525 -168.475 ;
        RECT 86.195 -170.165 86.525 -169.835 ;
        RECT 86.195 -171.525 86.525 -171.195 ;
        RECT 86.195 -172.885 86.525 -172.555 ;
        RECT 86.195 -174.245 86.525 -173.915 ;
        RECT 86.195 -175.605 86.525 -175.275 ;
        RECT 86.195 -176.965 86.525 -176.635 ;
        RECT 86.195 -178.325 86.525 -177.995 ;
        RECT 86.195 -179.685 86.525 -179.355 ;
        RECT 86.195 -181.045 86.525 -180.715 ;
        RECT 86.195 -182.405 86.525 -182.075 ;
        RECT 86.195 -183.765 86.525 -183.435 ;
        RECT 86.195 -185.125 86.525 -184.795 ;
        RECT 86.195 -186.485 86.525 -186.155 ;
        RECT 86.195 -187.845 86.525 -187.515 ;
        RECT 86.195 -189.205 86.525 -188.875 ;
        RECT 86.195 -190.565 86.525 -190.235 ;
        RECT 86.195 -191.925 86.525 -191.595 ;
        RECT 86.195 -193.285 86.525 -192.955 ;
        RECT 86.195 -194.645 86.525 -194.315 ;
        RECT 86.195 -196.005 86.525 -195.675 ;
        RECT 86.195 -197.365 86.525 -197.035 ;
        RECT 86.195 -198.725 86.525 -198.395 ;
        RECT 86.195 -200.085 86.525 -199.755 ;
        RECT 86.195 -201.445 86.525 -201.115 ;
        RECT 86.195 -202.805 86.525 -202.475 ;
        RECT 86.195 -204.165 86.525 -203.835 ;
        RECT 86.195 -205.525 86.525 -205.195 ;
        RECT 86.195 -206.885 86.525 -206.555 ;
        RECT 86.195 -208.245 86.525 -207.915 ;
        RECT 86.195 -209.605 86.525 -209.275 ;
        RECT 86.195 -210.965 86.525 -210.635 ;
        RECT 86.195 -212.325 86.525 -211.995 ;
        RECT 86.195 -213.685 86.525 -213.355 ;
        RECT 86.195 -215.045 86.525 -214.715 ;
        RECT 86.195 -216.405 86.525 -216.075 ;
        RECT 86.195 -217.765 86.525 -217.435 ;
        RECT 86.195 -219.125 86.525 -218.795 ;
        RECT 86.195 -221.37 86.525 -220.24 ;
        RECT 86.2 -221.485 86.52 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.555 129.8 87.885 130.93 ;
        RECT 87.555 127.675 87.885 128.005 ;
        RECT 87.555 126.315 87.885 126.645 ;
        RECT 87.555 124.955 87.885 125.285 ;
        RECT 87.555 123.595 87.885 123.925 ;
        RECT 87.56 123.595 87.88 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.555 -122.565 87.885 -122.235 ;
        RECT 87.555 -123.925 87.885 -123.595 ;
        RECT 87.555 -125.285 87.885 -124.955 ;
        RECT 87.555 -126.645 87.885 -126.315 ;
        RECT 87.555 -128.005 87.885 -127.675 ;
        RECT 87.555 -129.365 87.885 -129.035 ;
        RECT 87.555 -130.725 87.885 -130.395 ;
        RECT 87.555 -132.085 87.885 -131.755 ;
        RECT 87.555 -133.445 87.885 -133.115 ;
        RECT 87.555 -134.805 87.885 -134.475 ;
        RECT 87.555 -136.165 87.885 -135.835 ;
        RECT 87.555 -137.525 87.885 -137.195 ;
        RECT 87.555 -138.885 87.885 -138.555 ;
        RECT 87.555 -140.245 87.885 -139.915 ;
        RECT 87.555 -141.605 87.885 -141.275 ;
        RECT 87.555 -142.965 87.885 -142.635 ;
        RECT 87.555 -144.325 87.885 -143.995 ;
        RECT 87.555 -145.685 87.885 -145.355 ;
        RECT 87.555 -147.045 87.885 -146.715 ;
        RECT 87.555 -148.405 87.885 -148.075 ;
        RECT 87.555 -149.765 87.885 -149.435 ;
        RECT 87.555 -151.125 87.885 -150.795 ;
        RECT 87.555 -152.485 87.885 -152.155 ;
        RECT 87.555 -153.845 87.885 -153.515 ;
        RECT 87.555 -155.205 87.885 -154.875 ;
        RECT 87.555 -156.565 87.885 -156.235 ;
        RECT 87.555 -157.925 87.885 -157.595 ;
        RECT 87.555 -159.285 87.885 -158.955 ;
        RECT 87.555 -160.645 87.885 -160.315 ;
        RECT 87.555 -162.005 87.885 -161.675 ;
        RECT 87.555 -163.365 87.885 -163.035 ;
        RECT 87.555 -164.725 87.885 -164.395 ;
        RECT 87.555 -166.085 87.885 -165.755 ;
        RECT 87.555 -167.445 87.885 -167.115 ;
        RECT 87.555 -168.805 87.885 -168.475 ;
        RECT 87.555 -170.165 87.885 -169.835 ;
        RECT 87.555 -171.525 87.885 -171.195 ;
        RECT 87.555 -172.885 87.885 -172.555 ;
        RECT 87.555 -174.245 87.885 -173.915 ;
        RECT 87.555 -175.605 87.885 -175.275 ;
        RECT 87.555 -176.965 87.885 -176.635 ;
        RECT 87.555 -178.325 87.885 -177.995 ;
        RECT 87.555 -179.685 87.885 -179.355 ;
        RECT 87.555 -181.045 87.885 -180.715 ;
        RECT 87.555 -182.405 87.885 -182.075 ;
        RECT 87.555 -183.765 87.885 -183.435 ;
        RECT 87.555 -185.125 87.885 -184.795 ;
        RECT 87.555 -186.485 87.885 -186.155 ;
        RECT 87.555 -187.845 87.885 -187.515 ;
        RECT 87.555 -189.205 87.885 -188.875 ;
        RECT 87.555 -190.565 87.885 -190.235 ;
        RECT 87.555 -191.925 87.885 -191.595 ;
        RECT 87.555 -193.285 87.885 -192.955 ;
        RECT 87.555 -194.645 87.885 -194.315 ;
        RECT 87.555 -196.005 87.885 -195.675 ;
        RECT 87.555 -197.365 87.885 -197.035 ;
        RECT 87.555 -198.725 87.885 -198.395 ;
        RECT 87.555 -200.085 87.885 -199.755 ;
        RECT 87.555 -201.445 87.885 -201.115 ;
        RECT 87.555 -202.805 87.885 -202.475 ;
        RECT 87.555 -204.165 87.885 -203.835 ;
        RECT 87.555 -205.525 87.885 -205.195 ;
        RECT 87.555 -206.885 87.885 -206.555 ;
        RECT 87.555 -208.245 87.885 -207.915 ;
        RECT 87.555 -209.605 87.885 -209.275 ;
        RECT 87.555 -210.965 87.885 -210.635 ;
        RECT 87.555 -212.325 87.885 -211.995 ;
        RECT 87.555 -213.685 87.885 -213.355 ;
        RECT 87.555 -215.045 87.885 -214.715 ;
        RECT 87.555 -216.405 87.885 -216.075 ;
        RECT 87.555 -217.765 87.885 -217.435 ;
        RECT 87.555 -219.125 87.885 -218.795 ;
        RECT 87.555 -221.37 87.885 -220.24 ;
        RECT 87.56 -221.485 87.88 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.71 -121.535 89.04 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.915 129.8 89.245 130.93 ;
        RECT 88.915 127.675 89.245 128.005 ;
        RECT 88.915 126.315 89.245 126.645 ;
        RECT 88.915 124.955 89.245 125.285 ;
        RECT 88.915 123.595 89.245 123.925 ;
        RECT 88.92 123.595 89.24 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.275 129.8 90.605 130.93 ;
        RECT 90.275 127.675 90.605 128.005 ;
        RECT 90.275 126.315 90.605 126.645 ;
        RECT 90.275 124.955 90.605 125.285 ;
        RECT 90.275 123.595 90.605 123.925 ;
        RECT 90.28 123.595 90.6 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.275 -1.525 90.605 -1.195 ;
        RECT 90.275 -2.885 90.605 -2.555 ;
        RECT 90.28 -3.56 90.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.275 -118.485 90.605 -118.155 ;
        RECT 90.275 -119.845 90.605 -119.515 ;
        RECT 90.275 -121.205 90.605 -120.875 ;
        RECT 90.275 -122.565 90.605 -122.235 ;
        RECT 90.275 -123.925 90.605 -123.595 ;
        RECT 90.275 -125.285 90.605 -124.955 ;
        RECT 90.275 -126.645 90.605 -126.315 ;
        RECT 90.275 -128.005 90.605 -127.675 ;
        RECT 90.275 -129.365 90.605 -129.035 ;
        RECT 90.275 -130.725 90.605 -130.395 ;
        RECT 90.275 -132.085 90.605 -131.755 ;
        RECT 90.275 -133.445 90.605 -133.115 ;
        RECT 90.275 -134.805 90.605 -134.475 ;
        RECT 90.275 -136.165 90.605 -135.835 ;
        RECT 90.275 -137.525 90.605 -137.195 ;
        RECT 90.275 -138.885 90.605 -138.555 ;
        RECT 90.275 -140.245 90.605 -139.915 ;
        RECT 90.275 -141.605 90.605 -141.275 ;
        RECT 90.275 -142.965 90.605 -142.635 ;
        RECT 90.275 -144.325 90.605 -143.995 ;
        RECT 90.275 -145.685 90.605 -145.355 ;
        RECT 90.275 -147.045 90.605 -146.715 ;
        RECT 90.275 -148.405 90.605 -148.075 ;
        RECT 90.275 -149.765 90.605 -149.435 ;
        RECT 90.275 -151.125 90.605 -150.795 ;
        RECT 90.275 -152.485 90.605 -152.155 ;
        RECT 90.275 -153.845 90.605 -153.515 ;
        RECT 90.275 -155.205 90.605 -154.875 ;
        RECT 90.275 -156.565 90.605 -156.235 ;
        RECT 90.275 -157.925 90.605 -157.595 ;
        RECT 90.275 -159.285 90.605 -158.955 ;
        RECT 90.275 -160.645 90.605 -160.315 ;
        RECT 90.275 -162.005 90.605 -161.675 ;
        RECT 90.275 -163.365 90.605 -163.035 ;
        RECT 90.275 -164.725 90.605 -164.395 ;
        RECT 90.275 -166.085 90.605 -165.755 ;
        RECT 90.275 -167.445 90.605 -167.115 ;
        RECT 90.275 -168.805 90.605 -168.475 ;
        RECT 90.275 -170.165 90.605 -169.835 ;
        RECT 90.275 -171.525 90.605 -171.195 ;
        RECT 90.275 -172.885 90.605 -172.555 ;
        RECT 90.275 -174.245 90.605 -173.915 ;
        RECT 90.275 -175.605 90.605 -175.275 ;
        RECT 90.275 -176.965 90.605 -176.635 ;
        RECT 90.275 -178.325 90.605 -177.995 ;
        RECT 90.275 -179.685 90.605 -179.355 ;
        RECT 90.275 -181.045 90.605 -180.715 ;
        RECT 90.275 -182.405 90.605 -182.075 ;
        RECT 90.275 -183.765 90.605 -183.435 ;
        RECT 90.275 -185.125 90.605 -184.795 ;
        RECT 90.275 -186.485 90.605 -186.155 ;
        RECT 90.275 -187.845 90.605 -187.515 ;
        RECT 90.275 -189.205 90.605 -188.875 ;
        RECT 90.275 -190.565 90.605 -190.235 ;
        RECT 90.275 -191.925 90.605 -191.595 ;
        RECT 90.275 -193.285 90.605 -192.955 ;
        RECT 90.275 -194.645 90.605 -194.315 ;
        RECT 90.275 -196.005 90.605 -195.675 ;
        RECT 90.275 -197.365 90.605 -197.035 ;
        RECT 90.275 -198.725 90.605 -198.395 ;
        RECT 90.275 -200.085 90.605 -199.755 ;
        RECT 90.275 -201.445 90.605 -201.115 ;
        RECT 90.275 -202.805 90.605 -202.475 ;
        RECT 90.275 -204.165 90.605 -203.835 ;
        RECT 90.275 -205.525 90.605 -205.195 ;
        RECT 90.275 -206.885 90.605 -206.555 ;
        RECT 90.275 -208.245 90.605 -207.915 ;
        RECT 90.275 -209.605 90.605 -209.275 ;
        RECT 90.275 -210.965 90.605 -210.635 ;
        RECT 90.275 -212.325 90.605 -211.995 ;
        RECT 90.275 -213.685 90.605 -213.355 ;
        RECT 90.275 -215.045 90.605 -214.715 ;
        RECT 90.275 -216.405 90.605 -216.075 ;
        RECT 90.275 -217.765 90.605 -217.435 ;
        RECT 90.275 -219.125 90.605 -218.795 ;
        RECT 90.275 -221.37 90.605 -220.24 ;
        RECT 90.28 -221.485 90.6 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.635 129.8 91.965 130.93 ;
        RECT 91.635 127.675 91.965 128.005 ;
        RECT 91.635 126.315 91.965 126.645 ;
        RECT 91.635 124.955 91.965 125.285 ;
        RECT 91.635 123.595 91.965 123.925 ;
        RECT 91.64 123.595 91.96 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.635 -1.525 91.965 -1.195 ;
        RECT 91.635 -2.885 91.965 -2.555 ;
        RECT 91.64 -3.56 91.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.995 129.8 93.325 130.93 ;
        RECT 92.995 127.675 93.325 128.005 ;
        RECT 92.995 126.315 93.325 126.645 ;
        RECT 92.995 124.955 93.325 125.285 ;
        RECT 92.995 123.595 93.325 123.925 ;
        RECT 93 123.595 93.32 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.995 -1.525 93.325 -1.195 ;
        RECT 92.995 -2.885 93.325 -2.555 ;
        RECT 93 -3.56 93.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.995 -118.485 93.325 -118.155 ;
        RECT 92.995 -119.845 93.325 -119.515 ;
        RECT 92.995 -121.205 93.325 -120.875 ;
        RECT 92.995 -122.565 93.325 -122.235 ;
        RECT 92.995 -123.925 93.325 -123.595 ;
        RECT 92.995 -125.285 93.325 -124.955 ;
        RECT 92.995 -126.645 93.325 -126.315 ;
        RECT 92.995 -128.005 93.325 -127.675 ;
        RECT 92.995 -129.365 93.325 -129.035 ;
        RECT 92.995 -130.725 93.325 -130.395 ;
        RECT 92.995 -132.085 93.325 -131.755 ;
        RECT 92.995 -133.445 93.325 -133.115 ;
        RECT 92.995 -134.805 93.325 -134.475 ;
        RECT 92.995 -136.165 93.325 -135.835 ;
        RECT 92.995 -137.525 93.325 -137.195 ;
        RECT 92.995 -138.885 93.325 -138.555 ;
        RECT 92.995 -140.245 93.325 -139.915 ;
        RECT 92.995 -141.605 93.325 -141.275 ;
        RECT 92.995 -142.965 93.325 -142.635 ;
        RECT 92.995 -144.325 93.325 -143.995 ;
        RECT 92.995 -145.685 93.325 -145.355 ;
        RECT 92.995 -147.045 93.325 -146.715 ;
        RECT 92.995 -148.405 93.325 -148.075 ;
        RECT 92.995 -149.765 93.325 -149.435 ;
        RECT 92.995 -151.125 93.325 -150.795 ;
        RECT 92.995 -152.485 93.325 -152.155 ;
        RECT 92.995 -153.845 93.325 -153.515 ;
        RECT 92.995 -155.205 93.325 -154.875 ;
        RECT 92.995 -156.565 93.325 -156.235 ;
        RECT 92.995 -157.925 93.325 -157.595 ;
        RECT 92.995 -159.285 93.325 -158.955 ;
        RECT 92.995 -160.645 93.325 -160.315 ;
        RECT 92.995 -162.005 93.325 -161.675 ;
        RECT 92.995 -163.365 93.325 -163.035 ;
        RECT 92.995 -164.725 93.325 -164.395 ;
        RECT 92.995 -166.085 93.325 -165.755 ;
        RECT 92.995 -167.445 93.325 -167.115 ;
        RECT 92.995 -168.805 93.325 -168.475 ;
        RECT 92.995 -170.165 93.325 -169.835 ;
        RECT 92.995 -171.525 93.325 -171.195 ;
        RECT 92.995 -172.885 93.325 -172.555 ;
        RECT 92.995 -174.245 93.325 -173.915 ;
        RECT 92.995 -175.605 93.325 -175.275 ;
        RECT 92.995 -176.965 93.325 -176.635 ;
        RECT 92.995 -178.325 93.325 -177.995 ;
        RECT 92.995 -179.685 93.325 -179.355 ;
        RECT 92.995 -181.045 93.325 -180.715 ;
        RECT 92.995 -182.405 93.325 -182.075 ;
        RECT 92.995 -183.765 93.325 -183.435 ;
        RECT 92.995 -185.125 93.325 -184.795 ;
        RECT 92.995 -186.485 93.325 -186.155 ;
        RECT 92.995 -187.845 93.325 -187.515 ;
        RECT 92.995 -189.205 93.325 -188.875 ;
        RECT 92.995 -190.565 93.325 -190.235 ;
        RECT 92.995 -191.925 93.325 -191.595 ;
        RECT 92.995 -193.285 93.325 -192.955 ;
        RECT 92.995 -194.645 93.325 -194.315 ;
        RECT 92.995 -196.005 93.325 -195.675 ;
        RECT 92.995 -197.365 93.325 -197.035 ;
        RECT 92.995 -198.725 93.325 -198.395 ;
        RECT 92.995 -200.085 93.325 -199.755 ;
        RECT 92.995 -201.445 93.325 -201.115 ;
        RECT 92.995 -202.805 93.325 -202.475 ;
        RECT 92.995 -204.165 93.325 -203.835 ;
        RECT 92.995 -205.525 93.325 -205.195 ;
        RECT 92.995 -206.885 93.325 -206.555 ;
        RECT 92.995 -208.245 93.325 -207.915 ;
        RECT 92.995 -209.605 93.325 -209.275 ;
        RECT 92.995 -210.965 93.325 -210.635 ;
        RECT 92.995 -212.325 93.325 -211.995 ;
        RECT 92.995 -213.685 93.325 -213.355 ;
        RECT 92.995 -215.045 93.325 -214.715 ;
        RECT 92.995 -216.405 93.325 -216.075 ;
        RECT 92.995 -217.765 93.325 -217.435 ;
        RECT 92.995 -219.125 93.325 -218.795 ;
        RECT 92.995 -221.37 93.325 -220.24 ;
        RECT 93 -221.485 93.32 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.355 129.8 94.685 130.93 ;
        RECT 94.355 127.675 94.685 128.005 ;
        RECT 94.355 126.315 94.685 126.645 ;
        RECT 94.355 124.955 94.685 125.285 ;
        RECT 94.355 123.595 94.685 123.925 ;
        RECT 94.36 123.595 94.68 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.355 -122.565 94.685 -122.235 ;
        RECT 94.355 -123.925 94.685 -123.595 ;
        RECT 94.355 -125.285 94.685 -124.955 ;
        RECT 94.355 -126.645 94.685 -126.315 ;
        RECT 94.355 -128.005 94.685 -127.675 ;
        RECT 94.355 -129.365 94.685 -129.035 ;
        RECT 94.355 -130.725 94.685 -130.395 ;
        RECT 94.355 -132.085 94.685 -131.755 ;
        RECT 94.355 -133.445 94.685 -133.115 ;
        RECT 94.355 -134.805 94.685 -134.475 ;
        RECT 94.355 -136.165 94.685 -135.835 ;
        RECT 94.355 -137.525 94.685 -137.195 ;
        RECT 94.355 -138.885 94.685 -138.555 ;
        RECT 94.355 -140.245 94.685 -139.915 ;
        RECT 94.355 -141.605 94.685 -141.275 ;
        RECT 94.355 -142.965 94.685 -142.635 ;
        RECT 94.355 -144.325 94.685 -143.995 ;
        RECT 94.355 -145.685 94.685 -145.355 ;
        RECT 94.355 -147.045 94.685 -146.715 ;
        RECT 94.355 -148.405 94.685 -148.075 ;
        RECT 94.355 -149.765 94.685 -149.435 ;
        RECT 94.355 -151.125 94.685 -150.795 ;
        RECT 94.355 -152.485 94.685 -152.155 ;
        RECT 94.355 -153.845 94.685 -153.515 ;
        RECT 94.355 -155.205 94.685 -154.875 ;
        RECT 94.355 -156.565 94.685 -156.235 ;
        RECT 94.355 -157.925 94.685 -157.595 ;
        RECT 94.355 -159.285 94.685 -158.955 ;
        RECT 94.355 -160.645 94.685 -160.315 ;
        RECT 94.355 -162.005 94.685 -161.675 ;
        RECT 94.355 -163.365 94.685 -163.035 ;
        RECT 94.355 -164.725 94.685 -164.395 ;
        RECT 94.355 -166.085 94.685 -165.755 ;
        RECT 94.355 -167.445 94.685 -167.115 ;
        RECT 94.355 -168.805 94.685 -168.475 ;
        RECT 94.355 -170.165 94.685 -169.835 ;
        RECT 94.355 -171.525 94.685 -171.195 ;
        RECT 94.355 -172.885 94.685 -172.555 ;
        RECT 94.355 -174.245 94.685 -173.915 ;
        RECT 94.355 -175.605 94.685 -175.275 ;
        RECT 94.355 -176.965 94.685 -176.635 ;
        RECT 94.355 -178.325 94.685 -177.995 ;
        RECT 94.355 -179.685 94.685 -179.355 ;
        RECT 94.355 -181.045 94.685 -180.715 ;
        RECT 94.355 -182.405 94.685 -182.075 ;
        RECT 94.355 -183.765 94.685 -183.435 ;
        RECT 94.355 -185.125 94.685 -184.795 ;
        RECT 94.355 -186.485 94.685 -186.155 ;
        RECT 94.355 -187.845 94.685 -187.515 ;
        RECT 94.355 -189.205 94.685 -188.875 ;
        RECT 94.355 -190.565 94.685 -190.235 ;
        RECT 94.355 -191.925 94.685 -191.595 ;
        RECT 94.355 -193.285 94.685 -192.955 ;
        RECT 94.355 -194.645 94.685 -194.315 ;
        RECT 94.355 -196.005 94.685 -195.675 ;
        RECT 94.355 -197.365 94.685 -197.035 ;
        RECT 94.355 -198.725 94.685 -198.395 ;
        RECT 94.355 -200.085 94.685 -199.755 ;
        RECT 94.355 -201.445 94.685 -201.115 ;
        RECT 94.355 -202.805 94.685 -202.475 ;
        RECT 94.355 -204.165 94.685 -203.835 ;
        RECT 94.355 -205.525 94.685 -205.195 ;
        RECT 94.355 -206.885 94.685 -206.555 ;
        RECT 94.355 -208.245 94.685 -207.915 ;
        RECT 94.355 -209.605 94.685 -209.275 ;
        RECT 94.355 -210.965 94.685 -210.635 ;
        RECT 94.355 -212.325 94.685 -211.995 ;
        RECT 94.355 -213.685 94.685 -213.355 ;
        RECT 94.355 -215.045 94.685 -214.715 ;
        RECT 94.355 -216.405 94.685 -216.075 ;
        RECT 94.355 -217.765 94.685 -217.435 ;
        RECT 94.355 -219.125 94.685 -218.795 ;
        RECT 94.355 -221.37 94.685 -220.24 ;
        RECT 94.36 -221.485 94.68 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.81 -121.535 95.14 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.715 129.8 96.045 130.93 ;
        RECT 95.715 127.675 96.045 128.005 ;
        RECT 95.715 126.315 96.045 126.645 ;
        RECT 95.715 124.955 96.045 125.285 ;
        RECT 95.715 123.595 96.045 123.925 ;
        RECT 95.72 123.595 96.04 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.715 -1.525 96.045 -1.195 ;
        RECT 95.715 -2.885 96.045 -2.555 ;
        RECT 95.72 -3.56 96.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.075 129.8 97.405 130.93 ;
        RECT 97.075 127.675 97.405 128.005 ;
        RECT 97.075 126.315 97.405 126.645 ;
        RECT 97.075 124.955 97.405 125.285 ;
        RECT 97.075 123.595 97.405 123.925 ;
        RECT 97.08 123.595 97.4 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.075 -1.525 97.405 -1.195 ;
        RECT 97.075 -2.885 97.405 -2.555 ;
        RECT 97.08 -3.56 97.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.435 129.8 98.765 130.93 ;
        RECT 98.435 127.675 98.765 128.005 ;
        RECT 98.435 126.315 98.765 126.645 ;
        RECT 98.435 124.955 98.765 125.285 ;
        RECT 98.435 123.595 98.765 123.925 ;
        RECT 98.44 123.595 98.76 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.435 -1.525 98.765 -1.195 ;
        RECT 98.435 -2.885 98.765 -2.555 ;
        RECT 98.44 -3.56 98.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.435 -118.485 98.765 -118.155 ;
        RECT 98.435 -119.845 98.765 -119.515 ;
        RECT 98.435 -121.205 98.765 -120.875 ;
        RECT 98.435 -122.565 98.765 -122.235 ;
        RECT 98.435 -123.925 98.765 -123.595 ;
        RECT 98.435 -125.285 98.765 -124.955 ;
        RECT 98.435 -126.645 98.765 -126.315 ;
        RECT 98.435 -128.005 98.765 -127.675 ;
        RECT 98.435 -129.365 98.765 -129.035 ;
        RECT 98.435 -130.725 98.765 -130.395 ;
        RECT 98.435 -132.085 98.765 -131.755 ;
        RECT 98.435 -133.445 98.765 -133.115 ;
        RECT 98.435 -134.805 98.765 -134.475 ;
        RECT 98.435 -136.165 98.765 -135.835 ;
        RECT 98.435 -137.525 98.765 -137.195 ;
        RECT 98.435 -138.885 98.765 -138.555 ;
        RECT 98.435 -140.245 98.765 -139.915 ;
        RECT 98.435 -141.605 98.765 -141.275 ;
        RECT 98.435 -142.965 98.765 -142.635 ;
        RECT 98.435 -144.325 98.765 -143.995 ;
        RECT 98.435 -145.685 98.765 -145.355 ;
        RECT 98.435 -147.045 98.765 -146.715 ;
        RECT 98.435 -148.405 98.765 -148.075 ;
        RECT 98.435 -149.765 98.765 -149.435 ;
        RECT 98.435 -151.125 98.765 -150.795 ;
        RECT 98.435 -152.485 98.765 -152.155 ;
        RECT 98.435 -153.845 98.765 -153.515 ;
        RECT 98.435 -155.205 98.765 -154.875 ;
        RECT 98.435 -156.565 98.765 -156.235 ;
        RECT 98.435 -157.925 98.765 -157.595 ;
        RECT 98.435 -159.285 98.765 -158.955 ;
        RECT 98.435 -160.645 98.765 -160.315 ;
        RECT 98.435 -162.005 98.765 -161.675 ;
        RECT 98.435 -163.365 98.765 -163.035 ;
        RECT 98.435 -164.725 98.765 -164.395 ;
        RECT 98.435 -166.085 98.765 -165.755 ;
        RECT 98.435 -167.445 98.765 -167.115 ;
        RECT 98.435 -168.805 98.765 -168.475 ;
        RECT 98.435 -170.165 98.765 -169.835 ;
        RECT 98.435 -171.525 98.765 -171.195 ;
        RECT 98.435 -172.885 98.765 -172.555 ;
        RECT 98.435 -174.245 98.765 -173.915 ;
        RECT 98.435 -175.605 98.765 -175.275 ;
        RECT 98.435 -176.965 98.765 -176.635 ;
        RECT 98.435 -178.325 98.765 -177.995 ;
        RECT 98.435 -179.685 98.765 -179.355 ;
        RECT 98.435 -181.045 98.765 -180.715 ;
        RECT 98.435 -182.405 98.765 -182.075 ;
        RECT 98.435 -183.765 98.765 -183.435 ;
        RECT 98.435 -185.125 98.765 -184.795 ;
        RECT 98.435 -186.485 98.765 -186.155 ;
        RECT 98.435 -187.845 98.765 -187.515 ;
        RECT 98.435 -189.205 98.765 -188.875 ;
        RECT 98.435 -190.565 98.765 -190.235 ;
        RECT 98.435 -191.925 98.765 -191.595 ;
        RECT 98.435 -193.285 98.765 -192.955 ;
        RECT 98.435 -194.645 98.765 -194.315 ;
        RECT 98.435 -196.005 98.765 -195.675 ;
        RECT 98.435 -197.365 98.765 -197.035 ;
        RECT 98.435 -198.725 98.765 -198.395 ;
        RECT 98.435 -200.085 98.765 -199.755 ;
        RECT 98.435 -201.445 98.765 -201.115 ;
        RECT 98.435 -202.805 98.765 -202.475 ;
        RECT 98.435 -204.165 98.765 -203.835 ;
        RECT 98.435 -205.525 98.765 -205.195 ;
        RECT 98.435 -206.885 98.765 -206.555 ;
        RECT 98.435 -208.245 98.765 -207.915 ;
        RECT 98.435 -209.605 98.765 -209.275 ;
        RECT 98.435 -210.965 98.765 -210.635 ;
        RECT 98.435 -212.325 98.765 -211.995 ;
        RECT 98.435 -213.685 98.765 -213.355 ;
        RECT 98.435 -215.045 98.765 -214.715 ;
        RECT 98.435 -216.405 98.765 -216.075 ;
        RECT 98.435 -217.765 98.765 -217.435 ;
        RECT 98.435 -219.125 98.765 -218.795 ;
        RECT 98.435 -221.37 98.765 -220.24 ;
        RECT 98.44 -221.485 98.76 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.795 129.8 100.125 130.93 ;
        RECT 99.795 127.675 100.125 128.005 ;
        RECT 99.795 126.315 100.125 126.645 ;
        RECT 99.795 124.955 100.125 125.285 ;
        RECT 99.795 123.595 100.125 123.925 ;
        RECT 99.8 123.595 100.12 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.795 -122.565 100.125 -122.235 ;
        RECT 99.795 -123.925 100.125 -123.595 ;
        RECT 99.795 -125.285 100.125 -124.955 ;
        RECT 99.795 -126.645 100.125 -126.315 ;
        RECT 99.795 -128.005 100.125 -127.675 ;
        RECT 99.795 -129.365 100.125 -129.035 ;
        RECT 99.795 -130.725 100.125 -130.395 ;
        RECT 99.795 -132.085 100.125 -131.755 ;
        RECT 99.795 -133.445 100.125 -133.115 ;
        RECT 99.795 -134.805 100.125 -134.475 ;
        RECT 99.795 -136.165 100.125 -135.835 ;
        RECT 99.795 -137.525 100.125 -137.195 ;
        RECT 99.795 -138.885 100.125 -138.555 ;
        RECT 99.795 -140.245 100.125 -139.915 ;
        RECT 99.795 -141.605 100.125 -141.275 ;
        RECT 99.795 -142.965 100.125 -142.635 ;
        RECT 99.795 -144.325 100.125 -143.995 ;
        RECT 99.795 -145.685 100.125 -145.355 ;
        RECT 99.795 -147.045 100.125 -146.715 ;
        RECT 99.795 -148.405 100.125 -148.075 ;
        RECT 99.795 -149.765 100.125 -149.435 ;
        RECT 99.795 -151.125 100.125 -150.795 ;
        RECT 99.795 -152.485 100.125 -152.155 ;
        RECT 99.795 -153.845 100.125 -153.515 ;
        RECT 99.795 -155.205 100.125 -154.875 ;
        RECT 99.795 -156.565 100.125 -156.235 ;
        RECT 99.795 -157.925 100.125 -157.595 ;
        RECT 99.795 -159.285 100.125 -158.955 ;
        RECT 99.795 -160.645 100.125 -160.315 ;
        RECT 99.795 -162.005 100.125 -161.675 ;
        RECT 99.795 -163.365 100.125 -163.035 ;
        RECT 99.795 -164.725 100.125 -164.395 ;
        RECT 99.795 -166.085 100.125 -165.755 ;
        RECT 99.795 -167.445 100.125 -167.115 ;
        RECT 99.795 -168.805 100.125 -168.475 ;
        RECT 99.795 -170.165 100.125 -169.835 ;
        RECT 99.795 -171.525 100.125 -171.195 ;
        RECT 99.795 -172.885 100.125 -172.555 ;
        RECT 99.795 -174.245 100.125 -173.915 ;
        RECT 99.795 -175.605 100.125 -175.275 ;
        RECT 99.795 -176.965 100.125 -176.635 ;
        RECT 99.795 -178.325 100.125 -177.995 ;
        RECT 99.795 -179.685 100.125 -179.355 ;
        RECT 99.795 -181.045 100.125 -180.715 ;
        RECT 99.795 -182.405 100.125 -182.075 ;
        RECT 99.795 -183.765 100.125 -183.435 ;
        RECT 99.795 -185.125 100.125 -184.795 ;
        RECT 99.795 -186.485 100.125 -186.155 ;
        RECT 99.795 -187.845 100.125 -187.515 ;
        RECT 99.795 -189.205 100.125 -188.875 ;
        RECT 99.795 -190.565 100.125 -190.235 ;
        RECT 99.795 -191.925 100.125 -191.595 ;
        RECT 99.795 -193.285 100.125 -192.955 ;
        RECT 99.795 -194.645 100.125 -194.315 ;
        RECT 99.795 -196.005 100.125 -195.675 ;
        RECT 99.795 -197.365 100.125 -197.035 ;
        RECT 99.795 -198.725 100.125 -198.395 ;
        RECT 99.795 -200.085 100.125 -199.755 ;
        RECT 99.795 -201.445 100.125 -201.115 ;
        RECT 99.795 -202.805 100.125 -202.475 ;
        RECT 99.795 -204.165 100.125 -203.835 ;
        RECT 99.795 -205.525 100.125 -205.195 ;
        RECT 99.795 -206.885 100.125 -206.555 ;
        RECT 99.795 -208.245 100.125 -207.915 ;
        RECT 99.795 -209.605 100.125 -209.275 ;
        RECT 99.795 -210.965 100.125 -210.635 ;
        RECT 99.795 -212.325 100.125 -211.995 ;
        RECT 99.795 -213.685 100.125 -213.355 ;
        RECT 99.795 -215.045 100.125 -214.715 ;
        RECT 99.795 -216.405 100.125 -216.075 ;
        RECT 99.795 -217.765 100.125 -217.435 ;
        RECT 99.795 -219.125 100.125 -218.795 ;
        RECT 99.795 -221.37 100.125 -220.24 ;
        RECT 99.8 -221.485 100.12 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.91 -121.535 101.24 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.155 129.8 101.485 130.93 ;
        RECT 101.155 127.675 101.485 128.005 ;
        RECT 101.155 126.315 101.485 126.645 ;
        RECT 101.155 124.955 101.485 125.285 ;
        RECT 101.155 123.595 101.485 123.925 ;
        RECT 101.16 123.595 101.48 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.515 129.8 102.845 130.93 ;
        RECT 102.515 127.675 102.845 128.005 ;
        RECT 102.515 126.315 102.845 126.645 ;
        RECT 102.515 124.955 102.845 125.285 ;
        RECT 102.515 123.595 102.845 123.925 ;
        RECT 102.52 123.595 102.84 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.515 -1.525 102.845 -1.195 ;
        RECT 102.515 -2.885 102.845 -2.555 ;
        RECT 102.52 -3.56 102.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.515 -118.485 102.845 -118.155 ;
        RECT 102.515 -119.845 102.845 -119.515 ;
        RECT 102.515 -121.205 102.845 -120.875 ;
        RECT 102.515 -122.565 102.845 -122.235 ;
        RECT 102.515 -123.925 102.845 -123.595 ;
        RECT 102.515 -125.285 102.845 -124.955 ;
        RECT 102.515 -126.645 102.845 -126.315 ;
        RECT 102.515 -128.005 102.845 -127.675 ;
        RECT 102.515 -129.365 102.845 -129.035 ;
        RECT 102.515 -130.725 102.845 -130.395 ;
        RECT 102.515 -132.085 102.845 -131.755 ;
        RECT 102.515 -133.445 102.845 -133.115 ;
        RECT 102.515 -134.805 102.845 -134.475 ;
        RECT 102.515 -136.165 102.845 -135.835 ;
        RECT 102.515 -137.525 102.845 -137.195 ;
        RECT 102.515 -138.885 102.845 -138.555 ;
        RECT 102.515 -140.245 102.845 -139.915 ;
        RECT 102.515 -141.605 102.845 -141.275 ;
        RECT 102.515 -142.965 102.845 -142.635 ;
        RECT 102.515 -144.325 102.845 -143.995 ;
        RECT 102.515 -145.685 102.845 -145.355 ;
        RECT 102.515 -147.045 102.845 -146.715 ;
        RECT 102.515 -148.405 102.845 -148.075 ;
        RECT 102.515 -149.765 102.845 -149.435 ;
        RECT 102.515 -151.125 102.845 -150.795 ;
        RECT 102.515 -152.485 102.845 -152.155 ;
        RECT 102.515 -153.845 102.845 -153.515 ;
        RECT 102.515 -155.205 102.845 -154.875 ;
        RECT 102.515 -156.565 102.845 -156.235 ;
        RECT 102.515 -157.925 102.845 -157.595 ;
        RECT 102.515 -159.285 102.845 -158.955 ;
        RECT 102.515 -160.645 102.845 -160.315 ;
        RECT 102.515 -162.005 102.845 -161.675 ;
        RECT 102.515 -163.365 102.845 -163.035 ;
        RECT 102.515 -164.725 102.845 -164.395 ;
        RECT 102.515 -166.085 102.845 -165.755 ;
        RECT 102.515 -167.445 102.845 -167.115 ;
        RECT 102.515 -168.805 102.845 -168.475 ;
        RECT 102.515 -170.165 102.845 -169.835 ;
        RECT 102.515 -171.525 102.845 -171.195 ;
        RECT 102.515 -172.885 102.845 -172.555 ;
        RECT 102.515 -174.245 102.845 -173.915 ;
        RECT 102.515 -175.605 102.845 -175.275 ;
        RECT 102.515 -176.965 102.845 -176.635 ;
        RECT 102.515 -178.325 102.845 -177.995 ;
        RECT 102.515 -179.685 102.845 -179.355 ;
        RECT 102.515 -181.045 102.845 -180.715 ;
        RECT 102.515 -182.405 102.845 -182.075 ;
        RECT 102.515 -183.765 102.845 -183.435 ;
        RECT 102.515 -185.125 102.845 -184.795 ;
        RECT 102.515 -186.485 102.845 -186.155 ;
        RECT 102.515 -187.845 102.845 -187.515 ;
        RECT 102.515 -189.205 102.845 -188.875 ;
        RECT 102.515 -190.565 102.845 -190.235 ;
        RECT 102.515 -191.925 102.845 -191.595 ;
        RECT 102.515 -193.285 102.845 -192.955 ;
        RECT 102.515 -194.645 102.845 -194.315 ;
        RECT 102.515 -196.005 102.845 -195.675 ;
        RECT 102.515 -197.365 102.845 -197.035 ;
        RECT 102.515 -198.725 102.845 -198.395 ;
        RECT 102.515 -200.085 102.845 -199.755 ;
        RECT 102.515 -201.445 102.845 -201.115 ;
        RECT 102.515 -202.805 102.845 -202.475 ;
        RECT 102.515 -204.165 102.845 -203.835 ;
        RECT 102.515 -205.525 102.845 -205.195 ;
        RECT 102.515 -206.885 102.845 -206.555 ;
        RECT 102.515 -208.245 102.845 -207.915 ;
        RECT 102.515 -209.605 102.845 -209.275 ;
        RECT 102.515 -210.965 102.845 -210.635 ;
        RECT 102.515 -212.325 102.845 -211.995 ;
        RECT 102.515 -213.685 102.845 -213.355 ;
        RECT 102.515 -215.045 102.845 -214.715 ;
        RECT 102.515 -216.405 102.845 -216.075 ;
        RECT 102.515 -217.765 102.845 -217.435 ;
        RECT 102.515 -219.125 102.845 -218.795 ;
        RECT 102.515 -221.37 102.845 -220.24 ;
        RECT 102.52 -221.485 102.84 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.875 129.8 104.205 130.93 ;
        RECT 103.875 127.675 104.205 128.005 ;
        RECT 103.875 126.315 104.205 126.645 ;
        RECT 103.875 124.955 104.205 125.285 ;
        RECT 103.875 123.595 104.205 123.925 ;
        RECT 103.88 123.595 104.2 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.875 -1.525 104.205 -1.195 ;
        RECT 103.875 -2.885 104.205 -2.555 ;
        RECT 103.88 -3.56 104.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.235 129.8 105.565 130.93 ;
        RECT 105.235 127.675 105.565 128.005 ;
        RECT 105.235 126.315 105.565 126.645 ;
        RECT 105.235 124.955 105.565 125.285 ;
        RECT 105.235 123.595 105.565 123.925 ;
        RECT 105.24 123.595 105.56 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.235 -1.525 105.565 -1.195 ;
        RECT 105.235 -2.885 105.565 -2.555 ;
        RECT 105.24 -3.56 105.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.235 -179.685 105.565 -179.355 ;
        RECT 105.235 -181.045 105.565 -180.715 ;
        RECT 105.235 -182.405 105.565 -182.075 ;
        RECT 105.235 -183.765 105.565 -183.435 ;
        RECT 105.235 -185.125 105.565 -184.795 ;
        RECT 105.235 -186.485 105.565 -186.155 ;
        RECT 105.235 -187.845 105.565 -187.515 ;
        RECT 105.235 -189.205 105.565 -188.875 ;
        RECT 105.235 -190.565 105.565 -190.235 ;
        RECT 105.235 -191.925 105.565 -191.595 ;
        RECT 105.235 -193.285 105.565 -192.955 ;
        RECT 105.235 -194.645 105.565 -194.315 ;
        RECT 105.235 -196.005 105.565 -195.675 ;
        RECT 105.235 -197.365 105.565 -197.035 ;
        RECT 105.235 -198.725 105.565 -198.395 ;
        RECT 105.235 -200.085 105.565 -199.755 ;
        RECT 105.235 -201.445 105.565 -201.115 ;
        RECT 105.235 -202.805 105.565 -202.475 ;
        RECT 105.235 -204.165 105.565 -203.835 ;
        RECT 105.235 -205.525 105.565 -205.195 ;
        RECT 105.235 -206.885 105.565 -206.555 ;
        RECT 105.235 -208.245 105.565 -207.915 ;
        RECT 105.235 -209.605 105.565 -209.275 ;
        RECT 105.235 -210.965 105.565 -210.635 ;
        RECT 105.235 -212.325 105.565 -211.995 ;
        RECT 105.235 -213.685 105.565 -213.355 ;
        RECT 105.235 -215.045 105.565 -214.715 ;
        RECT 105.235 -216.405 105.565 -216.075 ;
        RECT 105.235 -217.765 105.565 -217.435 ;
        RECT 105.235 -219.125 105.565 -218.795 ;
        RECT 105.235 -221.37 105.565 -220.24 ;
        RECT 105.24 -221.485 105.56 -118.155 ;
        RECT 105.235 -118.485 105.565 -118.155 ;
        RECT 105.235 -119.845 105.565 -119.515 ;
        RECT 105.235 -121.205 105.565 -120.875 ;
        RECT 105.235 -122.565 105.565 -122.235 ;
        RECT 105.235 -123.925 105.565 -123.595 ;
        RECT 105.235 -125.285 105.565 -124.955 ;
        RECT 105.235 -126.645 105.565 -126.315 ;
        RECT 105.235 -128.005 105.565 -127.675 ;
        RECT 105.235 -129.365 105.565 -129.035 ;
        RECT 105.235 -130.725 105.565 -130.395 ;
        RECT 105.235 -132.085 105.565 -131.755 ;
        RECT 105.235 -133.445 105.565 -133.115 ;
        RECT 105.235 -134.805 105.565 -134.475 ;
        RECT 105.235 -136.165 105.565 -135.835 ;
        RECT 105.235 -137.525 105.565 -137.195 ;
        RECT 105.235 -138.885 105.565 -138.555 ;
        RECT 105.235 -140.245 105.565 -139.915 ;
        RECT 105.235 -141.605 105.565 -141.275 ;
        RECT 105.235 -142.965 105.565 -142.635 ;
        RECT 105.235 -144.325 105.565 -143.995 ;
        RECT 105.235 -145.685 105.565 -145.355 ;
        RECT 105.235 -147.045 105.565 -146.715 ;
        RECT 105.235 -148.405 105.565 -148.075 ;
        RECT 105.235 -149.765 105.565 -149.435 ;
        RECT 105.235 -151.125 105.565 -150.795 ;
        RECT 105.235 -152.485 105.565 -152.155 ;
        RECT 105.235 -153.845 105.565 -153.515 ;
        RECT 105.235 -155.205 105.565 -154.875 ;
        RECT 105.235 -156.565 105.565 -156.235 ;
        RECT 105.235 -157.925 105.565 -157.595 ;
        RECT 105.235 -159.285 105.565 -158.955 ;
        RECT 105.235 -160.645 105.565 -160.315 ;
        RECT 105.235 -162.005 105.565 -161.675 ;
        RECT 105.235 -163.365 105.565 -163.035 ;
        RECT 105.235 -164.725 105.565 -164.395 ;
        RECT 105.235 -166.085 105.565 -165.755 ;
        RECT 105.235 -167.445 105.565 -167.115 ;
        RECT 105.235 -168.805 105.565 -168.475 ;
        RECT 105.235 -170.165 105.565 -169.835 ;
        RECT 105.235 -171.525 105.565 -171.195 ;
        RECT 105.235 -172.885 105.565 -172.555 ;
        RECT 105.235 -174.245 105.565 -173.915 ;
        RECT 105.235 -175.605 105.565 -175.275 ;
        RECT 105.235 -176.965 105.565 -176.635 ;
        RECT 105.235 -178.325 105.565 -177.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.11 -121.535 52.44 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.195 129.8 52.525 130.93 ;
        RECT 52.195 127.675 52.525 128.005 ;
        RECT 52.195 126.315 52.525 126.645 ;
        RECT 52.195 124.955 52.525 125.285 ;
        RECT 52.195 123.595 52.525 123.925 ;
        RECT 52.2 123.595 52.52 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.555 129.8 53.885 130.93 ;
        RECT 53.555 127.675 53.885 128.005 ;
        RECT 53.555 126.315 53.885 126.645 ;
        RECT 53.555 124.955 53.885 125.285 ;
        RECT 53.555 123.595 53.885 123.925 ;
        RECT 53.56 123.595 53.88 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.555 -1.525 53.885 -1.195 ;
        RECT 53.555 -2.885 53.885 -2.555 ;
        RECT 53.56 -3.56 53.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.555 -118.485 53.885 -118.155 ;
        RECT 53.555 -119.845 53.885 -119.515 ;
        RECT 53.555 -121.205 53.885 -120.875 ;
        RECT 53.555 -122.565 53.885 -122.235 ;
        RECT 53.555 -123.925 53.885 -123.595 ;
        RECT 53.555 -125.285 53.885 -124.955 ;
        RECT 53.555 -126.645 53.885 -126.315 ;
        RECT 53.555 -128.005 53.885 -127.675 ;
        RECT 53.555 -129.365 53.885 -129.035 ;
        RECT 53.555 -130.725 53.885 -130.395 ;
        RECT 53.555 -132.085 53.885 -131.755 ;
        RECT 53.555 -133.445 53.885 -133.115 ;
        RECT 53.555 -134.805 53.885 -134.475 ;
        RECT 53.555 -136.165 53.885 -135.835 ;
        RECT 53.555 -137.525 53.885 -137.195 ;
        RECT 53.555 -138.885 53.885 -138.555 ;
        RECT 53.555 -140.245 53.885 -139.915 ;
        RECT 53.555 -141.605 53.885 -141.275 ;
        RECT 53.555 -142.965 53.885 -142.635 ;
        RECT 53.555 -144.325 53.885 -143.995 ;
        RECT 53.555 -145.685 53.885 -145.355 ;
        RECT 53.555 -147.045 53.885 -146.715 ;
        RECT 53.555 -148.405 53.885 -148.075 ;
        RECT 53.555 -149.765 53.885 -149.435 ;
        RECT 53.555 -151.125 53.885 -150.795 ;
        RECT 53.555 -152.485 53.885 -152.155 ;
        RECT 53.555 -153.845 53.885 -153.515 ;
        RECT 53.555 -155.205 53.885 -154.875 ;
        RECT 53.555 -156.565 53.885 -156.235 ;
        RECT 53.555 -157.925 53.885 -157.595 ;
        RECT 53.555 -159.285 53.885 -158.955 ;
        RECT 53.555 -160.645 53.885 -160.315 ;
        RECT 53.555 -162.005 53.885 -161.675 ;
        RECT 53.555 -163.365 53.885 -163.035 ;
        RECT 53.555 -164.725 53.885 -164.395 ;
        RECT 53.555 -166.085 53.885 -165.755 ;
        RECT 53.555 -167.445 53.885 -167.115 ;
        RECT 53.555 -168.805 53.885 -168.475 ;
        RECT 53.555 -170.165 53.885 -169.835 ;
        RECT 53.555 -171.525 53.885 -171.195 ;
        RECT 53.555 -172.885 53.885 -172.555 ;
        RECT 53.555 -174.245 53.885 -173.915 ;
        RECT 53.555 -175.605 53.885 -175.275 ;
        RECT 53.555 -176.965 53.885 -176.635 ;
        RECT 53.555 -178.325 53.885 -177.995 ;
        RECT 53.555 -179.685 53.885 -179.355 ;
        RECT 53.555 -181.045 53.885 -180.715 ;
        RECT 53.555 -182.405 53.885 -182.075 ;
        RECT 53.555 -183.765 53.885 -183.435 ;
        RECT 53.555 -185.125 53.885 -184.795 ;
        RECT 53.555 -186.485 53.885 -186.155 ;
        RECT 53.555 -187.845 53.885 -187.515 ;
        RECT 53.555 -189.205 53.885 -188.875 ;
        RECT 53.555 -190.565 53.885 -190.235 ;
        RECT 53.555 -191.925 53.885 -191.595 ;
        RECT 53.555 -193.285 53.885 -192.955 ;
        RECT 53.555 -194.645 53.885 -194.315 ;
        RECT 53.555 -196.005 53.885 -195.675 ;
        RECT 53.555 -197.365 53.885 -197.035 ;
        RECT 53.555 -198.725 53.885 -198.395 ;
        RECT 53.555 -200.085 53.885 -199.755 ;
        RECT 53.555 -201.445 53.885 -201.115 ;
        RECT 53.555 -202.805 53.885 -202.475 ;
        RECT 53.555 -204.165 53.885 -203.835 ;
        RECT 53.555 -205.525 53.885 -205.195 ;
        RECT 53.555 -206.885 53.885 -206.555 ;
        RECT 53.555 -208.245 53.885 -207.915 ;
        RECT 53.555 -209.605 53.885 -209.275 ;
        RECT 53.555 -210.965 53.885 -210.635 ;
        RECT 53.555 -212.325 53.885 -211.995 ;
        RECT 53.555 -213.685 53.885 -213.355 ;
        RECT 53.555 -215.045 53.885 -214.715 ;
        RECT 53.555 -216.405 53.885 -216.075 ;
        RECT 53.555 -217.765 53.885 -217.435 ;
        RECT 53.555 -219.125 53.885 -218.795 ;
        RECT 53.555 -221.37 53.885 -220.24 ;
        RECT 53.56 -221.485 53.88 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.915 129.8 55.245 130.93 ;
        RECT 54.915 127.675 55.245 128.005 ;
        RECT 54.915 126.315 55.245 126.645 ;
        RECT 54.915 124.955 55.245 125.285 ;
        RECT 54.915 123.595 55.245 123.925 ;
        RECT 54.92 123.595 55.24 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.915 -1.525 55.245 -1.195 ;
        RECT 54.915 -2.885 55.245 -2.555 ;
        RECT 54.92 -3.56 55.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.275 129.8 56.605 130.93 ;
        RECT 56.275 127.675 56.605 128.005 ;
        RECT 56.275 126.315 56.605 126.645 ;
        RECT 56.275 124.955 56.605 125.285 ;
        RECT 56.275 123.595 56.605 123.925 ;
        RECT 56.28 123.595 56.6 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.275 -1.525 56.605 -1.195 ;
        RECT 56.275 -2.885 56.605 -2.555 ;
        RECT 56.28 -3.56 56.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.275 -118.485 56.605 -118.155 ;
        RECT 56.275 -119.845 56.605 -119.515 ;
        RECT 56.275 -121.205 56.605 -120.875 ;
        RECT 56.275 -122.565 56.605 -122.235 ;
        RECT 56.275 -123.925 56.605 -123.595 ;
        RECT 56.275 -125.285 56.605 -124.955 ;
        RECT 56.275 -126.645 56.605 -126.315 ;
        RECT 56.275 -128.005 56.605 -127.675 ;
        RECT 56.275 -129.365 56.605 -129.035 ;
        RECT 56.275 -130.725 56.605 -130.395 ;
        RECT 56.275 -132.085 56.605 -131.755 ;
        RECT 56.275 -133.445 56.605 -133.115 ;
        RECT 56.275 -134.805 56.605 -134.475 ;
        RECT 56.275 -136.165 56.605 -135.835 ;
        RECT 56.275 -137.525 56.605 -137.195 ;
        RECT 56.275 -138.885 56.605 -138.555 ;
        RECT 56.275 -140.245 56.605 -139.915 ;
        RECT 56.275 -141.605 56.605 -141.275 ;
        RECT 56.275 -142.965 56.605 -142.635 ;
        RECT 56.275 -144.325 56.605 -143.995 ;
        RECT 56.275 -145.685 56.605 -145.355 ;
        RECT 56.275 -147.045 56.605 -146.715 ;
        RECT 56.275 -148.405 56.605 -148.075 ;
        RECT 56.275 -149.765 56.605 -149.435 ;
        RECT 56.275 -151.125 56.605 -150.795 ;
        RECT 56.275 -152.485 56.605 -152.155 ;
        RECT 56.275 -153.845 56.605 -153.515 ;
        RECT 56.275 -155.205 56.605 -154.875 ;
        RECT 56.275 -156.565 56.605 -156.235 ;
        RECT 56.275 -157.925 56.605 -157.595 ;
        RECT 56.275 -159.285 56.605 -158.955 ;
        RECT 56.275 -160.645 56.605 -160.315 ;
        RECT 56.275 -162.005 56.605 -161.675 ;
        RECT 56.275 -163.365 56.605 -163.035 ;
        RECT 56.275 -164.725 56.605 -164.395 ;
        RECT 56.275 -166.085 56.605 -165.755 ;
        RECT 56.275 -167.445 56.605 -167.115 ;
        RECT 56.275 -168.805 56.605 -168.475 ;
        RECT 56.275 -170.165 56.605 -169.835 ;
        RECT 56.275 -171.525 56.605 -171.195 ;
        RECT 56.275 -172.885 56.605 -172.555 ;
        RECT 56.275 -174.245 56.605 -173.915 ;
        RECT 56.275 -175.605 56.605 -175.275 ;
        RECT 56.275 -176.965 56.605 -176.635 ;
        RECT 56.275 -178.325 56.605 -177.995 ;
        RECT 56.275 -179.685 56.605 -179.355 ;
        RECT 56.275 -181.045 56.605 -180.715 ;
        RECT 56.275 -182.405 56.605 -182.075 ;
        RECT 56.275 -183.765 56.605 -183.435 ;
        RECT 56.275 -185.125 56.605 -184.795 ;
        RECT 56.275 -186.485 56.605 -186.155 ;
        RECT 56.275 -187.845 56.605 -187.515 ;
        RECT 56.275 -189.205 56.605 -188.875 ;
        RECT 56.275 -190.565 56.605 -190.235 ;
        RECT 56.275 -191.925 56.605 -191.595 ;
        RECT 56.275 -193.285 56.605 -192.955 ;
        RECT 56.275 -194.645 56.605 -194.315 ;
        RECT 56.275 -196.005 56.605 -195.675 ;
        RECT 56.275 -197.365 56.605 -197.035 ;
        RECT 56.275 -198.725 56.605 -198.395 ;
        RECT 56.275 -200.085 56.605 -199.755 ;
        RECT 56.275 -201.445 56.605 -201.115 ;
        RECT 56.275 -202.805 56.605 -202.475 ;
        RECT 56.275 -204.165 56.605 -203.835 ;
        RECT 56.275 -205.525 56.605 -205.195 ;
        RECT 56.275 -206.885 56.605 -206.555 ;
        RECT 56.275 -208.245 56.605 -207.915 ;
        RECT 56.275 -209.605 56.605 -209.275 ;
        RECT 56.275 -210.965 56.605 -210.635 ;
        RECT 56.275 -212.325 56.605 -211.995 ;
        RECT 56.275 -213.685 56.605 -213.355 ;
        RECT 56.275 -215.045 56.605 -214.715 ;
        RECT 56.275 -216.405 56.605 -216.075 ;
        RECT 56.275 -217.765 56.605 -217.435 ;
        RECT 56.275 -219.125 56.605 -218.795 ;
        RECT 56.275 -221.37 56.605 -220.24 ;
        RECT 56.28 -221.485 56.6 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.635 129.8 57.965 130.93 ;
        RECT 57.635 127.675 57.965 128.005 ;
        RECT 57.635 126.315 57.965 126.645 ;
        RECT 57.635 124.955 57.965 125.285 ;
        RECT 57.635 123.595 57.965 123.925 ;
        RECT 57.64 123.595 57.96 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.635 -122.565 57.965 -122.235 ;
        RECT 57.635 -123.925 57.965 -123.595 ;
        RECT 57.635 -125.285 57.965 -124.955 ;
        RECT 57.635 -126.645 57.965 -126.315 ;
        RECT 57.635 -128.005 57.965 -127.675 ;
        RECT 57.635 -129.365 57.965 -129.035 ;
        RECT 57.635 -130.725 57.965 -130.395 ;
        RECT 57.635 -132.085 57.965 -131.755 ;
        RECT 57.635 -133.445 57.965 -133.115 ;
        RECT 57.635 -134.805 57.965 -134.475 ;
        RECT 57.635 -136.165 57.965 -135.835 ;
        RECT 57.635 -137.525 57.965 -137.195 ;
        RECT 57.635 -138.885 57.965 -138.555 ;
        RECT 57.635 -140.245 57.965 -139.915 ;
        RECT 57.635 -141.605 57.965 -141.275 ;
        RECT 57.635 -142.965 57.965 -142.635 ;
        RECT 57.635 -144.325 57.965 -143.995 ;
        RECT 57.635 -145.685 57.965 -145.355 ;
        RECT 57.635 -147.045 57.965 -146.715 ;
        RECT 57.635 -148.405 57.965 -148.075 ;
        RECT 57.635 -149.765 57.965 -149.435 ;
        RECT 57.635 -151.125 57.965 -150.795 ;
        RECT 57.635 -152.485 57.965 -152.155 ;
        RECT 57.635 -153.845 57.965 -153.515 ;
        RECT 57.635 -155.205 57.965 -154.875 ;
        RECT 57.635 -156.565 57.965 -156.235 ;
        RECT 57.635 -157.925 57.965 -157.595 ;
        RECT 57.635 -159.285 57.965 -158.955 ;
        RECT 57.635 -160.645 57.965 -160.315 ;
        RECT 57.635 -162.005 57.965 -161.675 ;
        RECT 57.635 -163.365 57.965 -163.035 ;
        RECT 57.635 -164.725 57.965 -164.395 ;
        RECT 57.635 -166.085 57.965 -165.755 ;
        RECT 57.635 -167.445 57.965 -167.115 ;
        RECT 57.635 -168.805 57.965 -168.475 ;
        RECT 57.635 -170.165 57.965 -169.835 ;
        RECT 57.635 -171.525 57.965 -171.195 ;
        RECT 57.635 -172.885 57.965 -172.555 ;
        RECT 57.635 -174.245 57.965 -173.915 ;
        RECT 57.635 -175.605 57.965 -175.275 ;
        RECT 57.635 -176.965 57.965 -176.635 ;
        RECT 57.635 -178.325 57.965 -177.995 ;
        RECT 57.635 -179.685 57.965 -179.355 ;
        RECT 57.635 -181.045 57.965 -180.715 ;
        RECT 57.635 -182.405 57.965 -182.075 ;
        RECT 57.635 -183.765 57.965 -183.435 ;
        RECT 57.635 -185.125 57.965 -184.795 ;
        RECT 57.635 -186.485 57.965 -186.155 ;
        RECT 57.635 -187.845 57.965 -187.515 ;
        RECT 57.635 -189.205 57.965 -188.875 ;
        RECT 57.635 -190.565 57.965 -190.235 ;
        RECT 57.635 -191.925 57.965 -191.595 ;
        RECT 57.635 -193.285 57.965 -192.955 ;
        RECT 57.635 -194.645 57.965 -194.315 ;
        RECT 57.635 -196.005 57.965 -195.675 ;
        RECT 57.635 -197.365 57.965 -197.035 ;
        RECT 57.635 -198.725 57.965 -198.395 ;
        RECT 57.635 -200.085 57.965 -199.755 ;
        RECT 57.635 -201.445 57.965 -201.115 ;
        RECT 57.635 -202.805 57.965 -202.475 ;
        RECT 57.635 -204.165 57.965 -203.835 ;
        RECT 57.635 -205.525 57.965 -205.195 ;
        RECT 57.635 -206.885 57.965 -206.555 ;
        RECT 57.635 -208.245 57.965 -207.915 ;
        RECT 57.635 -209.605 57.965 -209.275 ;
        RECT 57.635 -210.965 57.965 -210.635 ;
        RECT 57.635 -212.325 57.965 -211.995 ;
        RECT 57.635 -213.685 57.965 -213.355 ;
        RECT 57.635 -215.045 57.965 -214.715 ;
        RECT 57.635 -216.405 57.965 -216.075 ;
        RECT 57.635 -217.765 57.965 -217.435 ;
        RECT 57.635 -219.125 57.965 -218.795 ;
        RECT 57.635 -221.37 57.965 -220.24 ;
        RECT 57.64 -221.485 57.96 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.21 -121.535 58.54 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.995 129.8 59.325 130.93 ;
        RECT 58.995 127.675 59.325 128.005 ;
        RECT 58.995 126.315 59.325 126.645 ;
        RECT 58.995 124.955 59.325 125.285 ;
        RECT 58.995 123.595 59.325 123.925 ;
        RECT 59 123.595 59.32 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.995 -1.525 59.325 -1.195 ;
        RECT 58.995 -2.885 59.325 -2.555 ;
        RECT 59 -3.56 59.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.355 129.8 60.685 130.93 ;
        RECT 60.355 127.675 60.685 128.005 ;
        RECT 60.355 126.315 60.685 126.645 ;
        RECT 60.355 124.955 60.685 125.285 ;
        RECT 60.355 123.595 60.685 123.925 ;
        RECT 60.36 123.595 60.68 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.355 -1.525 60.685 -1.195 ;
        RECT 60.355 -2.885 60.685 -2.555 ;
        RECT 60.36 -3.56 60.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.715 129.8 62.045 130.93 ;
        RECT 61.715 127.675 62.045 128.005 ;
        RECT 61.715 126.315 62.045 126.645 ;
        RECT 61.715 124.955 62.045 125.285 ;
        RECT 61.715 123.595 62.045 123.925 ;
        RECT 61.72 123.595 62.04 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.715 -1.525 62.045 -1.195 ;
        RECT 61.715 -2.885 62.045 -2.555 ;
        RECT 61.72 -3.56 62.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.715 -118.485 62.045 -118.155 ;
        RECT 61.715 -119.845 62.045 -119.515 ;
        RECT 61.715 -121.205 62.045 -120.875 ;
        RECT 61.715 -122.565 62.045 -122.235 ;
        RECT 61.715 -123.925 62.045 -123.595 ;
        RECT 61.715 -125.285 62.045 -124.955 ;
        RECT 61.715 -126.645 62.045 -126.315 ;
        RECT 61.715 -128.005 62.045 -127.675 ;
        RECT 61.715 -129.365 62.045 -129.035 ;
        RECT 61.715 -130.725 62.045 -130.395 ;
        RECT 61.715 -132.085 62.045 -131.755 ;
        RECT 61.715 -133.445 62.045 -133.115 ;
        RECT 61.715 -134.805 62.045 -134.475 ;
        RECT 61.715 -136.165 62.045 -135.835 ;
        RECT 61.715 -137.525 62.045 -137.195 ;
        RECT 61.715 -138.885 62.045 -138.555 ;
        RECT 61.715 -140.245 62.045 -139.915 ;
        RECT 61.715 -141.605 62.045 -141.275 ;
        RECT 61.715 -142.965 62.045 -142.635 ;
        RECT 61.715 -144.325 62.045 -143.995 ;
        RECT 61.715 -145.685 62.045 -145.355 ;
        RECT 61.715 -147.045 62.045 -146.715 ;
        RECT 61.715 -148.405 62.045 -148.075 ;
        RECT 61.715 -149.765 62.045 -149.435 ;
        RECT 61.715 -151.125 62.045 -150.795 ;
        RECT 61.715 -152.485 62.045 -152.155 ;
        RECT 61.715 -153.845 62.045 -153.515 ;
        RECT 61.715 -155.205 62.045 -154.875 ;
        RECT 61.715 -156.565 62.045 -156.235 ;
        RECT 61.715 -157.925 62.045 -157.595 ;
        RECT 61.715 -159.285 62.045 -158.955 ;
        RECT 61.715 -160.645 62.045 -160.315 ;
        RECT 61.715 -162.005 62.045 -161.675 ;
        RECT 61.715 -163.365 62.045 -163.035 ;
        RECT 61.715 -164.725 62.045 -164.395 ;
        RECT 61.715 -166.085 62.045 -165.755 ;
        RECT 61.715 -167.445 62.045 -167.115 ;
        RECT 61.715 -168.805 62.045 -168.475 ;
        RECT 61.715 -170.165 62.045 -169.835 ;
        RECT 61.715 -171.525 62.045 -171.195 ;
        RECT 61.715 -172.885 62.045 -172.555 ;
        RECT 61.715 -174.245 62.045 -173.915 ;
        RECT 61.715 -175.605 62.045 -175.275 ;
        RECT 61.715 -176.965 62.045 -176.635 ;
        RECT 61.715 -178.325 62.045 -177.995 ;
        RECT 61.715 -179.685 62.045 -179.355 ;
        RECT 61.715 -181.045 62.045 -180.715 ;
        RECT 61.715 -182.405 62.045 -182.075 ;
        RECT 61.715 -183.765 62.045 -183.435 ;
        RECT 61.715 -185.125 62.045 -184.795 ;
        RECT 61.715 -186.485 62.045 -186.155 ;
        RECT 61.715 -187.845 62.045 -187.515 ;
        RECT 61.715 -189.205 62.045 -188.875 ;
        RECT 61.715 -190.565 62.045 -190.235 ;
        RECT 61.715 -191.925 62.045 -191.595 ;
        RECT 61.715 -193.285 62.045 -192.955 ;
        RECT 61.715 -194.645 62.045 -194.315 ;
        RECT 61.715 -196.005 62.045 -195.675 ;
        RECT 61.715 -197.365 62.045 -197.035 ;
        RECT 61.715 -198.725 62.045 -198.395 ;
        RECT 61.715 -200.085 62.045 -199.755 ;
        RECT 61.715 -201.445 62.045 -201.115 ;
        RECT 61.715 -202.805 62.045 -202.475 ;
        RECT 61.715 -204.165 62.045 -203.835 ;
        RECT 61.715 -205.525 62.045 -205.195 ;
        RECT 61.715 -206.885 62.045 -206.555 ;
        RECT 61.715 -208.245 62.045 -207.915 ;
        RECT 61.715 -209.605 62.045 -209.275 ;
        RECT 61.715 -210.965 62.045 -210.635 ;
        RECT 61.715 -212.325 62.045 -211.995 ;
        RECT 61.715 -213.685 62.045 -213.355 ;
        RECT 61.715 -215.045 62.045 -214.715 ;
        RECT 61.715 -216.405 62.045 -216.075 ;
        RECT 61.715 -217.765 62.045 -217.435 ;
        RECT 61.715 -219.125 62.045 -218.795 ;
        RECT 61.715 -221.37 62.045 -220.24 ;
        RECT 61.72 -221.485 62.04 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.075 129.8 63.405 130.93 ;
        RECT 63.075 127.675 63.405 128.005 ;
        RECT 63.075 126.315 63.405 126.645 ;
        RECT 63.075 124.955 63.405 125.285 ;
        RECT 63.075 123.595 63.405 123.925 ;
        RECT 63.08 123.595 63.4 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.075 -122.565 63.405 -122.235 ;
        RECT 63.075 -123.925 63.405 -123.595 ;
        RECT 63.075 -125.285 63.405 -124.955 ;
        RECT 63.075 -126.645 63.405 -126.315 ;
        RECT 63.075 -128.005 63.405 -127.675 ;
        RECT 63.075 -129.365 63.405 -129.035 ;
        RECT 63.075 -130.725 63.405 -130.395 ;
        RECT 63.075 -132.085 63.405 -131.755 ;
        RECT 63.075 -133.445 63.405 -133.115 ;
        RECT 63.075 -134.805 63.405 -134.475 ;
        RECT 63.075 -136.165 63.405 -135.835 ;
        RECT 63.075 -137.525 63.405 -137.195 ;
        RECT 63.075 -138.885 63.405 -138.555 ;
        RECT 63.075 -140.245 63.405 -139.915 ;
        RECT 63.075 -141.605 63.405 -141.275 ;
        RECT 63.075 -142.965 63.405 -142.635 ;
        RECT 63.075 -144.325 63.405 -143.995 ;
        RECT 63.075 -145.685 63.405 -145.355 ;
        RECT 63.075 -147.045 63.405 -146.715 ;
        RECT 63.075 -148.405 63.405 -148.075 ;
        RECT 63.075 -149.765 63.405 -149.435 ;
        RECT 63.075 -151.125 63.405 -150.795 ;
        RECT 63.075 -152.485 63.405 -152.155 ;
        RECT 63.075 -153.845 63.405 -153.515 ;
        RECT 63.075 -155.205 63.405 -154.875 ;
        RECT 63.075 -156.565 63.405 -156.235 ;
        RECT 63.075 -157.925 63.405 -157.595 ;
        RECT 63.075 -159.285 63.405 -158.955 ;
        RECT 63.075 -160.645 63.405 -160.315 ;
        RECT 63.075 -162.005 63.405 -161.675 ;
        RECT 63.075 -163.365 63.405 -163.035 ;
        RECT 63.075 -164.725 63.405 -164.395 ;
        RECT 63.075 -166.085 63.405 -165.755 ;
        RECT 63.075 -167.445 63.405 -167.115 ;
        RECT 63.075 -168.805 63.405 -168.475 ;
        RECT 63.075 -170.165 63.405 -169.835 ;
        RECT 63.075 -171.525 63.405 -171.195 ;
        RECT 63.075 -172.885 63.405 -172.555 ;
        RECT 63.075 -174.245 63.405 -173.915 ;
        RECT 63.075 -175.605 63.405 -175.275 ;
        RECT 63.075 -176.965 63.405 -176.635 ;
        RECT 63.075 -178.325 63.405 -177.995 ;
        RECT 63.075 -179.685 63.405 -179.355 ;
        RECT 63.075 -181.045 63.405 -180.715 ;
        RECT 63.075 -182.405 63.405 -182.075 ;
        RECT 63.075 -183.765 63.405 -183.435 ;
        RECT 63.075 -185.125 63.405 -184.795 ;
        RECT 63.075 -186.485 63.405 -186.155 ;
        RECT 63.075 -187.845 63.405 -187.515 ;
        RECT 63.075 -189.205 63.405 -188.875 ;
        RECT 63.075 -190.565 63.405 -190.235 ;
        RECT 63.075 -191.925 63.405 -191.595 ;
        RECT 63.075 -193.285 63.405 -192.955 ;
        RECT 63.075 -194.645 63.405 -194.315 ;
        RECT 63.075 -196.005 63.405 -195.675 ;
        RECT 63.075 -197.365 63.405 -197.035 ;
        RECT 63.075 -198.725 63.405 -198.395 ;
        RECT 63.075 -200.085 63.405 -199.755 ;
        RECT 63.075 -201.445 63.405 -201.115 ;
        RECT 63.075 -202.805 63.405 -202.475 ;
        RECT 63.075 -204.165 63.405 -203.835 ;
        RECT 63.075 -205.525 63.405 -205.195 ;
        RECT 63.075 -206.885 63.405 -206.555 ;
        RECT 63.075 -208.245 63.405 -207.915 ;
        RECT 63.075 -209.605 63.405 -209.275 ;
        RECT 63.075 -210.965 63.405 -210.635 ;
        RECT 63.075 -212.325 63.405 -211.995 ;
        RECT 63.075 -213.685 63.405 -213.355 ;
        RECT 63.075 -215.045 63.405 -214.715 ;
        RECT 63.075 -216.405 63.405 -216.075 ;
        RECT 63.075 -217.765 63.405 -217.435 ;
        RECT 63.075 -219.125 63.405 -218.795 ;
        RECT 63.075 -221.37 63.405 -220.24 ;
        RECT 63.08 -221.485 63.4 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.31 -121.535 64.64 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.435 129.8 64.765 130.93 ;
        RECT 64.435 127.675 64.765 128.005 ;
        RECT 64.435 126.315 64.765 126.645 ;
        RECT 64.435 124.955 64.765 125.285 ;
        RECT 64.435 123.595 64.765 123.925 ;
        RECT 64.44 123.595 64.76 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.795 129.8 66.125 130.93 ;
        RECT 65.795 127.675 66.125 128.005 ;
        RECT 65.795 126.315 66.125 126.645 ;
        RECT 65.795 124.955 66.125 125.285 ;
        RECT 65.795 123.595 66.125 123.925 ;
        RECT 65.8 123.595 66.12 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.795 -1.525 66.125 -1.195 ;
        RECT 65.795 -2.885 66.125 -2.555 ;
        RECT 65.8 -3.56 66.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.795 -118.485 66.125 -118.155 ;
        RECT 65.795 -119.845 66.125 -119.515 ;
        RECT 65.795 -121.205 66.125 -120.875 ;
        RECT 65.795 -122.565 66.125 -122.235 ;
        RECT 65.795 -123.925 66.125 -123.595 ;
        RECT 65.795 -125.285 66.125 -124.955 ;
        RECT 65.795 -126.645 66.125 -126.315 ;
        RECT 65.795 -128.005 66.125 -127.675 ;
        RECT 65.795 -129.365 66.125 -129.035 ;
        RECT 65.795 -130.725 66.125 -130.395 ;
        RECT 65.795 -132.085 66.125 -131.755 ;
        RECT 65.795 -133.445 66.125 -133.115 ;
        RECT 65.795 -134.805 66.125 -134.475 ;
        RECT 65.795 -136.165 66.125 -135.835 ;
        RECT 65.795 -137.525 66.125 -137.195 ;
        RECT 65.795 -138.885 66.125 -138.555 ;
        RECT 65.795 -140.245 66.125 -139.915 ;
        RECT 65.795 -141.605 66.125 -141.275 ;
        RECT 65.795 -142.965 66.125 -142.635 ;
        RECT 65.795 -144.325 66.125 -143.995 ;
        RECT 65.795 -145.685 66.125 -145.355 ;
        RECT 65.795 -147.045 66.125 -146.715 ;
        RECT 65.795 -148.405 66.125 -148.075 ;
        RECT 65.795 -149.765 66.125 -149.435 ;
        RECT 65.795 -151.125 66.125 -150.795 ;
        RECT 65.795 -152.485 66.125 -152.155 ;
        RECT 65.795 -153.845 66.125 -153.515 ;
        RECT 65.795 -155.205 66.125 -154.875 ;
        RECT 65.795 -156.565 66.125 -156.235 ;
        RECT 65.795 -157.925 66.125 -157.595 ;
        RECT 65.795 -159.285 66.125 -158.955 ;
        RECT 65.795 -160.645 66.125 -160.315 ;
        RECT 65.795 -162.005 66.125 -161.675 ;
        RECT 65.795 -163.365 66.125 -163.035 ;
        RECT 65.795 -164.725 66.125 -164.395 ;
        RECT 65.795 -166.085 66.125 -165.755 ;
        RECT 65.795 -167.445 66.125 -167.115 ;
        RECT 65.795 -168.805 66.125 -168.475 ;
        RECT 65.795 -170.165 66.125 -169.835 ;
        RECT 65.795 -171.525 66.125 -171.195 ;
        RECT 65.795 -172.885 66.125 -172.555 ;
        RECT 65.795 -174.245 66.125 -173.915 ;
        RECT 65.795 -175.605 66.125 -175.275 ;
        RECT 65.795 -176.965 66.125 -176.635 ;
        RECT 65.795 -178.325 66.125 -177.995 ;
        RECT 65.795 -179.685 66.125 -179.355 ;
        RECT 65.795 -181.045 66.125 -180.715 ;
        RECT 65.795 -182.405 66.125 -182.075 ;
        RECT 65.795 -183.765 66.125 -183.435 ;
        RECT 65.795 -185.125 66.125 -184.795 ;
        RECT 65.795 -186.485 66.125 -186.155 ;
        RECT 65.795 -187.845 66.125 -187.515 ;
        RECT 65.795 -189.205 66.125 -188.875 ;
        RECT 65.795 -190.565 66.125 -190.235 ;
        RECT 65.795 -191.925 66.125 -191.595 ;
        RECT 65.795 -193.285 66.125 -192.955 ;
        RECT 65.795 -194.645 66.125 -194.315 ;
        RECT 65.795 -196.005 66.125 -195.675 ;
        RECT 65.795 -197.365 66.125 -197.035 ;
        RECT 65.795 -198.725 66.125 -198.395 ;
        RECT 65.795 -200.085 66.125 -199.755 ;
        RECT 65.795 -201.445 66.125 -201.115 ;
        RECT 65.795 -202.805 66.125 -202.475 ;
        RECT 65.795 -204.165 66.125 -203.835 ;
        RECT 65.795 -205.525 66.125 -205.195 ;
        RECT 65.795 -206.885 66.125 -206.555 ;
        RECT 65.795 -208.245 66.125 -207.915 ;
        RECT 65.795 -209.605 66.125 -209.275 ;
        RECT 65.795 -210.965 66.125 -210.635 ;
        RECT 65.795 -212.325 66.125 -211.995 ;
        RECT 65.795 -213.685 66.125 -213.355 ;
        RECT 65.795 -215.045 66.125 -214.715 ;
        RECT 65.795 -216.405 66.125 -216.075 ;
        RECT 65.795 -217.765 66.125 -217.435 ;
        RECT 65.795 -219.125 66.125 -218.795 ;
        RECT 65.795 -221.37 66.125 -220.24 ;
        RECT 65.8 -221.485 66.12 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.155 129.8 67.485 130.93 ;
        RECT 67.155 127.675 67.485 128.005 ;
        RECT 67.155 126.315 67.485 126.645 ;
        RECT 67.155 124.955 67.485 125.285 ;
        RECT 67.155 123.595 67.485 123.925 ;
        RECT 67.16 123.595 67.48 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.155 -1.525 67.485 -1.195 ;
        RECT 67.155 -2.885 67.485 -2.555 ;
        RECT 67.16 -3.56 67.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.515 129.8 68.845 130.93 ;
        RECT 68.515 127.675 68.845 128.005 ;
        RECT 68.515 126.315 68.845 126.645 ;
        RECT 68.515 124.955 68.845 125.285 ;
        RECT 68.515 123.595 68.845 123.925 ;
        RECT 68.52 123.595 68.84 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.515 -1.525 68.845 -1.195 ;
        RECT 68.515 -2.885 68.845 -2.555 ;
        RECT 68.52 -3.56 68.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.515 -118.485 68.845 -118.155 ;
        RECT 68.515 -119.845 68.845 -119.515 ;
        RECT 68.515 -121.205 68.845 -120.875 ;
        RECT 68.515 -122.565 68.845 -122.235 ;
        RECT 68.515 -123.925 68.845 -123.595 ;
        RECT 68.515 -125.285 68.845 -124.955 ;
        RECT 68.515 -126.645 68.845 -126.315 ;
        RECT 68.515 -128.005 68.845 -127.675 ;
        RECT 68.515 -129.365 68.845 -129.035 ;
        RECT 68.515 -130.725 68.845 -130.395 ;
        RECT 68.515 -132.085 68.845 -131.755 ;
        RECT 68.515 -133.445 68.845 -133.115 ;
        RECT 68.515 -134.805 68.845 -134.475 ;
        RECT 68.515 -136.165 68.845 -135.835 ;
        RECT 68.515 -137.525 68.845 -137.195 ;
        RECT 68.515 -138.885 68.845 -138.555 ;
        RECT 68.515 -140.245 68.845 -139.915 ;
        RECT 68.515 -141.605 68.845 -141.275 ;
        RECT 68.515 -142.965 68.845 -142.635 ;
        RECT 68.515 -144.325 68.845 -143.995 ;
        RECT 68.515 -145.685 68.845 -145.355 ;
        RECT 68.515 -147.045 68.845 -146.715 ;
        RECT 68.515 -148.405 68.845 -148.075 ;
        RECT 68.515 -149.765 68.845 -149.435 ;
        RECT 68.515 -151.125 68.845 -150.795 ;
        RECT 68.515 -152.485 68.845 -152.155 ;
        RECT 68.515 -153.845 68.845 -153.515 ;
        RECT 68.515 -155.205 68.845 -154.875 ;
        RECT 68.515 -156.565 68.845 -156.235 ;
        RECT 68.515 -157.925 68.845 -157.595 ;
        RECT 68.515 -159.285 68.845 -158.955 ;
        RECT 68.515 -160.645 68.845 -160.315 ;
        RECT 68.515 -162.005 68.845 -161.675 ;
        RECT 68.515 -163.365 68.845 -163.035 ;
        RECT 68.515 -164.725 68.845 -164.395 ;
        RECT 68.515 -166.085 68.845 -165.755 ;
        RECT 68.515 -167.445 68.845 -167.115 ;
        RECT 68.515 -168.805 68.845 -168.475 ;
        RECT 68.515 -170.165 68.845 -169.835 ;
        RECT 68.515 -171.525 68.845 -171.195 ;
        RECT 68.515 -172.885 68.845 -172.555 ;
        RECT 68.515 -174.245 68.845 -173.915 ;
        RECT 68.515 -175.605 68.845 -175.275 ;
        RECT 68.515 -176.965 68.845 -176.635 ;
        RECT 68.515 -178.325 68.845 -177.995 ;
        RECT 68.515 -179.685 68.845 -179.355 ;
        RECT 68.515 -181.045 68.845 -180.715 ;
        RECT 68.515 -182.405 68.845 -182.075 ;
        RECT 68.515 -183.765 68.845 -183.435 ;
        RECT 68.515 -185.125 68.845 -184.795 ;
        RECT 68.515 -186.485 68.845 -186.155 ;
        RECT 68.515 -187.845 68.845 -187.515 ;
        RECT 68.515 -189.205 68.845 -188.875 ;
        RECT 68.515 -190.565 68.845 -190.235 ;
        RECT 68.515 -191.925 68.845 -191.595 ;
        RECT 68.515 -193.285 68.845 -192.955 ;
        RECT 68.515 -194.645 68.845 -194.315 ;
        RECT 68.515 -196.005 68.845 -195.675 ;
        RECT 68.515 -197.365 68.845 -197.035 ;
        RECT 68.515 -198.725 68.845 -198.395 ;
        RECT 68.515 -200.085 68.845 -199.755 ;
        RECT 68.515 -201.445 68.845 -201.115 ;
        RECT 68.515 -202.805 68.845 -202.475 ;
        RECT 68.515 -204.165 68.845 -203.835 ;
        RECT 68.515 -205.525 68.845 -205.195 ;
        RECT 68.515 -206.885 68.845 -206.555 ;
        RECT 68.515 -208.245 68.845 -207.915 ;
        RECT 68.515 -209.605 68.845 -209.275 ;
        RECT 68.515 -210.965 68.845 -210.635 ;
        RECT 68.515 -212.325 68.845 -211.995 ;
        RECT 68.515 -213.685 68.845 -213.355 ;
        RECT 68.515 -215.045 68.845 -214.715 ;
        RECT 68.515 -216.405 68.845 -216.075 ;
        RECT 68.515 -217.765 68.845 -217.435 ;
        RECT 68.515 -219.125 68.845 -218.795 ;
        RECT 68.515 -221.37 68.845 -220.24 ;
        RECT 68.52 -221.485 68.84 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.875 129.8 70.205 130.93 ;
        RECT 69.875 127.675 70.205 128.005 ;
        RECT 69.875 126.315 70.205 126.645 ;
        RECT 69.875 124.955 70.205 125.285 ;
        RECT 69.875 123.595 70.205 123.925 ;
        RECT 69.88 123.595 70.2 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.875 -122.565 70.205 -122.235 ;
        RECT 69.875 -123.925 70.205 -123.595 ;
        RECT 69.875 -125.285 70.205 -124.955 ;
        RECT 69.875 -126.645 70.205 -126.315 ;
        RECT 69.875 -128.005 70.205 -127.675 ;
        RECT 69.875 -129.365 70.205 -129.035 ;
        RECT 69.875 -130.725 70.205 -130.395 ;
        RECT 69.875 -132.085 70.205 -131.755 ;
        RECT 69.875 -133.445 70.205 -133.115 ;
        RECT 69.875 -134.805 70.205 -134.475 ;
        RECT 69.875 -136.165 70.205 -135.835 ;
        RECT 69.875 -137.525 70.205 -137.195 ;
        RECT 69.875 -138.885 70.205 -138.555 ;
        RECT 69.875 -140.245 70.205 -139.915 ;
        RECT 69.875 -141.605 70.205 -141.275 ;
        RECT 69.875 -142.965 70.205 -142.635 ;
        RECT 69.875 -144.325 70.205 -143.995 ;
        RECT 69.875 -145.685 70.205 -145.355 ;
        RECT 69.875 -147.045 70.205 -146.715 ;
        RECT 69.875 -148.405 70.205 -148.075 ;
        RECT 69.875 -149.765 70.205 -149.435 ;
        RECT 69.875 -151.125 70.205 -150.795 ;
        RECT 69.875 -152.485 70.205 -152.155 ;
        RECT 69.875 -153.845 70.205 -153.515 ;
        RECT 69.875 -155.205 70.205 -154.875 ;
        RECT 69.875 -156.565 70.205 -156.235 ;
        RECT 69.875 -157.925 70.205 -157.595 ;
        RECT 69.875 -159.285 70.205 -158.955 ;
        RECT 69.875 -160.645 70.205 -160.315 ;
        RECT 69.875 -162.005 70.205 -161.675 ;
        RECT 69.875 -163.365 70.205 -163.035 ;
        RECT 69.875 -164.725 70.205 -164.395 ;
        RECT 69.875 -166.085 70.205 -165.755 ;
        RECT 69.875 -167.445 70.205 -167.115 ;
        RECT 69.875 -168.805 70.205 -168.475 ;
        RECT 69.875 -170.165 70.205 -169.835 ;
        RECT 69.875 -171.525 70.205 -171.195 ;
        RECT 69.875 -172.885 70.205 -172.555 ;
        RECT 69.875 -174.245 70.205 -173.915 ;
        RECT 69.875 -175.605 70.205 -175.275 ;
        RECT 69.875 -176.965 70.205 -176.635 ;
        RECT 69.875 -178.325 70.205 -177.995 ;
        RECT 69.875 -179.685 70.205 -179.355 ;
        RECT 69.875 -181.045 70.205 -180.715 ;
        RECT 69.875 -182.405 70.205 -182.075 ;
        RECT 69.875 -183.765 70.205 -183.435 ;
        RECT 69.875 -185.125 70.205 -184.795 ;
        RECT 69.875 -186.485 70.205 -186.155 ;
        RECT 69.875 -187.845 70.205 -187.515 ;
        RECT 69.875 -189.205 70.205 -188.875 ;
        RECT 69.875 -190.565 70.205 -190.235 ;
        RECT 69.875 -191.925 70.205 -191.595 ;
        RECT 69.875 -193.285 70.205 -192.955 ;
        RECT 69.875 -194.645 70.205 -194.315 ;
        RECT 69.875 -196.005 70.205 -195.675 ;
        RECT 69.875 -197.365 70.205 -197.035 ;
        RECT 69.875 -198.725 70.205 -198.395 ;
        RECT 69.875 -200.085 70.205 -199.755 ;
        RECT 69.875 -201.445 70.205 -201.115 ;
        RECT 69.875 -202.805 70.205 -202.475 ;
        RECT 69.875 -204.165 70.205 -203.835 ;
        RECT 69.875 -205.525 70.205 -205.195 ;
        RECT 69.875 -206.885 70.205 -206.555 ;
        RECT 69.875 -208.245 70.205 -207.915 ;
        RECT 69.875 -209.605 70.205 -209.275 ;
        RECT 69.875 -210.965 70.205 -210.635 ;
        RECT 69.875 -212.325 70.205 -211.995 ;
        RECT 69.875 -213.685 70.205 -213.355 ;
        RECT 69.875 -215.045 70.205 -214.715 ;
        RECT 69.875 -216.405 70.205 -216.075 ;
        RECT 69.875 -217.765 70.205 -217.435 ;
        RECT 69.875 -219.125 70.205 -218.795 ;
        RECT 69.875 -221.37 70.205 -220.24 ;
        RECT 69.88 -221.485 70.2 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.41 -121.535 70.74 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.235 129.8 71.565 130.93 ;
        RECT 71.235 127.675 71.565 128.005 ;
        RECT 71.235 126.315 71.565 126.645 ;
        RECT 71.235 124.955 71.565 125.285 ;
        RECT 71.235 123.595 71.565 123.925 ;
        RECT 71.24 123.595 71.56 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.235 -1.525 71.565 -1.195 ;
        RECT 71.235 -2.885 71.565 -2.555 ;
        RECT 71.24 -3.56 71.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.595 129.8 72.925 130.93 ;
        RECT 72.595 127.675 72.925 128.005 ;
        RECT 72.595 126.315 72.925 126.645 ;
        RECT 72.595 124.955 72.925 125.285 ;
        RECT 72.595 123.595 72.925 123.925 ;
        RECT 72.6 123.595 72.92 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.595 -1.525 72.925 -1.195 ;
        RECT 72.595 -2.885 72.925 -2.555 ;
        RECT 72.6 -3.56 72.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 129.8 74.285 130.93 ;
        RECT 73.955 127.675 74.285 128.005 ;
        RECT 73.955 126.315 74.285 126.645 ;
        RECT 73.955 124.955 74.285 125.285 ;
        RECT 73.955 123.595 74.285 123.925 ;
        RECT 73.96 123.595 74.28 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 -1.525 74.285 -1.195 ;
        RECT 73.955 -2.885 74.285 -2.555 ;
        RECT 73.96 -3.56 74.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 -118.485 74.285 -118.155 ;
        RECT 73.955 -119.845 74.285 -119.515 ;
        RECT 73.955 -121.205 74.285 -120.875 ;
        RECT 73.955 -122.565 74.285 -122.235 ;
        RECT 73.955 -123.925 74.285 -123.595 ;
        RECT 73.955 -125.285 74.285 -124.955 ;
        RECT 73.955 -126.645 74.285 -126.315 ;
        RECT 73.955 -128.005 74.285 -127.675 ;
        RECT 73.955 -129.365 74.285 -129.035 ;
        RECT 73.955 -130.725 74.285 -130.395 ;
        RECT 73.955 -132.085 74.285 -131.755 ;
        RECT 73.955 -133.445 74.285 -133.115 ;
        RECT 73.955 -134.805 74.285 -134.475 ;
        RECT 73.955 -136.165 74.285 -135.835 ;
        RECT 73.955 -137.525 74.285 -137.195 ;
        RECT 73.955 -138.885 74.285 -138.555 ;
        RECT 73.955 -140.245 74.285 -139.915 ;
        RECT 73.955 -141.605 74.285 -141.275 ;
        RECT 73.955 -142.965 74.285 -142.635 ;
        RECT 73.955 -144.325 74.285 -143.995 ;
        RECT 73.955 -145.685 74.285 -145.355 ;
        RECT 73.955 -147.045 74.285 -146.715 ;
        RECT 73.955 -148.405 74.285 -148.075 ;
        RECT 73.955 -149.765 74.285 -149.435 ;
        RECT 73.955 -151.125 74.285 -150.795 ;
        RECT 73.955 -152.485 74.285 -152.155 ;
        RECT 73.955 -153.845 74.285 -153.515 ;
        RECT 73.955 -155.205 74.285 -154.875 ;
        RECT 73.955 -156.565 74.285 -156.235 ;
        RECT 73.955 -157.925 74.285 -157.595 ;
        RECT 73.955 -159.285 74.285 -158.955 ;
        RECT 73.955 -160.645 74.285 -160.315 ;
        RECT 73.955 -162.005 74.285 -161.675 ;
        RECT 73.955 -163.365 74.285 -163.035 ;
        RECT 73.955 -164.725 74.285 -164.395 ;
        RECT 73.955 -166.085 74.285 -165.755 ;
        RECT 73.955 -167.445 74.285 -167.115 ;
        RECT 73.955 -168.805 74.285 -168.475 ;
        RECT 73.955 -170.165 74.285 -169.835 ;
        RECT 73.955 -171.525 74.285 -171.195 ;
        RECT 73.955 -172.885 74.285 -172.555 ;
        RECT 73.955 -174.245 74.285 -173.915 ;
        RECT 73.955 -175.605 74.285 -175.275 ;
        RECT 73.955 -176.965 74.285 -176.635 ;
        RECT 73.955 -178.325 74.285 -177.995 ;
        RECT 73.955 -179.685 74.285 -179.355 ;
        RECT 73.955 -181.045 74.285 -180.715 ;
        RECT 73.955 -182.405 74.285 -182.075 ;
        RECT 73.955 -183.765 74.285 -183.435 ;
        RECT 73.955 -185.125 74.285 -184.795 ;
        RECT 73.955 -186.485 74.285 -186.155 ;
        RECT 73.955 -187.845 74.285 -187.515 ;
        RECT 73.955 -189.205 74.285 -188.875 ;
        RECT 73.955 -190.565 74.285 -190.235 ;
        RECT 73.955 -191.925 74.285 -191.595 ;
        RECT 73.955 -193.285 74.285 -192.955 ;
        RECT 73.955 -194.645 74.285 -194.315 ;
        RECT 73.955 -196.005 74.285 -195.675 ;
        RECT 73.955 -197.365 74.285 -197.035 ;
        RECT 73.955 -198.725 74.285 -198.395 ;
        RECT 73.955 -200.085 74.285 -199.755 ;
        RECT 73.955 -201.445 74.285 -201.115 ;
        RECT 73.955 -202.805 74.285 -202.475 ;
        RECT 73.955 -204.165 74.285 -203.835 ;
        RECT 73.955 -205.525 74.285 -205.195 ;
        RECT 73.955 -206.885 74.285 -206.555 ;
        RECT 73.955 -208.245 74.285 -207.915 ;
        RECT 73.955 -209.605 74.285 -209.275 ;
        RECT 73.955 -210.965 74.285 -210.635 ;
        RECT 73.955 -212.325 74.285 -211.995 ;
        RECT 73.955 -213.685 74.285 -213.355 ;
        RECT 73.955 -215.045 74.285 -214.715 ;
        RECT 73.955 -216.405 74.285 -216.075 ;
        RECT 73.955 -217.765 74.285 -217.435 ;
        RECT 73.955 -219.125 74.285 -218.795 ;
        RECT 73.955 -221.37 74.285 -220.24 ;
        RECT 73.96 -221.485 74.28 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.315 129.8 75.645 130.93 ;
        RECT 75.315 127.675 75.645 128.005 ;
        RECT 75.315 126.315 75.645 126.645 ;
        RECT 75.315 124.955 75.645 125.285 ;
        RECT 75.315 123.595 75.645 123.925 ;
        RECT 75.32 123.595 75.64 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.315 -122.565 75.645 -122.235 ;
        RECT 75.315 -123.925 75.645 -123.595 ;
        RECT 75.315 -125.285 75.645 -124.955 ;
        RECT 75.315 -126.645 75.645 -126.315 ;
        RECT 75.315 -128.005 75.645 -127.675 ;
        RECT 75.315 -129.365 75.645 -129.035 ;
        RECT 75.315 -130.725 75.645 -130.395 ;
        RECT 75.315 -132.085 75.645 -131.755 ;
        RECT 75.315 -133.445 75.645 -133.115 ;
        RECT 75.315 -134.805 75.645 -134.475 ;
        RECT 75.315 -136.165 75.645 -135.835 ;
        RECT 75.315 -137.525 75.645 -137.195 ;
        RECT 75.315 -138.885 75.645 -138.555 ;
        RECT 75.315 -140.245 75.645 -139.915 ;
        RECT 75.315 -141.605 75.645 -141.275 ;
        RECT 75.315 -142.965 75.645 -142.635 ;
        RECT 75.315 -144.325 75.645 -143.995 ;
        RECT 75.315 -145.685 75.645 -145.355 ;
        RECT 75.315 -147.045 75.645 -146.715 ;
        RECT 75.315 -148.405 75.645 -148.075 ;
        RECT 75.315 -149.765 75.645 -149.435 ;
        RECT 75.315 -151.125 75.645 -150.795 ;
        RECT 75.315 -152.485 75.645 -152.155 ;
        RECT 75.315 -153.845 75.645 -153.515 ;
        RECT 75.315 -155.205 75.645 -154.875 ;
        RECT 75.315 -156.565 75.645 -156.235 ;
        RECT 75.315 -157.925 75.645 -157.595 ;
        RECT 75.315 -159.285 75.645 -158.955 ;
        RECT 75.315 -160.645 75.645 -160.315 ;
        RECT 75.315 -162.005 75.645 -161.675 ;
        RECT 75.315 -163.365 75.645 -163.035 ;
        RECT 75.315 -164.725 75.645 -164.395 ;
        RECT 75.315 -166.085 75.645 -165.755 ;
        RECT 75.315 -167.445 75.645 -167.115 ;
        RECT 75.315 -168.805 75.645 -168.475 ;
        RECT 75.315 -170.165 75.645 -169.835 ;
        RECT 75.315 -171.525 75.645 -171.195 ;
        RECT 75.315 -172.885 75.645 -172.555 ;
        RECT 75.315 -174.245 75.645 -173.915 ;
        RECT 75.315 -175.605 75.645 -175.275 ;
        RECT 75.315 -176.965 75.645 -176.635 ;
        RECT 75.315 -178.325 75.645 -177.995 ;
        RECT 75.315 -179.685 75.645 -179.355 ;
        RECT 75.315 -181.045 75.645 -180.715 ;
        RECT 75.315 -182.405 75.645 -182.075 ;
        RECT 75.315 -183.765 75.645 -183.435 ;
        RECT 75.315 -185.125 75.645 -184.795 ;
        RECT 75.315 -186.485 75.645 -186.155 ;
        RECT 75.315 -187.845 75.645 -187.515 ;
        RECT 75.315 -189.205 75.645 -188.875 ;
        RECT 75.315 -190.565 75.645 -190.235 ;
        RECT 75.315 -191.925 75.645 -191.595 ;
        RECT 75.315 -193.285 75.645 -192.955 ;
        RECT 75.315 -194.645 75.645 -194.315 ;
        RECT 75.315 -196.005 75.645 -195.675 ;
        RECT 75.315 -197.365 75.645 -197.035 ;
        RECT 75.315 -198.725 75.645 -198.395 ;
        RECT 75.315 -200.085 75.645 -199.755 ;
        RECT 75.315 -201.445 75.645 -201.115 ;
        RECT 75.315 -202.805 75.645 -202.475 ;
        RECT 75.315 -204.165 75.645 -203.835 ;
        RECT 75.315 -205.525 75.645 -205.195 ;
        RECT 75.315 -206.885 75.645 -206.555 ;
        RECT 75.315 -208.245 75.645 -207.915 ;
        RECT 75.315 -209.605 75.645 -209.275 ;
        RECT 75.315 -210.965 75.645 -210.635 ;
        RECT 75.315 -212.325 75.645 -211.995 ;
        RECT 75.315 -213.685 75.645 -213.355 ;
        RECT 75.315 -215.045 75.645 -214.715 ;
        RECT 75.315 -216.405 75.645 -216.075 ;
        RECT 75.315 -217.765 75.645 -217.435 ;
        RECT 75.315 -219.125 75.645 -218.795 ;
        RECT 75.315 -221.37 75.645 -220.24 ;
        RECT 75.32 -221.485 75.64 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.51 -121.535 76.84 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.675 129.8 77.005 130.93 ;
        RECT 76.675 127.675 77.005 128.005 ;
        RECT 76.675 126.315 77.005 126.645 ;
        RECT 76.675 124.955 77.005 125.285 ;
        RECT 76.675 123.595 77.005 123.925 ;
        RECT 76.68 123.595 77 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.035 129.8 78.365 130.93 ;
        RECT 78.035 127.675 78.365 128.005 ;
        RECT 78.035 126.315 78.365 126.645 ;
        RECT 78.035 124.955 78.365 125.285 ;
        RECT 78.035 123.595 78.365 123.925 ;
        RECT 78.04 123.595 78.36 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.035 -1.525 78.365 -1.195 ;
        RECT 78.035 -2.885 78.365 -2.555 ;
        RECT 78.04 -3.56 78.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.035 -178.325 78.365 -177.995 ;
        RECT 78.035 -179.685 78.365 -179.355 ;
        RECT 78.035 -181.045 78.365 -180.715 ;
        RECT 78.035 -182.405 78.365 -182.075 ;
        RECT 78.035 -183.765 78.365 -183.435 ;
        RECT 78.035 -185.125 78.365 -184.795 ;
        RECT 78.035 -186.485 78.365 -186.155 ;
        RECT 78.035 -187.845 78.365 -187.515 ;
        RECT 78.035 -189.205 78.365 -188.875 ;
        RECT 78.035 -190.565 78.365 -190.235 ;
        RECT 78.035 -191.925 78.365 -191.595 ;
        RECT 78.035 -193.285 78.365 -192.955 ;
        RECT 78.035 -194.645 78.365 -194.315 ;
        RECT 78.035 -196.005 78.365 -195.675 ;
        RECT 78.035 -197.365 78.365 -197.035 ;
        RECT 78.035 -198.725 78.365 -198.395 ;
        RECT 78.035 -200.085 78.365 -199.755 ;
        RECT 78.035 -201.445 78.365 -201.115 ;
        RECT 78.035 -202.805 78.365 -202.475 ;
        RECT 78.035 -204.165 78.365 -203.835 ;
        RECT 78.035 -205.525 78.365 -205.195 ;
        RECT 78.035 -206.885 78.365 -206.555 ;
        RECT 78.035 -208.245 78.365 -207.915 ;
        RECT 78.035 -209.605 78.365 -209.275 ;
        RECT 78.035 -210.965 78.365 -210.635 ;
        RECT 78.035 -212.325 78.365 -211.995 ;
        RECT 78.035 -213.685 78.365 -213.355 ;
        RECT 78.035 -215.045 78.365 -214.715 ;
        RECT 78.035 -216.405 78.365 -216.075 ;
        RECT 78.035 -217.765 78.365 -217.435 ;
        RECT 78.035 -219.125 78.365 -218.795 ;
        RECT 78.035 -221.37 78.365 -220.24 ;
        RECT 78.04 -221.485 78.36 -118.155 ;
        RECT 78.035 -118.485 78.365 -118.155 ;
        RECT 78.035 -119.845 78.365 -119.515 ;
        RECT 78.035 -121.205 78.365 -120.875 ;
        RECT 78.035 -122.565 78.365 -122.235 ;
        RECT 78.035 -123.925 78.365 -123.595 ;
        RECT 78.035 -125.285 78.365 -124.955 ;
        RECT 78.035 -126.645 78.365 -126.315 ;
        RECT 78.035 -128.005 78.365 -127.675 ;
        RECT 78.035 -129.365 78.365 -129.035 ;
        RECT 78.035 -130.725 78.365 -130.395 ;
        RECT 78.035 -132.085 78.365 -131.755 ;
        RECT 78.035 -133.445 78.365 -133.115 ;
        RECT 78.035 -134.805 78.365 -134.475 ;
        RECT 78.035 -136.165 78.365 -135.835 ;
        RECT 78.035 -137.525 78.365 -137.195 ;
        RECT 78.035 -138.885 78.365 -138.555 ;
        RECT 78.035 -140.245 78.365 -139.915 ;
        RECT 78.035 -141.605 78.365 -141.275 ;
        RECT 78.035 -142.965 78.365 -142.635 ;
        RECT 78.035 -144.325 78.365 -143.995 ;
        RECT 78.035 -145.685 78.365 -145.355 ;
        RECT 78.035 -147.045 78.365 -146.715 ;
        RECT 78.035 -148.405 78.365 -148.075 ;
        RECT 78.035 -149.765 78.365 -149.435 ;
        RECT 78.035 -151.125 78.365 -150.795 ;
        RECT 78.035 -152.485 78.365 -152.155 ;
        RECT 78.035 -153.845 78.365 -153.515 ;
        RECT 78.035 -155.205 78.365 -154.875 ;
        RECT 78.035 -156.565 78.365 -156.235 ;
        RECT 78.035 -157.925 78.365 -157.595 ;
        RECT 78.035 -159.285 78.365 -158.955 ;
        RECT 78.035 -160.645 78.365 -160.315 ;
        RECT 78.035 -162.005 78.365 -161.675 ;
        RECT 78.035 -163.365 78.365 -163.035 ;
        RECT 78.035 -164.725 78.365 -164.395 ;
        RECT 78.035 -166.085 78.365 -165.755 ;
        RECT 78.035 -167.445 78.365 -167.115 ;
        RECT 78.035 -168.805 78.365 -168.475 ;
        RECT 78.035 -170.165 78.365 -169.835 ;
        RECT 78.035 -171.525 78.365 -171.195 ;
        RECT 78.035 -172.885 78.365 -172.555 ;
        RECT 78.035 -174.245 78.365 -173.915 ;
        RECT 78.035 -175.605 78.365 -175.275 ;
        RECT 78.035 -176.965 78.365 -176.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.61 -121.535 21.94 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.275 129.8 22.605 130.93 ;
        RECT 22.275 127.675 22.605 128.005 ;
        RECT 22.275 126.315 22.605 126.645 ;
        RECT 22.275 124.955 22.605 125.285 ;
        RECT 22.275 123.595 22.605 123.925 ;
        RECT 22.28 123.595 22.6 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.635 129.8 23.965 130.93 ;
        RECT 23.635 127.675 23.965 128.005 ;
        RECT 23.635 126.315 23.965 126.645 ;
        RECT 23.635 124.955 23.965 125.285 ;
        RECT 23.635 123.595 23.965 123.925 ;
        RECT 23.64 123.595 23.96 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.635 -1.525 23.965 -1.195 ;
        RECT 23.635 -2.885 23.965 -2.555 ;
        RECT 23.64 -3.56 23.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.995 129.8 25.325 130.93 ;
        RECT 24.995 127.675 25.325 128.005 ;
        RECT 24.995 126.315 25.325 126.645 ;
        RECT 24.995 124.955 25.325 125.285 ;
        RECT 24.995 123.595 25.325 123.925 ;
        RECT 25 123.595 25.32 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.995 -1.525 25.325 -1.195 ;
        RECT 24.995 -2.885 25.325 -2.555 ;
        RECT 25 -3.56 25.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.995 -118.485 25.325 -118.155 ;
        RECT 24.995 -119.845 25.325 -119.515 ;
        RECT 24.995 -121.205 25.325 -120.875 ;
        RECT 24.995 -122.565 25.325 -122.235 ;
        RECT 24.995 -123.925 25.325 -123.595 ;
        RECT 24.995 -125.285 25.325 -124.955 ;
        RECT 24.995 -126.645 25.325 -126.315 ;
        RECT 24.995 -128.005 25.325 -127.675 ;
        RECT 24.995 -129.365 25.325 -129.035 ;
        RECT 24.995 -130.725 25.325 -130.395 ;
        RECT 24.995 -132.085 25.325 -131.755 ;
        RECT 24.995 -133.445 25.325 -133.115 ;
        RECT 24.995 -134.805 25.325 -134.475 ;
        RECT 24.995 -136.165 25.325 -135.835 ;
        RECT 24.995 -137.525 25.325 -137.195 ;
        RECT 24.995 -138.885 25.325 -138.555 ;
        RECT 24.995 -140.245 25.325 -139.915 ;
        RECT 24.995 -141.605 25.325 -141.275 ;
        RECT 24.995 -142.965 25.325 -142.635 ;
        RECT 24.995 -144.325 25.325 -143.995 ;
        RECT 24.995 -145.685 25.325 -145.355 ;
        RECT 24.995 -147.045 25.325 -146.715 ;
        RECT 24.995 -148.405 25.325 -148.075 ;
        RECT 24.995 -149.765 25.325 -149.435 ;
        RECT 24.995 -151.125 25.325 -150.795 ;
        RECT 24.995 -152.485 25.325 -152.155 ;
        RECT 24.995 -153.845 25.325 -153.515 ;
        RECT 24.995 -155.205 25.325 -154.875 ;
        RECT 24.995 -156.565 25.325 -156.235 ;
        RECT 24.995 -157.925 25.325 -157.595 ;
        RECT 24.995 -159.285 25.325 -158.955 ;
        RECT 24.995 -160.645 25.325 -160.315 ;
        RECT 24.995 -162.005 25.325 -161.675 ;
        RECT 24.995 -163.365 25.325 -163.035 ;
        RECT 24.995 -164.725 25.325 -164.395 ;
        RECT 24.995 -166.085 25.325 -165.755 ;
        RECT 24.995 -167.445 25.325 -167.115 ;
        RECT 24.995 -168.805 25.325 -168.475 ;
        RECT 24.995 -170.165 25.325 -169.835 ;
        RECT 24.995 -171.525 25.325 -171.195 ;
        RECT 24.995 -172.885 25.325 -172.555 ;
        RECT 24.995 -174.245 25.325 -173.915 ;
        RECT 24.995 -175.605 25.325 -175.275 ;
        RECT 24.995 -176.965 25.325 -176.635 ;
        RECT 24.995 -178.325 25.325 -177.995 ;
        RECT 24.995 -179.685 25.325 -179.355 ;
        RECT 24.995 -181.045 25.325 -180.715 ;
        RECT 24.995 -182.405 25.325 -182.075 ;
        RECT 24.995 -183.765 25.325 -183.435 ;
        RECT 24.995 -185.125 25.325 -184.795 ;
        RECT 24.995 -186.485 25.325 -186.155 ;
        RECT 24.995 -187.845 25.325 -187.515 ;
        RECT 24.995 -189.205 25.325 -188.875 ;
        RECT 24.995 -190.565 25.325 -190.235 ;
        RECT 24.995 -191.925 25.325 -191.595 ;
        RECT 24.995 -193.285 25.325 -192.955 ;
        RECT 24.995 -194.645 25.325 -194.315 ;
        RECT 24.995 -196.005 25.325 -195.675 ;
        RECT 24.995 -197.365 25.325 -197.035 ;
        RECT 24.995 -198.725 25.325 -198.395 ;
        RECT 24.995 -200.085 25.325 -199.755 ;
        RECT 24.995 -201.445 25.325 -201.115 ;
        RECT 24.995 -202.805 25.325 -202.475 ;
        RECT 24.995 -204.165 25.325 -203.835 ;
        RECT 24.995 -205.525 25.325 -205.195 ;
        RECT 24.995 -206.885 25.325 -206.555 ;
        RECT 24.995 -208.245 25.325 -207.915 ;
        RECT 24.995 -209.605 25.325 -209.275 ;
        RECT 24.995 -210.965 25.325 -210.635 ;
        RECT 24.995 -212.325 25.325 -211.995 ;
        RECT 24.995 -213.685 25.325 -213.355 ;
        RECT 24.995 -215.045 25.325 -214.715 ;
        RECT 24.995 -216.405 25.325 -216.075 ;
        RECT 24.995 -217.765 25.325 -217.435 ;
        RECT 24.995 -219.125 25.325 -218.795 ;
        RECT 24.995 -221.37 25.325 -220.24 ;
        RECT 25 -221.485 25.32 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.355 129.8 26.685 130.93 ;
        RECT 26.355 127.675 26.685 128.005 ;
        RECT 26.355 126.315 26.685 126.645 ;
        RECT 26.355 124.955 26.685 125.285 ;
        RECT 26.355 123.595 26.685 123.925 ;
        RECT 26.36 123.595 26.68 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.355 -1.525 26.685 -1.195 ;
        RECT 26.355 -2.885 26.685 -2.555 ;
        RECT 26.36 -3.56 26.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.355 -118.485 26.685 -118.155 ;
        RECT 26.355 -119.845 26.685 -119.515 ;
        RECT 26.355 -121.205 26.685 -120.875 ;
        RECT 26.355 -122.565 26.685 -122.235 ;
        RECT 26.355 -123.925 26.685 -123.595 ;
        RECT 26.355 -125.285 26.685 -124.955 ;
        RECT 26.355 -126.645 26.685 -126.315 ;
        RECT 26.355 -128.005 26.685 -127.675 ;
        RECT 26.355 -129.365 26.685 -129.035 ;
        RECT 26.355 -130.725 26.685 -130.395 ;
        RECT 26.355 -132.085 26.685 -131.755 ;
        RECT 26.355 -133.445 26.685 -133.115 ;
        RECT 26.355 -134.805 26.685 -134.475 ;
        RECT 26.355 -136.165 26.685 -135.835 ;
        RECT 26.355 -137.525 26.685 -137.195 ;
        RECT 26.355 -138.885 26.685 -138.555 ;
        RECT 26.355 -140.245 26.685 -139.915 ;
        RECT 26.355 -141.605 26.685 -141.275 ;
        RECT 26.355 -142.965 26.685 -142.635 ;
        RECT 26.355 -144.325 26.685 -143.995 ;
        RECT 26.355 -145.685 26.685 -145.355 ;
        RECT 26.355 -147.045 26.685 -146.715 ;
        RECT 26.355 -148.405 26.685 -148.075 ;
        RECT 26.355 -149.765 26.685 -149.435 ;
        RECT 26.355 -151.125 26.685 -150.795 ;
        RECT 26.355 -152.485 26.685 -152.155 ;
        RECT 26.355 -153.845 26.685 -153.515 ;
        RECT 26.355 -155.205 26.685 -154.875 ;
        RECT 26.355 -156.565 26.685 -156.235 ;
        RECT 26.355 -157.925 26.685 -157.595 ;
        RECT 26.355 -159.285 26.685 -158.955 ;
        RECT 26.355 -160.645 26.685 -160.315 ;
        RECT 26.355 -162.005 26.685 -161.675 ;
        RECT 26.355 -163.365 26.685 -163.035 ;
        RECT 26.355 -164.725 26.685 -164.395 ;
        RECT 26.355 -166.085 26.685 -165.755 ;
        RECT 26.355 -167.445 26.685 -167.115 ;
        RECT 26.355 -168.805 26.685 -168.475 ;
        RECT 26.355 -170.165 26.685 -169.835 ;
        RECT 26.355 -171.525 26.685 -171.195 ;
        RECT 26.355 -172.885 26.685 -172.555 ;
        RECT 26.355 -174.245 26.685 -173.915 ;
        RECT 26.355 -175.605 26.685 -175.275 ;
        RECT 26.355 -176.965 26.685 -176.635 ;
        RECT 26.355 -178.325 26.685 -177.995 ;
        RECT 26.355 -179.685 26.685 -179.355 ;
        RECT 26.355 -181.045 26.685 -180.715 ;
        RECT 26.355 -182.405 26.685 -182.075 ;
        RECT 26.355 -183.765 26.685 -183.435 ;
        RECT 26.355 -185.125 26.685 -184.795 ;
        RECT 26.355 -186.485 26.685 -186.155 ;
        RECT 26.355 -187.845 26.685 -187.515 ;
        RECT 26.355 -189.205 26.685 -188.875 ;
        RECT 26.355 -190.565 26.685 -190.235 ;
        RECT 26.355 -191.925 26.685 -191.595 ;
        RECT 26.355 -193.285 26.685 -192.955 ;
        RECT 26.355 -194.645 26.685 -194.315 ;
        RECT 26.355 -196.005 26.685 -195.675 ;
        RECT 26.355 -197.365 26.685 -197.035 ;
        RECT 26.355 -198.725 26.685 -198.395 ;
        RECT 26.355 -200.085 26.685 -199.755 ;
        RECT 26.355 -201.445 26.685 -201.115 ;
        RECT 26.355 -202.805 26.685 -202.475 ;
        RECT 26.355 -204.165 26.685 -203.835 ;
        RECT 26.355 -205.525 26.685 -205.195 ;
        RECT 26.355 -206.885 26.685 -206.555 ;
        RECT 26.355 -208.245 26.685 -207.915 ;
        RECT 26.355 -209.605 26.685 -209.275 ;
        RECT 26.355 -210.965 26.685 -210.635 ;
        RECT 26.355 -212.325 26.685 -211.995 ;
        RECT 26.355 -213.685 26.685 -213.355 ;
        RECT 26.355 -215.045 26.685 -214.715 ;
        RECT 26.355 -216.405 26.685 -216.075 ;
        RECT 26.355 -217.765 26.685 -217.435 ;
        RECT 26.355 -219.125 26.685 -218.795 ;
        RECT 26.355 -221.37 26.685 -220.24 ;
        RECT 26.36 -221.485 26.68 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.71 -121.535 28.04 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.715 129.8 28.045 130.93 ;
        RECT 27.715 127.675 28.045 128.005 ;
        RECT 27.715 126.315 28.045 126.645 ;
        RECT 27.715 124.955 28.045 125.285 ;
        RECT 27.715 123.595 28.045 123.925 ;
        RECT 27.72 123.595 28.04 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.715 -122.565 28.045 -122.235 ;
        RECT 27.715 -123.925 28.045 -123.595 ;
        RECT 27.715 -125.285 28.045 -124.955 ;
        RECT 27.715 -126.645 28.045 -126.315 ;
        RECT 27.715 -128.005 28.045 -127.675 ;
        RECT 27.715 -129.365 28.045 -129.035 ;
        RECT 27.715 -130.725 28.045 -130.395 ;
        RECT 27.715 -132.085 28.045 -131.755 ;
        RECT 27.715 -133.445 28.045 -133.115 ;
        RECT 27.715 -134.805 28.045 -134.475 ;
        RECT 27.715 -136.165 28.045 -135.835 ;
        RECT 27.715 -137.525 28.045 -137.195 ;
        RECT 27.715 -138.885 28.045 -138.555 ;
        RECT 27.715 -140.245 28.045 -139.915 ;
        RECT 27.715 -141.605 28.045 -141.275 ;
        RECT 27.715 -142.965 28.045 -142.635 ;
        RECT 27.715 -144.325 28.045 -143.995 ;
        RECT 27.715 -145.685 28.045 -145.355 ;
        RECT 27.715 -147.045 28.045 -146.715 ;
        RECT 27.715 -148.405 28.045 -148.075 ;
        RECT 27.715 -149.765 28.045 -149.435 ;
        RECT 27.715 -151.125 28.045 -150.795 ;
        RECT 27.715 -152.485 28.045 -152.155 ;
        RECT 27.715 -153.845 28.045 -153.515 ;
        RECT 27.715 -155.205 28.045 -154.875 ;
        RECT 27.715 -156.565 28.045 -156.235 ;
        RECT 27.715 -157.925 28.045 -157.595 ;
        RECT 27.715 -159.285 28.045 -158.955 ;
        RECT 27.715 -160.645 28.045 -160.315 ;
        RECT 27.715 -162.005 28.045 -161.675 ;
        RECT 27.715 -163.365 28.045 -163.035 ;
        RECT 27.715 -164.725 28.045 -164.395 ;
        RECT 27.715 -166.085 28.045 -165.755 ;
        RECT 27.715 -167.445 28.045 -167.115 ;
        RECT 27.715 -168.805 28.045 -168.475 ;
        RECT 27.715 -170.165 28.045 -169.835 ;
        RECT 27.715 -171.525 28.045 -171.195 ;
        RECT 27.715 -172.885 28.045 -172.555 ;
        RECT 27.715 -174.245 28.045 -173.915 ;
        RECT 27.715 -175.605 28.045 -175.275 ;
        RECT 27.715 -176.965 28.045 -176.635 ;
        RECT 27.715 -178.325 28.045 -177.995 ;
        RECT 27.715 -179.685 28.045 -179.355 ;
        RECT 27.715 -181.045 28.045 -180.715 ;
        RECT 27.715 -182.405 28.045 -182.075 ;
        RECT 27.715 -183.765 28.045 -183.435 ;
        RECT 27.715 -185.125 28.045 -184.795 ;
        RECT 27.715 -186.485 28.045 -186.155 ;
        RECT 27.715 -187.845 28.045 -187.515 ;
        RECT 27.715 -189.205 28.045 -188.875 ;
        RECT 27.715 -190.565 28.045 -190.235 ;
        RECT 27.715 -191.925 28.045 -191.595 ;
        RECT 27.715 -193.285 28.045 -192.955 ;
        RECT 27.715 -194.645 28.045 -194.315 ;
        RECT 27.715 -196.005 28.045 -195.675 ;
        RECT 27.715 -197.365 28.045 -197.035 ;
        RECT 27.715 -198.725 28.045 -198.395 ;
        RECT 27.715 -200.085 28.045 -199.755 ;
        RECT 27.715 -201.445 28.045 -201.115 ;
        RECT 27.715 -202.805 28.045 -202.475 ;
        RECT 27.715 -204.165 28.045 -203.835 ;
        RECT 27.715 -205.525 28.045 -205.195 ;
        RECT 27.715 -206.885 28.045 -206.555 ;
        RECT 27.715 -208.245 28.045 -207.915 ;
        RECT 27.715 -209.605 28.045 -209.275 ;
        RECT 27.715 -210.965 28.045 -210.635 ;
        RECT 27.715 -212.325 28.045 -211.995 ;
        RECT 27.715 -213.685 28.045 -213.355 ;
        RECT 27.715 -215.045 28.045 -214.715 ;
        RECT 27.715 -216.405 28.045 -216.075 ;
        RECT 27.715 -217.765 28.045 -217.435 ;
        RECT 27.715 -219.125 28.045 -218.795 ;
        RECT 27.715 -221.37 28.045 -220.24 ;
        RECT 27.72 -221.485 28.04 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.075 129.8 29.405 130.93 ;
        RECT 29.075 127.675 29.405 128.005 ;
        RECT 29.075 126.315 29.405 126.645 ;
        RECT 29.075 124.955 29.405 125.285 ;
        RECT 29.075 123.595 29.405 123.925 ;
        RECT 29.08 123.595 29.4 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.075 -1.525 29.405 -1.195 ;
        RECT 29.075 -2.885 29.405 -2.555 ;
        RECT 29.08 -3.56 29.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.435 129.8 30.765 130.93 ;
        RECT 30.435 127.675 30.765 128.005 ;
        RECT 30.435 126.315 30.765 126.645 ;
        RECT 30.435 124.955 30.765 125.285 ;
        RECT 30.435 123.595 30.765 123.925 ;
        RECT 30.44 123.595 30.76 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.435 -1.525 30.765 -1.195 ;
        RECT 30.435 -2.885 30.765 -2.555 ;
        RECT 30.44 -3.56 30.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.795 129.8 32.125 130.93 ;
        RECT 31.795 127.675 32.125 128.005 ;
        RECT 31.795 126.315 32.125 126.645 ;
        RECT 31.795 124.955 32.125 125.285 ;
        RECT 31.795 123.595 32.125 123.925 ;
        RECT 31.8 123.595 32.12 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.795 -1.525 32.125 -1.195 ;
        RECT 31.795 -2.885 32.125 -2.555 ;
        RECT 31.8 -3.56 32.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.795 -118.485 32.125 -118.155 ;
        RECT 31.795 -119.845 32.125 -119.515 ;
        RECT 31.795 -121.205 32.125 -120.875 ;
        RECT 31.795 -122.565 32.125 -122.235 ;
        RECT 31.795 -123.925 32.125 -123.595 ;
        RECT 31.795 -125.285 32.125 -124.955 ;
        RECT 31.795 -126.645 32.125 -126.315 ;
        RECT 31.795 -128.005 32.125 -127.675 ;
        RECT 31.795 -129.365 32.125 -129.035 ;
        RECT 31.795 -130.725 32.125 -130.395 ;
        RECT 31.795 -132.085 32.125 -131.755 ;
        RECT 31.795 -133.445 32.125 -133.115 ;
        RECT 31.795 -134.805 32.125 -134.475 ;
        RECT 31.795 -136.165 32.125 -135.835 ;
        RECT 31.795 -137.525 32.125 -137.195 ;
        RECT 31.795 -138.885 32.125 -138.555 ;
        RECT 31.795 -140.245 32.125 -139.915 ;
        RECT 31.795 -141.605 32.125 -141.275 ;
        RECT 31.795 -142.965 32.125 -142.635 ;
        RECT 31.795 -144.325 32.125 -143.995 ;
        RECT 31.795 -145.685 32.125 -145.355 ;
        RECT 31.795 -147.045 32.125 -146.715 ;
        RECT 31.795 -148.405 32.125 -148.075 ;
        RECT 31.795 -149.765 32.125 -149.435 ;
        RECT 31.795 -151.125 32.125 -150.795 ;
        RECT 31.795 -152.485 32.125 -152.155 ;
        RECT 31.795 -153.845 32.125 -153.515 ;
        RECT 31.795 -155.205 32.125 -154.875 ;
        RECT 31.795 -156.565 32.125 -156.235 ;
        RECT 31.795 -157.925 32.125 -157.595 ;
        RECT 31.795 -159.285 32.125 -158.955 ;
        RECT 31.795 -160.645 32.125 -160.315 ;
        RECT 31.795 -162.005 32.125 -161.675 ;
        RECT 31.795 -163.365 32.125 -163.035 ;
        RECT 31.795 -164.725 32.125 -164.395 ;
        RECT 31.795 -166.085 32.125 -165.755 ;
        RECT 31.795 -167.445 32.125 -167.115 ;
        RECT 31.795 -168.805 32.125 -168.475 ;
        RECT 31.795 -170.165 32.125 -169.835 ;
        RECT 31.795 -171.525 32.125 -171.195 ;
        RECT 31.795 -172.885 32.125 -172.555 ;
        RECT 31.795 -174.245 32.125 -173.915 ;
        RECT 31.795 -175.605 32.125 -175.275 ;
        RECT 31.795 -176.965 32.125 -176.635 ;
        RECT 31.795 -178.325 32.125 -177.995 ;
        RECT 31.795 -179.685 32.125 -179.355 ;
        RECT 31.795 -181.045 32.125 -180.715 ;
        RECT 31.795 -182.405 32.125 -182.075 ;
        RECT 31.795 -183.765 32.125 -183.435 ;
        RECT 31.795 -185.125 32.125 -184.795 ;
        RECT 31.795 -186.485 32.125 -186.155 ;
        RECT 31.795 -187.845 32.125 -187.515 ;
        RECT 31.795 -189.205 32.125 -188.875 ;
        RECT 31.795 -190.565 32.125 -190.235 ;
        RECT 31.795 -191.925 32.125 -191.595 ;
        RECT 31.795 -193.285 32.125 -192.955 ;
        RECT 31.795 -194.645 32.125 -194.315 ;
        RECT 31.795 -196.005 32.125 -195.675 ;
        RECT 31.795 -197.365 32.125 -197.035 ;
        RECT 31.795 -198.725 32.125 -198.395 ;
        RECT 31.795 -200.085 32.125 -199.755 ;
        RECT 31.795 -201.445 32.125 -201.115 ;
        RECT 31.795 -202.805 32.125 -202.475 ;
        RECT 31.795 -204.165 32.125 -203.835 ;
        RECT 31.795 -205.525 32.125 -205.195 ;
        RECT 31.795 -206.885 32.125 -206.555 ;
        RECT 31.795 -208.245 32.125 -207.915 ;
        RECT 31.795 -209.605 32.125 -209.275 ;
        RECT 31.795 -210.965 32.125 -210.635 ;
        RECT 31.795 -212.325 32.125 -211.995 ;
        RECT 31.795 -213.685 32.125 -213.355 ;
        RECT 31.795 -215.045 32.125 -214.715 ;
        RECT 31.795 -216.405 32.125 -216.075 ;
        RECT 31.795 -217.765 32.125 -217.435 ;
        RECT 31.795 -219.125 32.125 -218.795 ;
        RECT 31.795 -221.37 32.125 -220.24 ;
        RECT 31.8 -221.485 32.12 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.155 129.8 33.485 130.93 ;
        RECT 33.155 127.675 33.485 128.005 ;
        RECT 33.155 126.315 33.485 126.645 ;
        RECT 33.155 124.955 33.485 125.285 ;
        RECT 33.155 123.595 33.485 123.925 ;
        RECT 33.16 123.595 33.48 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.155 -122.565 33.485 -122.235 ;
        RECT 33.155 -123.925 33.485 -123.595 ;
        RECT 33.155 -125.285 33.485 -124.955 ;
        RECT 33.155 -126.645 33.485 -126.315 ;
        RECT 33.155 -128.005 33.485 -127.675 ;
        RECT 33.155 -129.365 33.485 -129.035 ;
        RECT 33.155 -130.725 33.485 -130.395 ;
        RECT 33.155 -132.085 33.485 -131.755 ;
        RECT 33.155 -133.445 33.485 -133.115 ;
        RECT 33.155 -134.805 33.485 -134.475 ;
        RECT 33.155 -136.165 33.485 -135.835 ;
        RECT 33.155 -137.525 33.485 -137.195 ;
        RECT 33.155 -138.885 33.485 -138.555 ;
        RECT 33.155 -140.245 33.485 -139.915 ;
        RECT 33.155 -141.605 33.485 -141.275 ;
        RECT 33.155 -142.965 33.485 -142.635 ;
        RECT 33.155 -144.325 33.485 -143.995 ;
        RECT 33.155 -145.685 33.485 -145.355 ;
        RECT 33.155 -147.045 33.485 -146.715 ;
        RECT 33.155 -148.405 33.485 -148.075 ;
        RECT 33.155 -149.765 33.485 -149.435 ;
        RECT 33.155 -151.125 33.485 -150.795 ;
        RECT 33.155 -152.485 33.485 -152.155 ;
        RECT 33.155 -153.845 33.485 -153.515 ;
        RECT 33.155 -155.205 33.485 -154.875 ;
        RECT 33.155 -156.565 33.485 -156.235 ;
        RECT 33.155 -157.925 33.485 -157.595 ;
        RECT 33.155 -159.285 33.485 -158.955 ;
        RECT 33.155 -160.645 33.485 -160.315 ;
        RECT 33.155 -162.005 33.485 -161.675 ;
        RECT 33.155 -163.365 33.485 -163.035 ;
        RECT 33.155 -164.725 33.485 -164.395 ;
        RECT 33.155 -166.085 33.485 -165.755 ;
        RECT 33.155 -167.445 33.485 -167.115 ;
        RECT 33.155 -168.805 33.485 -168.475 ;
        RECT 33.155 -170.165 33.485 -169.835 ;
        RECT 33.155 -171.525 33.485 -171.195 ;
        RECT 33.155 -172.885 33.485 -172.555 ;
        RECT 33.155 -174.245 33.485 -173.915 ;
        RECT 33.155 -175.605 33.485 -175.275 ;
        RECT 33.155 -176.965 33.485 -176.635 ;
        RECT 33.155 -178.325 33.485 -177.995 ;
        RECT 33.155 -179.685 33.485 -179.355 ;
        RECT 33.155 -181.045 33.485 -180.715 ;
        RECT 33.155 -182.405 33.485 -182.075 ;
        RECT 33.155 -183.765 33.485 -183.435 ;
        RECT 33.155 -185.125 33.485 -184.795 ;
        RECT 33.155 -186.485 33.485 -186.155 ;
        RECT 33.155 -187.845 33.485 -187.515 ;
        RECT 33.155 -189.205 33.485 -188.875 ;
        RECT 33.155 -190.565 33.485 -190.235 ;
        RECT 33.155 -191.925 33.485 -191.595 ;
        RECT 33.155 -193.285 33.485 -192.955 ;
        RECT 33.155 -194.645 33.485 -194.315 ;
        RECT 33.155 -196.005 33.485 -195.675 ;
        RECT 33.155 -197.365 33.485 -197.035 ;
        RECT 33.155 -198.725 33.485 -198.395 ;
        RECT 33.155 -200.085 33.485 -199.755 ;
        RECT 33.155 -201.445 33.485 -201.115 ;
        RECT 33.155 -202.805 33.485 -202.475 ;
        RECT 33.155 -204.165 33.485 -203.835 ;
        RECT 33.155 -205.525 33.485 -205.195 ;
        RECT 33.155 -206.885 33.485 -206.555 ;
        RECT 33.155 -208.245 33.485 -207.915 ;
        RECT 33.155 -209.605 33.485 -209.275 ;
        RECT 33.155 -210.965 33.485 -210.635 ;
        RECT 33.155 -212.325 33.485 -211.995 ;
        RECT 33.155 -213.685 33.485 -213.355 ;
        RECT 33.155 -215.045 33.485 -214.715 ;
        RECT 33.155 -216.405 33.485 -216.075 ;
        RECT 33.155 -217.765 33.485 -217.435 ;
        RECT 33.155 -219.125 33.485 -218.795 ;
        RECT 33.155 -221.37 33.485 -220.24 ;
        RECT 33.16 -221.485 33.48 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.81 -121.535 34.14 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.515 129.8 34.845 130.93 ;
        RECT 34.515 127.675 34.845 128.005 ;
        RECT 34.515 126.315 34.845 126.645 ;
        RECT 34.515 124.955 34.845 125.285 ;
        RECT 34.515 123.595 34.845 123.925 ;
        RECT 34.52 123.595 34.84 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.515 -1.525 34.845 -1.195 ;
        RECT 34.515 -2.885 34.845 -2.555 ;
        RECT 34.52 -3.56 34.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.875 129.8 36.205 130.93 ;
        RECT 35.875 127.675 36.205 128.005 ;
        RECT 35.875 126.315 36.205 126.645 ;
        RECT 35.875 124.955 36.205 125.285 ;
        RECT 35.875 123.595 36.205 123.925 ;
        RECT 35.88 123.595 36.2 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.875 -1.525 36.205 -1.195 ;
        RECT 35.875 -2.885 36.205 -2.555 ;
        RECT 35.88 -3.56 36.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.235 129.8 37.565 130.93 ;
        RECT 37.235 127.675 37.565 128.005 ;
        RECT 37.235 126.315 37.565 126.645 ;
        RECT 37.235 124.955 37.565 125.285 ;
        RECT 37.235 123.595 37.565 123.925 ;
        RECT 37.24 123.595 37.56 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.235 -1.525 37.565 -1.195 ;
        RECT 37.235 -2.885 37.565 -2.555 ;
        RECT 37.24 -3.56 37.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.235 -118.485 37.565 -118.155 ;
        RECT 37.235 -119.845 37.565 -119.515 ;
        RECT 37.235 -121.205 37.565 -120.875 ;
        RECT 37.235 -122.565 37.565 -122.235 ;
        RECT 37.235 -123.925 37.565 -123.595 ;
        RECT 37.235 -125.285 37.565 -124.955 ;
        RECT 37.235 -126.645 37.565 -126.315 ;
        RECT 37.235 -128.005 37.565 -127.675 ;
        RECT 37.235 -129.365 37.565 -129.035 ;
        RECT 37.235 -130.725 37.565 -130.395 ;
        RECT 37.235 -132.085 37.565 -131.755 ;
        RECT 37.235 -133.445 37.565 -133.115 ;
        RECT 37.235 -134.805 37.565 -134.475 ;
        RECT 37.235 -136.165 37.565 -135.835 ;
        RECT 37.235 -137.525 37.565 -137.195 ;
        RECT 37.235 -138.885 37.565 -138.555 ;
        RECT 37.235 -140.245 37.565 -139.915 ;
        RECT 37.235 -141.605 37.565 -141.275 ;
        RECT 37.235 -142.965 37.565 -142.635 ;
        RECT 37.235 -144.325 37.565 -143.995 ;
        RECT 37.235 -145.685 37.565 -145.355 ;
        RECT 37.235 -147.045 37.565 -146.715 ;
        RECT 37.235 -148.405 37.565 -148.075 ;
        RECT 37.235 -149.765 37.565 -149.435 ;
        RECT 37.235 -151.125 37.565 -150.795 ;
        RECT 37.235 -152.485 37.565 -152.155 ;
        RECT 37.235 -153.845 37.565 -153.515 ;
        RECT 37.235 -155.205 37.565 -154.875 ;
        RECT 37.235 -156.565 37.565 -156.235 ;
        RECT 37.235 -157.925 37.565 -157.595 ;
        RECT 37.235 -159.285 37.565 -158.955 ;
        RECT 37.235 -160.645 37.565 -160.315 ;
        RECT 37.235 -162.005 37.565 -161.675 ;
        RECT 37.235 -163.365 37.565 -163.035 ;
        RECT 37.235 -164.725 37.565 -164.395 ;
        RECT 37.235 -166.085 37.565 -165.755 ;
        RECT 37.235 -167.445 37.565 -167.115 ;
        RECT 37.235 -168.805 37.565 -168.475 ;
        RECT 37.235 -170.165 37.565 -169.835 ;
        RECT 37.235 -171.525 37.565 -171.195 ;
        RECT 37.235 -172.885 37.565 -172.555 ;
        RECT 37.235 -174.245 37.565 -173.915 ;
        RECT 37.235 -175.605 37.565 -175.275 ;
        RECT 37.235 -176.965 37.565 -176.635 ;
        RECT 37.235 -178.325 37.565 -177.995 ;
        RECT 37.235 -179.685 37.565 -179.355 ;
        RECT 37.235 -181.045 37.565 -180.715 ;
        RECT 37.235 -182.405 37.565 -182.075 ;
        RECT 37.235 -183.765 37.565 -183.435 ;
        RECT 37.235 -185.125 37.565 -184.795 ;
        RECT 37.235 -186.485 37.565 -186.155 ;
        RECT 37.235 -187.845 37.565 -187.515 ;
        RECT 37.235 -189.205 37.565 -188.875 ;
        RECT 37.235 -190.565 37.565 -190.235 ;
        RECT 37.235 -191.925 37.565 -191.595 ;
        RECT 37.235 -193.285 37.565 -192.955 ;
        RECT 37.235 -194.645 37.565 -194.315 ;
        RECT 37.235 -196.005 37.565 -195.675 ;
        RECT 37.235 -197.365 37.565 -197.035 ;
        RECT 37.235 -198.725 37.565 -198.395 ;
        RECT 37.235 -200.085 37.565 -199.755 ;
        RECT 37.235 -201.445 37.565 -201.115 ;
        RECT 37.235 -202.805 37.565 -202.475 ;
        RECT 37.235 -204.165 37.565 -203.835 ;
        RECT 37.235 -205.525 37.565 -205.195 ;
        RECT 37.235 -206.885 37.565 -206.555 ;
        RECT 37.235 -208.245 37.565 -207.915 ;
        RECT 37.235 -209.605 37.565 -209.275 ;
        RECT 37.235 -210.965 37.565 -210.635 ;
        RECT 37.235 -212.325 37.565 -211.995 ;
        RECT 37.235 -213.685 37.565 -213.355 ;
        RECT 37.235 -215.045 37.565 -214.715 ;
        RECT 37.235 -216.405 37.565 -216.075 ;
        RECT 37.235 -217.765 37.565 -217.435 ;
        RECT 37.235 -219.125 37.565 -218.795 ;
        RECT 37.235 -221.37 37.565 -220.24 ;
        RECT 37.24 -221.485 37.56 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.595 129.8 38.925 130.93 ;
        RECT 38.595 127.675 38.925 128.005 ;
        RECT 38.595 126.315 38.925 126.645 ;
        RECT 38.595 124.955 38.925 125.285 ;
        RECT 38.595 123.595 38.925 123.925 ;
        RECT 38.6 123.595 38.92 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.595 -122.565 38.925 -122.235 ;
        RECT 38.595 -123.925 38.925 -123.595 ;
        RECT 38.595 -125.285 38.925 -124.955 ;
        RECT 38.595 -126.645 38.925 -126.315 ;
        RECT 38.595 -128.005 38.925 -127.675 ;
        RECT 38.595 -129.365 38.925 -129.035 ;
        RECT 38.595 -130.725 38.925 -130.395 ;
        RECT 38.595 -132.085 38.925 -131.755 ;
        RECT 38.595 -133.445 38.925 -133.115 ;
        RECT 38.595 -134.805 38.925 -134.475 ;
        RECT 38.595 -136.165 38.925 -135.835 ;
        RECT 38.595 -137.525 38.925 -137.195 ;
        RECT 38.595 -138.885 38.925 -138.555 ;
        RECT 38.595 -140.245 38.925 -139.915 ;
        RECT 38.595 -141.605 38.925 -141.275 ;
        RECT 38.595 -142.965 38.925 -142.635 ;
        RECT 38.595 -144.325 38.925 -143.995 ;
        RECT 38.595 -145.685 38.925 -145.355 ;
        RECT 38.595 -147.045 38.925 -146.715 ;
        RECT 38.595 -148.405 38.925 -148.075 ;
        RECT 38.595 -149.765 38.925 -149.435 ;
        RECT 38.595 -151.125 38.925 -150.795 ;
        RECT 38.595 -152.485 38.925 -152.155 ;
        RECT 38.595 -153.845 38.925 -153.515 ;
        RECT 38.595 -155.205 38.925 -154.875 ;
        RECT 38.595 -156.565 38.925 -156.235 ;
        RECT 38.595 -157.925 38.925 -157.595 ;
        RECT 38.595 -159.285 38.925 -158.955 ;
        RECT 38.595 -160.645 38.925 -160.315 ;
        RECT 38.595 -162.005 38.925 -161.675 ;
        RECT 38.595 -163.365 38.925 -163.035 ;
        RECT 38.595 -164.725 38.925 -164.395 ;
        RECT 38.595 -166.085 38.925 -165.755 ;
        RECT 38.595 -167.445 38.925 -167.115 ;
        RECT 38.595 -168.805 38.925 -168.475 ;
        RECT 38.595 -170.165 38.925 -169.835 ;
        RECT 38.595 -171.525 38.925 -171.195 ;
        RECT 38.595 -172.885 38.925 -172.555 ;
        RECT 38.595 -174.245 38.925 -173.915 ;
        RECT 38.595 -175.605 38.925 -175.275 ;
        RECT 38.595 -176.965 38.925 -176.635 ;
        RECT 38.595 -178.325 38.925 -177.995 ;
        RECT 38.595 -179.685 38.925 -179.355 ;
        RECT 38.595 -181.045 38.925 -180.715 ;
        RECT 38.595 -182.405 38.925 -182.075 ;
        RECT 38.595 -183.765 38.925 -183.435 ;
        RECT 38.595 -185.125 38.925 -184.795 ;
        RECT 38.595 -186.485 38.925 -186.155 ;
        RECT 38.595 -187.845 38.925 -187.515 ;
        RECT 38.595 -189.205 38.925 -188.875 ;
        RECT 38.595 -190.565 38.925 -190.235 ;
        RECT 38.595 -191.925 38.925 -191.595 ;
        RECT 38.595 -193.285 38.925 -192.955 ;
        RECT 38.595 -194.645 38.925 -194.315 ;
        RECT 38.595 -196.005 38.925 -195.675 ;
        RECT 38.595 -197.365 38.925 -197.035 ;
        RECT 38.595 -198.725 38.925 -198.395 ;
        RECT 38.595 -200.085 38.925 -199.755 ;
        RECT 38.595 -201.445 38.925 -201.115 ;
        RECT 38.595 -202.805 38.925 -202.475 ;
        RECT 38.595 -204.165 38.925 -203.835 ;
        RECT 38.595 -205.525 38.925 -205.195 ;
        RECT 38.595 -206.885 38.925 -206.555 ;
        RECT 38.595 -208.245 38.925 -207.915 ;
        RECT 38.595 -209.605 38.925 -209.275 ;
        RECT 38.595 -210.965 38.925 -210.635 ;
        RECT 38.595 -212.325 38.925 -211.995 ;
        RECT 38.595 -213.685 38.925 -213.355 ;
        RECT 38.595 -215.045 38.925 -214.715 ;
        RECT 38.595 -216.405 38.925 -216.075 ;
        RECT 38.595 -217.765 38.925 -217.435 ;
        RECT 38.595 -219.125 38.925 -218.795 ;
        RECT 38.595 -221.37 38.925 -220.24 ;
        RECT 38.6 -221.485 38.92 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.91 -121.535 40.24 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.955 129.8 40.285 130.93 ;
        RECT 39.955 127.675 40.285 128.005 ;
        RECT 39.955 126.315 40.285 126.645 ;
        RECT 39.955 124.955 40.285 125.285 ;
        RECT 39.955 123.595 40.285 123.925 ;
        RECT 39.96 123.595 40.28 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.315 129.8 41.645 130.93 ;
        RECT 41.315 127.675 41.645 128.005 ;
        RECT 41.315 126.315 41.645 126.645 ;
        RECT 41.315 124.955 41.645 125.285 ;
        RECT 41.315 123.595 41.645 123.925 ;
        RECT 41.32 123.595 41.64 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.315 -1.525 41.645 -1.195 ;
        RECT 41.315 -2.885 41.645 -2.555 ;
        RECT 41.32 -3.56 41.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.675 129.8 43.005 130.93 ;
        RECT 42.675 127.675 43.005 128.005 ;
        RECT 42.675 126.315 43.005 126.645 ;
        RECT 42.675 124.955 43.005 125.285 ;
        RECT 42.675 123.595 43.005 123.925 ;
        RECT 42.68 123.595 43 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.675 -1.525 43.005 -1.195 ;
        RECT 42.675 -2.885 43.005 -2.555 ;
        RECT 42.68 -3.56 43 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.035 129.8 44.365 130.93 ;
        RECT 44.035 127.675 44.365 128.005 ;
        RECT 44.035 126.315 44.365 126.645 ;
        RECT 44.035 124.955 44.365 125.285 ;
        RECT 44.035 123.595 44.365 123.925 ;
        RECT 44.04 123.595 44.36 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.035 -1.525 44.365 -1.195 ;
        RECT 44.035 -2.885 44.365 -2.555 ;
        RECT 44.04 -3.56 44.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.035 -118.485 44.365 -118.155 ;
        RECT 44.035 -119.845 44.365 -119.515 ;
        RECT 44.035 -121.205 44.365 -120.875 ;
        RECT 44.035 -122.565 44.365 -122.235 ;
        RECT 44.035 -123.925 44.365 -123.595 ;
        RECT 44.035 -125.285 44.365 -124.955 ;
        RECT 44.035 -126.645 44.365 -126.315 ;
        RECT 44.035 -128.005 44.365 -127.675 ;
        RECT 44.035 -129.365 44.365 -129.035 ;
        RECT 44.035 -130.725 44.365 -130.395 ;
        RECT 44.035 -132.085 44.365 -131.755 ;
        RECT 44.035 -133.445 44.365 -133.115 ;
        RECT 44.035 -134.805 44.365 -134.475 ;
        RECT 44.035 -136.165 44.365 -135.835 ;
        RECT 44.035 -137.525 44.365 -137.195 ;
        RECT 44.035 -138.885 44.365 -138.555 ;
        RECT 44.035 -140.245 44.365 -139.915 ;
        RECT 44.035 -141.605 44.365 -141.275 ;
        RECT 44.035 -142.965 44.365 -142.635 ;
        RECT 44.035 -144.325 44.365 -143.995 ;
        RECT 44.035 -145.685 44.365 -145.355 ;
        RECT 44.035 -147.045 44.365 -146.715 ;
        RECT 44.035 -148.405 44.365 -148.075 ;
        RECT 44.035 -149.765 44.365 -149.435 ;
        RECT 44.035 -151.125 44.365 -150.795 ;
        RECT 44.035 -152.485 44.365 -152.155 ;
        RECT 44.035 -153.845 44.365 -153.515 ;
        RECT 44.035 -155.205 44.365 -154.875 ;
        RECT 44.035 -156.565 44.365 -156.235 ;
        RECT 44.035 -157.925 44.365 -157.595 ;
        RECT 44.035 -159.285 44.365 -158.955 ;
        RECT 44.035 -160.645 44.365 -160.315 ;
        RECT 44.035 -162.005 44.365 -161.675 ;
        RECT 44.035 -163.365 44.365 -163.035 ;
        RECT 44.035 -164.725 44.365 -164.395 ;
        RECT 44.035 -166.085 44.365 -165.755 ;
        RECT 44.035 -167.445 44.365 -167.115 ;
        RECT 44.035 -168.805 44.365 -168.475 ;
        RECT 44.035 -170.165 44.365 -169.835 ;
        RECT 44.035 -171.525 44.365 -171.195 ;
        RECT 44.035 -172.885 44.365 -172.555 ;
        RECT 44.035 -174.245 44.365 -173.915 ;
        RECT 44.035 -175.605 44.365 -175.275 ;
        RECT 44.035 -176.965 44.365 -176.635 ;
        RECT 44.035 -178.325 44.365 -177.995 ;
        RECT 44.035 -179.685 44.365 -179.355 ;
        RECT 44.035 -181.045 44.365 -180.715 ;
        RECT 44.035 -182.405 44.365 -182.075 ;
        RECT 44.035 -183.765 44.365 -183.435 ;
        RECT 44.035 -185.125 44.365 -184.795 ;
        RECT 44.035 -186.485 44.365 -186.155 ;
        RECT 44.035 -187.845 44.365 -187.515 ;
        RECT 44.035 -189.205 44.365 -188.875 ;
        RECT 44.035 -190.565 44.365 -190.235 ;
        RECT 44.035 -191.925 44.365 -191.595 ;
        RECT 44.035 -193.285 44.365 -192.955 ;
        RECT 44.035 -194.645 44.365 -194.315 ;
        RECT 44.035 -196.005 44.365 -195.675 ;
        RECT 44.035 -197.365 44.365 -197.035 ;
        RECT 44.035 -198.725 44.365 -198.395 ;
        RECT 44.035 -200.085 44.365 -199.755 ;
        RECT 44.035 -201.445 44.365 -201.115 ;
        RECT 44.035 -202.805 44.365 -202.475 ;
        RECT 44.035 -204.165 44.365 -203.835 ;
        RECT 44.035 -205.525 44.365 -205.195 ;
        RECT 44.035 -206.885 44.365 -206.555 ;
        RECT 44.035 -208.245 44.365 -207.915 ;
        RECT 44.035 -209.605 44.365 -209.275 ;
        RECT 44.035 -210.965 44.365 -210.635 ;
        RECT 44.035 -212.325 44.365 -211.995 ;
        RECT 44.035 -213.685 44.365 -213.355 ;
        RECT 44.035 -215.045 44.365 -214.715 ;
        RECT 44.035 -216.405 44.365 -216.075 ;
        RECT 44.035 -217.765 44.365 -217.435 ;
        RECT 44.035 -219.125 44.365 -218.795 ;
        RECT 44.035 -221.37 44.365 -220.24 ;
        RECT 44.04 -221.485 44.36 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.395 129.8 45.725 130.93 ;
        RECT 45.395 127.675 45.725 128.005 ;
        RECT 45.395 126.315 45.725 126.645 ;
        RECT 45.395 124.955 45.725 125.285 ;
        RECT 45.395 123.595 45.725 123.925 ;
        RECT 45.4 123.595 45.72 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.395 -122.565 45.725 -122.235 ;
        RECT 45.395 -123.925 45.725 -123.595 ;
        RECT 45.395 -125.285 45.725 -124.955 ;
        RECT 45.395 -126.645 45.725 -126.315 ;
        RECT 45.395 -128.005 45.725 -127.675 ;
        RECT 45.395 -129.365 45.725 -129.035 ;
        RECT 45.395 -130.725 45.725 -130.395 ;
        RECT 45.395 -132.085 45.725 -131.755 ;
        RECT 45.395 -133.445 45.725 -133.115 ;
        RECT 45.395 -134.805 45.725 -134.475 ;
        RECT 45.395 -136.165 45.725 -135.835 ;
        RECT 45.395 -137.525 45.725 -137.195 ;
        RECT 45.395 -138.885 45.725 -138.555 ;
        RECT 45.395 -140.245 45.725 -139.915 ;
        RECT 45.395 -141.605 45.725 -141.275 ;
        RECT 45.395 -142.965 45.725 -142.635 ;
        RECT 45.395 -144.325 45.725 -143.995 ;
        RECT 45.395 -145.685 45.725 -145.355 ;
        RECT 45.395 -147.045 45.725 -146.715 ;
        RECT 45.395 -148.405 45.725 -148.075 ;
        RECT 45.395 -149.765 45.725 -149.435 ;
        RECT 45.395 -151.125 45.725 -150.795 ;
        RECT 45.395 -152.485 45.725 -152.155 ;
        RECT 45.395 -153.845 45.725 -153.515 ;
        RECT 45.395 -155.205 45.725 -154.875 ;
        RECT 45.395 -156.565 45.725 -156.235 ;
        RECT 45.395 -157.925 45.725 -157.595 ;
        RECT 45.395 -159.285 45.725 -158.955 ;
        RECT 45.395 -160.645 45.725 -160.315 ;
        RECT 45.395 -162.005 45.725 -161.675 ;
        RECT 45.395 -163.365 45.725 -163.035 ;
        RECT 45.395 -164.725 45.725 -164.395 ;
        RECT 45.395 -166.085 45.725 -165.755 ;
        RECT 45.395 -167.445 45.725 -167.115 ;
        RECT 45.395 -168.805 45.725 -168.475 ;
        RECT 45.395 -170.165 45.725 -169.835 ;
        RECT 45.395 -171.525 45.725 -171.195 ;
        RECT 45.395 -172.885 45.725 -172.555 ;
        RECT 45.395 -174.245 45.725 -173.915 ;
        RECT 45.395 -175.605 45.725 -175.275 ;
        RECT 45.395 -176.965 45.725 -176.635 ;
        RECT 45.395 -178.325 45.725 -177.995 ;
        RECT 45.395 -179.685 45.725 -179.355 ;
        RECT 45.395 -181.045 45.725 -180.715 ;
        RECT 45.395 -182.405 45.725 -182.075 ;
        RECT 45.395 -183.765 45.725 -183.435 ;
        RECT 45.395 -185.125 45.725 -184.795 ;
        RECT 45.395 -186.485 45.725 -186.155 ;
        RECT 45.395 -187.845 45.725 -187.515 ;
        RECT 45.395 -189.205 45.725 -188.875 ;
        RECT 45.395 -190.565 45.725 -190.235 ;
        RECT 45.395 -191.925 45.725 -191.595 ;
        RECT 45.395 -193.285 45.725 -192.955 ;
        RECT 45.395 -194.645 45.725 -194.315 ;
        RECT 45.395 -196.005 45.725 -195.675 ;
        RECT 45.395 -197.365 45.725 -197.035 ;
        RECT 45.395 -198.725 45.725 -198.395 ;
        RECT 45.395 -200.085 45.725 -199.755 ;
        RECT 45.395 -201.445 45.725 -201.115 ;
        RECT 45.395 -202.805 45.725 -202.475 ;
        RECT 45.395 -204.165 45.725 -203.835 ;
        RECT 45.395 -205.525 45.725 -205.195 ;
        RECT 45.395 -206.885 45.725 -206.555 ;
        RECT 45.395 -208.245 45.725 -207.915 ;
        RECT 45.395 -209.605 45.725 -209.275 ;
        RECT 45.395 -210.965 45.725 -210.635 ;
        RECT 45.395 -212.325 45.725 -211.995 ;
        RECT 45.395 -213.685 45.725 -213.355 ;
        RECT 45.395 -215.045 45.725 -214.715 ;
        RECT 45.395 -216.405 45.725 -216.075 ;
        RECT 45.395 -217.765 45.725 -217.435 ;
        RECT 45.395 -219.125 45.725 -218.795 ;
        RECT 45.395 -221.37 45.725 -220.24 ;
        RECT 45.4 -221.485 45.72 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.01 -121.535 46.34 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.755 129.8 47.085 130.93 ;
        RECT 46.755 127.675 47.085 128.005 ;
        RECT 46.755 126.315 47.085 126.645 ;
        RECT 46.755 124.955 47.085 125.285 ;
        RECT 46.755 123.595 47.085 123.925 ;
        RECT 46.76 123.595 47.08 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.755 -1.525 47.085 -1.195 ;
        RECT 46.755 -2.885 47.085 -2.555 ;
        RECT 46.76 -3.56 47.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.115 129.8 48.445 130.93 ;
        RECT 48.115 127.675 48.445 128.005 ;
        RECT 48.115 126.315 48.445 126.645 ;
        RECT 48.115 124.955 48.445 125.285 ;
        RECT 48.115 123.595 48.445 123.925 ;
        RECT 48.12 123.595 48.44 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.115 -1.525 48.445 -1.195 ;
        RECT 48.115 -2.885 48.445 -2.555 ;
        RECT 48.12 -3.56 48.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.475 129.8 49.805 130.93 ;
        RECT 49.475 127.675 49.805 128.005 ;
        RECT 49.475 126.315 49.805 126.645 ;
        RECT 49.475 124.955 49.805 125.285 ;
        RECT 49.475 123.595 49.805 123.925 ;
        RECT 49.48 123.595 49.8 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.475 -1.525 49.805 -1.195 ;
        RECT 49.475 -2.885 49.805 -2.555 ;
        RECT 49.48 -3.56 49.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.475 -118.485 49.805 -118.155 ;
        RECT 49.475 -119.845 49.805 -119.515 ;
        RECT 49.475 -121.205 49.805 -120.875 ;
        RECT 49.475 -122.565 49.805 -122.235 ;
        RECT 49.475 -123.925 49.805 -123.595 ;
        RECT 49.475 -125.285 49.805 -124.955 ;
        RECT 49.475 -126.645 49.805 -126.315 ;
        RECT 49.475 -128.005 49.805 -127.675 ;
        RECT 49.475 -129.365 49.805 -129.035 ;
        RECT 49.475 -130.725 49.805 -130.395 ;
        RECT 49.475 -132.085 49.805 -131.755 ;
        RECT 49.475 -133.445 49.805 -133.115 ;
        RECT 49.475 -134.805 49.805 -134.475 ;
        RECT 49.475 -136.165 49.805 -135.835 ;
        RECT 49.475 -137.525 49.805 -137.195 ;
        RECT 49.475 -138.885 49.805 -138.555 ;
        RECT 49.475 -140.245 49.805 -139.915 ;
        RECT 49.475 -141.605 49.805 -141.275 ;
        RECT 49.475 -142.965 49.805 -142.635 ;
        RECT 49.475 -144.325 49.805 -143.995 ;
        RECT 49.475 -145.685 49.805 -145.355 ;
        RECT 49.475 -147.045 49.805 -146.715 ;
        RECT 49.475 -148.405 49.805 -148.075 ;
        RECT 49.475 -149.765 49.805 -149.435 ;
        RECT 49.475 -151.125 49.805 -150.795 ;
        RECT 49.475 -152.485 49.805 -152.155 ;
        RECT 49.475 -153.845 49.805 -153.515 ;
        RECT 49.475 -155.205 49.805 -154.875 ;
        RECT 49.475 -156.565 49.805 -156.235 ;
        RECT 49.475 -157.925 49.805 -157.595 ;
        RECT 49.475 -159.285 49.805 -158.955 ;
        RECT 49.475 -160.645 49.805 -160.315 ;
        RECT 49.475 -162.005 49.805 -161.675 ;
        RECT 49.475 -163.365 49.805 -163.035 ;
        RECT 49.475 -164.725 49.805 -164.395 ;
        RECT 49.475 -166.085 49.805 -165.755 ;
        RECT 49.475 -167.445 49.805 -167.115 ;
        RECT 49.475 -168.805 49.805 -168.475 ;
        RECT 49.475 -170.165 49.805 -169.835 ;
        RECT 49.475 -171.525 49.805 -171.195 ;
        RECT 49.475 -172.885 49.805 -172.555 ;
        RECT 49.475 -174.245 49.805 -173.915 ;
        RECT 49.475 -175.605 49.805 -175.275 ;
        RECT 49.475 -176.965 49.805 -176.635 ;
        RECT 49.475 -178.325 49.805 -177.995 ;
        RECT 49.475 -179.685 49.805 -179.355 ;
        RECT 49.475 -181.045 49.805 -180.715 ;
        RECT 49.475 -182.405 49.805 -182.075 ;
        RECT 49.475 -183.765 49.805 -183.435 ;
        RECT 49.475 -185.125 49.805 -184.795 ;
        RECT 49.475 -186.485 49.805 -186.155 ;
        RECT 49.475 -187.845 49.805 -187.515 ;
        RECT 49.475 -189.205 49.805 -188.875 ;
        RECT 49.475 -190.565 49.805 -190.235 ;
        RECT 49.475 -191.925 49.805 -191.595 ;
        RECT 49.475 -193.285 49.805 -192.955 ;
        RECT 49.475 -194.645 49.805 -194.315 ;
        RECT 49.475 -196.005 49.805 -195.675 ;
        RECT 49.475 -197.365 49.805 -197.035 ;
        RECT 49.475 -198.725 49.805 -198.395 ;
        RECT 49.475 -200.085 49.805 -199.755 ;
        RECT 49.475 -201.445 49.805 -201.115 ;
        RECT 49.475 -202.805 49.805 -202.475 ;
        RECT 49.475 -204.165 49.805 -203.835 ;
        RECT 49.475 -205.525 49.805 -205.195 ;
        RECT 49.475 -206.885 49.805 -206.555 ;
        RECT 49.475 -208.245 49.805 -207.915 ;
        RECT 49.475 -209.605 49.805 -209.275 ;
        RECT 49.475 -210.965 49.805 -210.635 ;
        RECT 49.475 -212.325 49.805 -211.995 ;
        RECT 49.475 -213.685 49.805 -213.355 ;
        RECT 49.475 -215.045 49.805 -214.715 ;
        RECT 49.475 -216.405 49.805 -216.075 ;
        RECT 49.475 -217.765 49.805 -217.435 ;
        RECT 49.475 -219.125 49.805 -218.795 ;
        RECT 49.475 -221.37 49.805 -220.24 ;
        RECT 49.48 -221.485 49.8 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.835 129.8 51.165 130.93 ;
        RECT 50.835 127.675 51.165 128.005 ;
        RECT 50.835 126.315 51.165 126.645 ;
        RECT 50.835 124.955 51.165 125.285 ;
        RECT 50.835 123.595 51.165 123.925 ;
        RECT 50.84 123.595 51.16 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.835 -183.765 51.165 -183.435 ;
        RECT 50.835 -185.125 51.165 -184.795 ;
        RECT 50.835 -186.485 51.165 -186.155 ;
        RECT 50.835 -187.845 51.165 -187.515 ;
        RECT 50.835 -189.205 51.165 -188.875 ;
        RECT 50.835 -190.565 51.165 -190.235 ;
        RECT 50.835 -191.925 51.165 -191.595 ;
        RECT 50.835 -193.285 51.165 -192.955 ;
        RECT 50.835 -194.645 51.165 -194.315 ;
        RECT 50.835 -196.005 51.165 -195.675 ;
        RECT 50.835 -197.365 51.165 -197.035 ;
        RECT 50.835 -198.725 51.165 -198.395 ;
        RECT 50.835 -200.085 51.165 -199.755 ;
        RECT 50.835 -201.445 51.165 -201.115 ;
        RECT 50.835 -202.805 51.165 -202.475 ;
        RECT 50.835 -204.165 51.165 -203.835 ;
        RECT 50.835 -205.525 51.165 -205.195 ;
        RECT 50.835 -206.885 51.165 -206.555 ;
        RECT 50.835 -208.245 51.165 -207.915 ;
        RECT 50.835 -209.605 51.165 -209.275 ;
        RECT 50.835 -210.965 51.165 -210.635 ;
        RECT 50.835 -212.325 51.165 -211.995 ;
        RECT 50.835 -213.685 51.165 -213.355 ;
        RECT 50.835 -215.045 51.165 -214.715 ;
        RECT 50.835 -216.405 51.165 -216.075 ;
        RECT 50.835 -217.765 51.165 -217.435 ;
        RECT 50.835 -219.125 51.165 -218.795 ;
        RECT 50.835 -221.37 51.165 -220.24 ;
        RECT 50.84 -221.485 51.16 -122.235 ;
        RECT 50.835 -122.565 51.165 -122.235 ;
        RECT 50.835 -123.925 51.165 -123.595 ;
        RECT 50.835 -125.285 51.165 -124.955 ;
        RECT 50.835 -126.645 51.165 -126.315 ;
        RECT 50.835 -128.005 51.165 -127.675 ;
        RECT 50.835 -129.365 51.165 -129.035 ;
        RECT 50.835 -130.725 51.165 -130.395 ;
        RECT 50.835 -132.085 51.165 -131.755 ;
        RECT 50.835 -133.445 51.165 -133.115 ;
        RECT 50.835 -134.805 51.165 -134.475 ;
        RECT 50.835 -136.165 51.165 -135.835 ;
        RECT 50.835 -137.525 51.165 -137.195 ;
        RECT 50.835 -138.885 51.165 -138.555 ;
        RECT 50.835 -140.245 51.165 -139.915 ;
        RECT 50.835 -141.605 51.165 -141.275 ;
        RECT 50.835 -142.965 51.165 -142.635 ;
        RECT 50.835 -144.325 51.165 -143.995 ;
        RECT 50.835 -145.685 51.165 -145.355 ;
        RECT 50.835 -147.045 51.165 -146.715 ;
        RECT 50.835 -148.405 51.165 -148.075 ;
        RECT 50.835 -149.765 51.165 -149.435 ;
        RECT 50.835 -151.125 51.165 -150.795 ;
        RECT 50.835 -152.485 51.165 -152.155 ;
        RECT 50.835 -153.845 51.165 -153.515 ;
        RECT 50.835 -155.205 51.165 -154.875 ;
        RECT 50.835 -156.565 51.165 -156.235 ;
        RECT 50.835 -157.925 51.165 -157.595 ;
        RECT 50.835 -159.285 51.165 -158.955 ;
        RECT 50.835 -160.645 51.165 -160.315 ;
        RECT 50.835 -162.005 51.165 -161.675 ;
        RECT 50.835 -163.365 51.165 -163.035 ;
        RECT 50.835 -164.725 51.165 -164.395 ;
        RECT 50.835 -166.085 51.165 -165.755 ;
        RECT 50.835 -167.445 51.165 -167.115 ;
        RECT 50.835 -168.805 51.165 -168.475 ;
        RECT 50.835 -170.165 51.165 -169.835 ;
        RECT 50.835 -171.525 51.165 -171.195 ;
        RECT 50.835 -172.885 51.165 -172.555 ;
        RECT 50.835 -174.245 51.165 -173.915 ;
        RECT 50.835 -175.605 51.165 -175.275 ;
        RECT 50.835 -176.965 51.165 -176.635 ;
        RECT 50.835 -178.325 51.165 -177.995 ;
        RECT 50.835 -179.685 51.165 -179.355 ;
        RECT 50.835 -181.045 51.165 -180.715 ;
        RECT 50.835 -182.405 51.165 -182.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.515 129.8 0.845 130.93 ;
        RECT 0.515 127.675 0.845 128.005 ;
        RECT 0.515 126.315 0.845 126.645 ;
        RECT 0.515 124.955 0.845 125.285 ;
        RECT 0.515 123.595 0.845 123.925 ;
        RECT 0.52 123.595 0.84 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.515 -1.525 0.845 -1.195 ;
        RECT 0.515 -2.885 0.845 -2.555 ;
        RECT 0.52 -3.56 0.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.515 -118.485 0.845 -118.155 ;
        RECT 0.515 -119.845 0.845 -119.515 ;
        RECT 0.515 -121.205 0.845 -120.875 ;
        RECT 0.515 -122.565 0.845 -122.235 ;
        RECT 0.515 -123.925 0.845 -123.595 ;
        RECT 0.515 -125.285 0.845 -124.955 ;
        RECT 0.515 -126.645 0.845 -126.315 ;
        RECT 0.515 -128.005 0.845 -127.675 ;
        RECT 0.515 -129.365 0.845 -129.035 ;
        RECT 0.515 -130.725 0.845 -130.395 ;
        RECT 0.515 -132.085 0.845 -131.755 ;
        RECT 0.515 -133.445 0.845 -133.115 ;
        RECT 0.515 -134.805 0.845 -134.475 ;
        RECT 0.515 -136.165 0.845 -135.835 ;
        RECT 0.515 -137.525 0.845 -137.195 ;
        RECT 0.515 -138.885 0.845 -138.555 ;
        RECT 0.515 -140.245 0.845 -139.915 ;
        RECT 0.515 -141.605 0.845 -141.275 ;
        RECT 0.515 -142.965 0.845 -142.635 ;
        RECT 0.515 -144.325 0.845 -143.995 ;
        RECT 0.515 -145.685 0.845 -145.355 ;
        RECT 0.515 -147.045 0.845 -146.715 ;
        RECT 0.515 -148.405 0.845 -148.075 ;
        RECT 0.515 -149.765 0.845 -149.435 ;
        RECT 0.515 -151.125 0.845 -150.795 ;
        RECT 0.515 -152.485 0.845 -152.155 ;
        RECT 0.515 -153.845 0.845 -153.515 ;
        RECT 0.515 -155.205 0.845 -154.875 ;
        RECT 0.515 -156.565 0.845 -156.235 ;
        RECT 0.515 -157.925 0.845 -157.595 ;
        RECT 0.515 -159.285 0.845 -158.955 ;
        RECT 0.515 -160.645 0.845 -160.315 ;
        RECT 0.515 -162.005 0.845 -161.675 ;
        RECT 0.515 -163.365 0.845 -163.035 ;
        RECT 0.515 -164.725 0.845 -164.395 ;
        RECT 0.515 -166.085 0.845 -165.755 ;
        RECT 0.515 -167.445 0.845 -167.115 ;
        RECT 0.515 -168.805 0.845 -168.475 ;
        RECT 0.515 -170.165 0.845 -169.835 ;
        RECT 0.515 -171.525 0.845 -171.195 ;
        RECT 0.515 -172.885 0.845 -172.555 ;
        RECT 0.515 -174.245 0.845 -173.915 ;
        RECT 0.515 -175.605 0.845 -175.275 ;
        RECT 0.515 -176.965 0.845 -176.635 ;
        RECT 0.515 -178.325 0.845 -177.995 ;
        RECT 0.515 -179.685 0.845 -179.355 ;
        RECT 0.515 -181.045 0.845 -180.715 ;
        RECT 0.515 -182.405 0.845 -182.075 ;
        RECT 0.515 -183.765 0.845 -183.435 ;
        RECT 0.515 -185.125 0.845 -184.795 ;
        RECT 0.515 -186.485 0.845 -186.155 ;
        RECT 0.515 -187.845 0.845 -187.515 ;
        RECT 0.515 -189.205 0.845 -188.875 ;
        RECT 0.515 -190.565 0.845 -190.235 ;
        RECT 0.515 -191.925 0.845 -191.595 ;
        RECT 0.515 -193.285 0.845 -192.955 ;
        RECT 0.515 -194.645 0.845 -194.315 ;
        RECT 0.515 -196.005 0.845 -195.675 ;
        RECT 0.515 -197.365 0.845 -197.035 ;
        RECT 0.515 -198.725 0.845 -198.395 ;
        RECT 0.515 -200.085 0.845 -199.755 ;
        RECT 0.515 -201.445 0.845 -201.115 ;
        RECT 0.515 -202.805 0.845 -202.475 ;
        RECT 0.515 -204.165 0.845 -203.835 ;
        RECT 0.515 -205.525 0.845 -205.195 ;
        RECT 0.515 -206.885 0.845 -206.555 ;
        RECT 0.515 -208.245 0.845 -207.915 ;
        RECT 0.515 -209.605 0.845 -209.275 ;
        RECT 0.515 -210.965 0.845 -210.635 ;
        RECT 0.515 -212.325 0.845 -211.995 ;
        RECT 0.515 -213.685 0.845 -213.355 ;
        RECT 0.515 -215.045 0.845 -214.715 ;
        RECT 0.515 -216.405 0.845 -216.075 ;
        RECT 0.515 -217.765 0.845 -217.435 ;
        RECT 0.515 -219.125 0.845 -218.795 ;
        RECT 0.515 -221.37 0.845 -220.24 ;
        RECT 0.52 -221.485 0.84 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.875 129.8 2.205 130.93 ;
        RECT 1.875 127.675 2.205 128.005 ;
        RECT 1.875 126.315 2.205 126.645 ;
        RECT 1.875 124.955 2.205 125.285 ;
        RECT 1.875 123.595 2.205 123.925 ;
        RECT 1.88 123.595 2.2 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.875 -1.525 2.205 -1.195 ;
        RECT 1.875 -2.885 2.205 -2.555 ;
        RECT 1.88 -3.56 2.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.875 -118.485 2.205 -118.155 ;
        RECT 1.875 -119.845 2.205 -119.515 ;
        RECT 1.875 -121.205 2.205 -120.875 ;
        RECT 1.875 -122.565 2.205 -122.235 ;
        RECT 1.875 -123.925 2.205 -123.595 ;
        RECT 1.875 -125.285 2.205 -124.955 ;
        RECT 1.875 -126.645 2.205 -126.315 ;
        RECT 1.875 -128.005 2.205 -127.675 ;
        RECT 1.875 -129.365 2.205 -129.035 ;
        RECT 1.875 -130.725 2.205 -130.395 ;
        RECT 1.875 -132.085 2.205 -131.755 ;
        RECT 1.875 -133.445 2.205 -133.115 ;
        RECT 1.875 -134.805 2.205 -134.475 ;
        RECT 1.875 -136.165 2.205 -135.835 ;
        RECT 1.875 -137.525 2.205 -137.195 ;
        RECT 1.875 -138.885 2.205 -138.555 ;
        RECT 1.875 -140.245 2.205 -139.915 ;
        RECT 1.875 -141.605 2.205 -141.275 ;
        RECT 1.875 -142.965 2.205 -142.635 ;
        RECT 1.875 -144.325 2.205 -143.995 ;
        RECT 1.875 -145.685 2.205 -145.355 ;
        RECT 1.875 -147.045 2.205 -146.715 ;
        RECT 1.875 -148.405 2.205 -148.075 ;
        RECT 1.875 -149.765 2.205 -149.435 ;
        RECT 1.875 -151.125 2.205 -150.795 ;
        RECT 1.875 -152.485 2.205 -152.155 ;
        RECT 1.875 -153.845 2.205 -153.515 ;
        RECT 1.875 -155.205 2.205 -154.875 ;
        RECT 1.875 -156.565 2.205 -156.235 ;
        RECT 1.875 -157.925 2.205 -157.595 ;
        RECT 1.875 -159.285 2.205 -158.955 ;
        RECT 1.875 -160.645 2.205 -160.315 ;
        RECT 1.875 -162.005 2.205 -161.675 ;
        RECT 1.875 -163.365 2.205 -163.035 ;
        RECT 1.875 -164.725 2.205 -164.395 ;
        RECT 1.875 -166.085 2.205 -165.755 ;
        RECT 1.875 -167.445 2.205 -167.115 ;
        RECT 1.875 -168.805 2.205 -168.475 ;
        RECT 1.875 -170.165 2.205 -169.835 ;
        RECT 1.875 -171.525 2.205 -171.195 ;
        RECT 1.875 -172.885 2.205 -172.555 ;
        RECT 1.875 -174.245 2.205 -173.915 ;
        RECT 1.875 -175.605 2.205 -175.275 ;
        RECT 1.875 -176.965 2.205 -176.635 ;
        RECT 1.875 -178.325 2.205 -177.995 ;
        RECT 1.875 -179.685 2.205 -179.355 ;
        RECT 1.875 -181.045 2.205 -180.715 ;
        RECT 1.875 -182.405 2.205 -182.075 ;
        RECT 1.875 -183.765 2.205 -183.435 ;
        RECT 1.875 -185.125 2.205 -184.795 ;
        RECT 1.875 -186.485 2.205 -186.155 ;
        RECT 1.875 -187.845 2.205 -187.515 ;
        RECT 1.875 -189.205 2.205 -188.875 ;
        RECT 1.875 -190.565 2.205 -190.235 ;
        RECT 1.875 -191.925 2.205 -191.595 ;
        RECT 1.875 -193.285 2.205 -192.955 ;
        RECT 1.875 -194.645 2.205 -194.315 ;
        RECT 1.875 -196.005 2.205 -195.675 ;
        RECT 1.875 -197.365 2.205 -197.035 ;
        RECT 1.875 -198.725 2.205 -198.395 ;
        RECT 1.875 -200.085 2.205 -199.755 ;
        RECT 1.875 -201.445 2.205 -201.115 ;
        RECT 1.875 -202.805 2.205 -202.475 ;
        RECT 1.875 -204.165 2.205 -203.835 ;
        RECT 1.875 -205.525 2.205 -205.195 ;
        RECT 1.875 -206.885 2.205 -206.555 ;
        RECT 1.875 -208.245 2.205 -207.915 ;
        RECT 1.875 -209.605 2.205 -209.275 ;
        RECT 1.875 -210.965 2.205 -210.635 ;
        RECT 1.875 -212.325 2.205 -211.995 ;
        RECT 1.875 -213.685 2.205 -213.355 ;
        RECT 1.875 -215.045 2.205 -214.715 ;
        RECT 1.875 -216.405 2.205 -216.075 ;
        RECT 1.875 -217.765 2.205 -217.435 ;
        RECT 1.875 -219.125 2.205 -218.795 ;
        RECT 1.875 -221.37 2.205 -220.24 ;
        RECT 1.88 -221.485 2.2 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.235 129.8 3.565 130.93 ;
        RECT 3.235 127.675 3.565 128.005 ;
        RECT 3.235 126.315 3.565 126.645 ;
        RECT 3.235 124.955 3.565 125.285 ;
        RECT 3.235 123.595 3.565 123.925 ;
        RECT 3.24 123.595 3.56 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.235 -122.565 3.565 -122.235 ;
        RECT 3.235 -123.925 3.565 -123.595 ;
        RECT 3.235 -125.285 3.565 -124.955 ;
        RECT 3.235 -126.645 3.565 -126.315 ;
        RECT 3.235 -128.005 3.565 -127.675 ;
        RECT 3.235 -129.365 3.565 -129.035 ;
        RECT 3.235 -130.725 3.565 -130.395 ;
        RECT 3.235 -132.085 3.565 -131.755 ;
        RECT 3.235 -133.445 3.565 -133.115 ;
        RECT 3.235 -134.805 3.565 -134.475 ;
        RECT 3.235 -136.165 3.565 -135.835 ;
        RECT 3.235 -137.525 3.565 -137.195 ;
        RECT 3.235 -138.885 3.565 -138.555 ;
        RECT 3.235 -140.245 3.565 -139.915 ;
        RECT 3.235 -141.605 3.565 -141.275 ;
        RECT 3.235 -142.965 3.565 -142.635 ;
        RECT 3.235 -144.325 3.565 -143.995 ;
        RECT 3.235 -145.685 3.565 -145.355 ;
        RECT 3.235 -147.045 3.565 -146.715 ;
        RECT 3.235 -148.405 3.565 -148.075 ;
        RECT 3.235 -149.765 3.565 -149.435 ;
        RECT 3.235 -151.125 3.565 -150.795 ;
        RECT 3.235 -152.485 3.565 -152.155 ;
        RECT 3.235 -153.845 3.565 -153.515 ;
        RECT 3.235 -155.205 3.565 -154.875 ;
        RECT 3.235 -156.565 3.565 -156.235 ;
        RECT 3.235 -157.925 3.565 -157.595 ;
        RECT 3.235 -159.285 3.565 -158.955 ;
        RECT 3.235 -160.645 3.565 -160.315 ;
        RECT 3.235 -162.005 3.565 -161.675 ;
        RECT 3.235 -163.365 3.565 -163.035 ;
        RECT 3.235 -164.725 3.565 -164.395 ;
        RECT 3.235 -166.085 3.565 -165.755 ;
        RECT 3.235 -167.445 3.565 -167.115 ;
        RECT 3.235 -168.805 3.565 -168.475 ;
        RECT 3.235 -170.165 3.565 -169.835 ;
        RECT 3.235 -171.525 3.565 -171.195 ;
        RECT 3.235 -172.885 3.565 -172.555 ;
        RECT 3.235 -174.245 3.565 -173.915 ;
        RECT 3.235 -175.605 3.565 -175.275 ;
        RECT 3.235 -176.965 3.565 -176.635 ;
        RECT 3.235 -178.325 3.565 -177.995 ;
        RECT 3.235 -179.685 3.565 -179.355 ;
        RECT 3.235 -181.045 3.565 -180.715 ;
        RECT 3.235 -182.405 3.565 -182.075 ;
        RECT 3.235 -183.765 3.565 -183.435 ;
        RECT 3.235 -185.125 3.565 -184.795 ;
        RECT 3.235 -186.485 3.565 -186.155 ;
        RECT 3.235 -187.845 3.565 -187.515 ;
        RECT 3.235 -189.205 3.565 -188.875 ;
        RECT 3.235 -190.565 3.565 -190.235 ;
        RECT 3.235 -191.925 3.565 -191.595 ;
        RECT 3.235 -193.285 3.565 -192.955 ;
        RECT 3.235 -194.645 3.565 -194.315 ;
        RECT 3.235 -196.005 3.565 -195.675 ;
        RECT 3.235 -197.365 3.565 -197.035 ;
        RECT 3.235 -198.725 3.565 -198.395 ;
        RECT 3.235 -200.085 3.565 -199.755 ;
        RECT 3.235 -201.445 3.565 -201.115 ;
        RECT 3.235 -202.805 3.565 -202.475 ;
        RECT 3.235 -204.165 3.565 -203.835 ;
        RECT 3.235 -205.525 3.565 -205.195 ;
        RECT 3.235 -206.885 3.565 -206.555 ;
        RECT 3.235 -208.245 3.565 -207.915 ;
        RECT 3.235 -209.605 3.565 -209.275 ;
        RECT 3.235 -210.965 3.565 -210.635 ;
        RECT 3.235 -212.325 3.565 -211.995 ;
        RECT 3.235 -213.685 3.565 -213.355 ;
        RECT 3.235 -215.045 3.565 -214.715 ;
        RECT 3.235 -216.405 3.565 -216.075 ;
        RECT 3.235 -217.765 3.565 -217.435 ;
        RECT 3.235 -219.125 3.565 -218.795 ;
        RECT 3.235 -221.37 3.565 -220.24 ;
        RECT 3.24 -221.485 3.56 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.31 -121.535 3.64 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.595 129.8 4.925 130.93 ;
        RECT 4.595 127.675 4.925 128.005 ;
        RECT 4.595 126.315 4.925 126.645 ;
        RECT 4.595 124.955 4.925 125.285 ;
        RECT 4.595 123.595 4.925 123.925 ;
        RECT 4.6 123.595 4.92 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.595 -1.525 4.925 -1.195 ;
        RECT 4.595 -2.885 4.925 -2.555 ;
        RECT 4.6 -3.56 4.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.955 129.8 6.285 130.93 ;
        RECT 5.955 127.675 6.285 128.005 ;
        RECT 5.955 126.315 6.285 126.645 ;
        RECT 5.955 124.955 6.285 125.285 ;
        RECT 5.955 123.595 6.285 123.925 ;
        RECT 5.96 123.595 6.28 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.955 -1.525 6.285 -1.195 ;
        RECT 5.955 -2.885 6.285 -2.555 ;
        RECT 5.96 -3.56 6.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.315 129.8 7.645 130.93 ;
        RECT 7.315 127.675 7.645 128.005 ;
        RECT 7.315 126.315 7.645 126.645 ;
        RECT 7.315 124.955 7.645 125.285 ;
        RECT 7.315 123.595 7.645 123.925 ;
        RECT 7.32 123.595 7.64 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.315 -1.525 7.645 -1.195 ;
        RECT 7.315 -2.885 7.645 -2.555 ;
        RECT 7.32 -3.56 7.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.315 -118.485 7.645 -118.155 ;
        RECT 7.315 -119.845 7.645 -119.515 ;
        RECT 7.315 -121.205 7.645 -120.875 ;
        RECT 7.315 -122.565 7.645 -122.235 ;
        RECT 7.315 -123.925 7.645 -123.595 ;
        RECT 7.315 -125.285 7.645 -124.955 ;
        RECT 7.315 -126.645 7.645 -126.315 ;
        RECT 7.315 -128.005 7.645 -127.675 ;
        RECT 7.315 -129.365 7.645 -129.035 ;
        RECT 7.315 -130.725 7.645 -130.395 ;
        RECT 7.315 -132.085 7.645 -131.755 ;
        RECT 7.315 -133.445 7.645 -133.115 ;
        RECT 7.315 -134.805 7.645 -134.475 ;
        RECT 7.315 -136.165 7.645 -135.835 ;
        RECT 7.315 -137.525 7.645 -137.195 ;
        RECT 7.315 -138.885 7.645 -138.555 ;
        RECT 7.315 -140.245 7.645 -139.915 ;
        RECT 7.315 -141.605 7.645 -141.275 ;
        RECT 7.315 -142.965 7.645 -142.635 ;
        RECT 7.315 -144.325 7.645 -143.995 ;
        RECT 7.315 -145.685 7.645 -145.355 ;
        RECT 7.315 -147.045 7.645 -146.715 ;
        RECT 7.315 -148.405 7.645 -148.075 ;
        RECT 7.315 -149.765 7.645 -149.435 ;
        RECT 7.315 -151.125 7.645 -150.795 ;
        RECT 7.315 -152.485 7.645 -152.155 ;
        RECT 7.315 -153.845 7.645 -153.515 ;
        RECT 7.315 -155.205 7.645 -154.875 ;
        RECT 7.315 -156.565 7.645 -156.235 ;
        RECT 7.315 -157.925 7.645 -157.595 ;
        RECT 7.315 -159.285 7.645 -158.955 ;
        RECT 7.315 -160.645 7.645 -160.315 ;
        RECT 7.315 -162.005 7.645 -161.675 ;
        RECT 7.315 -163.365 7.645 -163.035 ;
        RECT 7.315 -164.725 7.645 -164.395 ;
        RECT 7.315 -166.085 7.645 -165.755 ;
        RECT 7.315 -167.445 7.645 -167.115 ;
        RECT 7.315 -168.805 7.645 -168.475 ;
        RECT 7.315 -170.165 7.645 -169.835 ;
        RECT 7.315 -171.525 7.645 -171.195 ;
        RECT 7.315 -172.885 7.645 -172.555 ;
        RECT 7.315 -174.245 7.645 -173.915 ;
        RECT 7.315 -175.605 7.645 -175.275 ;
        RECT 7.315 -176.965 7.645 -176.635 ;
        RECT 7.315 -178.325 7.645 -177.995 ;
        RECT 7.315 -179.685 7.645 -179.355 ;
        RECT 7.315 -181.045 7.645 -180.715 ;
        RECT 7.315 -182.405 7.645 -182.075 ;
        RECT 7.315 -183.765 7.645 -183.435 ;
        RECT 7.315 -185.125 7.645 -184.795 ;
        RECT 7.315 -186.485 7.645 -186.155 ;
        RECT 7.315 -187.845 7.645 -187.515 ;
        RECT 7.315 -189.205 7.645 -188.875 ;
        RECT 7.315 -190.565 7.645 -190.235 ;
        RECT 7.315 -191.925 7.645 -191.595 ;
        RECT 7.315 -193.285 7.645 -192.955 ;
        RECT 7.315 -194.645 7.645 -194.315 ;
        RECT 7.315 -196.005 7.645 -195.675 ;
        RECT 7.315 -197.365 7.645 -197.035 ;
        RECT 7.315 -198.725 7.645 -198.395 ;
        RECT 7.315 -200.085 7.645 -199.755 ;
        RECT 7.315 -201.445 7.645 -201.115 ;
        RECT 7.315 -202.805 7.645 -202.475 ;
        RECT 7.315 -204.165 7.645 -203.835 ;
        RECT 7.315 -205.525 7.645 -205.195 ;
        RECT 7.315 -206.885 7.645 -206.555 ;
        RECT 7.315 -208.245 7.645 -207.915 ;
        RECT 7.315 -209.605 7.645 -209.275 ;
        RECT 7.315 -210.965 7.645 -210.635 ;
        RECT 7.315 -212.325 7.645 -211.995 ;
        RECT 7.315 -213.685 7.645 -213.355 ;
        RECT 7.315 -215.045 7.645 -214.715 ;
        RECT 7.315 -216.405 7.645 -216.075 ;
        RECT 7.315 -217.765 7.645 -217.435 ;
        RECT 7.315 -219.125 7.645 -218.795 ;
        RECT 7.315 -221.37 7.645 -220.24 ;
        RECT 7.32 -221.485 7.64 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.675 129.8 9.005 130.93 ;
        RECT 8.675 127.675 9.005 128.005 ;
        RECT 8.675 126.315 9.005 126.645 ;
        RECT 8.675 124.955 9.005 125.285 ;
        RECT 8.675 123.595 9.005 123.925 ;
        RECT 8.68 123.595 9 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.675 -122.565 9.005 -122.235 ;
        RECT 8.675 -123.925 9.005 -123.595 ;
        RECT 8.675 -125.285 9.005 -124.955 ;
        RECT 8.675 -126.645 9.005 -126.315 ;
        RECT 8.675 -128.005 9.005 -127.675 ;
        RECT 8.675 -129.365 9.005 -129.035 ;
        RECT 8.675 -130.725 9.005 -130.395 ;
        RECT 8.675 -132.085 9.005 -131.755 ;
        RECT 8.675 -133.445 9.005 -133.115 ;
        RECT 8.675 -134.805 9.005 -134.475 ;
        RECT 8.675 -136.165 9.005 -135.835 ;
        RECT 8.675 -137.525 9.005 -137.195 ;
        RECT 8.675 -138.885 9.005 -138.555 ;
        RECT 8.675 -140.245 9.005 -139.915 ;
        RECT 8.675 -141.605 9.005 -141.275 ;
        RECT 8.675 -142.965 9.005 -142.635 ;
        RECT 8.675 -144.325 9.005 -143.995 ;
        RECT 8.675 -145.685 9.005 -145.355 ;
        RECT 8.675 -147.045 9.005 -146.715 ;
        RECT 8.675 -148.405 9.005 -148.075 ;
        RECT 8.675 -149.765 9.005 -149.435 ;
        RECT 8.675 -151.125 9.005 -150.795 ;
        RECT 8.675 -152.485 9.005 -152.155 ;
        RECT 8.675 -153.845 9.005 -153.515 ;
        RECT 8.675 -155.205 9.005 -154.875 ;
        RECT 8.675 -156.565 9.005 -156.235 ;
        RECT 8.675 -157.925 9.005 -157.595 ;
        RECT 8.675 -159.285 9.005 -158.955 ;
        RECT 8.675 -160.645 9.005 -160.315 ;
        RECT 8.675 -162.005 9.005 -161.675 ;
        RECT 8.675 -163.365 9.005 -163.035 ;
        RECT 8.675 -164.725 9.005 -164.395 ;
        RECT 8.675 -166.085 9.005 -165.755 ;
        RECT 8.675 -167.445 9.005 -167.115 ;
        RECT 8.675 -168.805 9.005 -168.475 ;
        RECT 8.675 -170.165 9.005 -169.835 ;
        RECT 8.675 -171.525 9.005 -171.195 ;
        RECT 8.675 -172.885 9.005 -172.555 ;
        RECT 8.675 -174.245 9.005 -173.915 ;
        RECT 8.675 -175.605 9.005 -175.275 ;
        RECT 8.675 -176.965 9.005 -176.635 ;
        RECT 8.675 -178.325 9.005 -177.995 ;
        RECT 8.675 -179.685 9.005 -179.355 ;
        RECT 8.675 -181.045 9.005 -180.715 ;
        RECT 8.675 -182.405 9.005 -182.075 ;
        RECT 8.675 -183.765 9.005 -183.435 ;
        RECT 8.675 -185.125 9.005 -184.795 ;
        RECT 8.675 -186.485 9.005 -186.155 ;
        RECT 8.675 -187.845 9.005 -187.515 ;
        RECT 8.675 -189.205 9.005 -188.875 ;
        RECT 8.675 -190.565 9.005 -190.235 ;
        RECT 8.675 -191.925 9.005 -191.595 ;
        RECT 8.675 -193.285 9.005 -192.955 ;
        RECT 8.675 -194.645 9.005 -194.315 ;
        RECT 8.675 -196.005 9.005 -195.675 ;
        RECT 8.675 -197.365 9.005 -197.035 ;
        RECT 8.675 -198.725 9.005 -198.395 ;
        RECT 8.675 -200.085 9.005 -199.755 ;
        RECT 8.675 -201.445 9.005 -201.115 ;
        RECT 8.675 -202.805 9.005 -202.475 ;
        RECT 8.675 -204.165 9.005 -203.835 ;
        RECT 8.675 -205.525 9.005 -205.195 ;
        RECT 8.675 -206.885 9.005 -206.555 ;
        RECT 8.675 -208.245 9.005 -207.915 ;
        RECT 8.675 -209.605 9.005 -209.275 ;
        RECT 8.675 -210.965 9.005 -210.635 ;
        RECT 8.675 -212.325 9.005 -211.995 ;
        RECT 8.675 -213.685 9.005 -213.355 ;
        RECT 8.675 -215.045 9.005 -214.715 ;
        RECT 8.675 -216.405 9.005 -216.075 ;
        RECT 8.675 -217.765 9.005 -217.435 ;
        RECT 8.675 -219.125 9.005 -218.795 ;
        RECT 8.675 -221.37 9.005 -220.24 ;
        RECT 8.68 -221.485 9 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.41 -121.535 9.74 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.035 129.8 10.365 130.93 ;
        RECT 10.035 127.675 10.365 128.005 ;
        RECT 10.035 126.315 10.365 126.645 ;
        RECT 10.035 124.955 10.365 125.285 ;
        RECT 10.035 123.595 10.365 123.925 ;
        RECT 10.04 123.595 10.36 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.395 129.8 11.725 130.93 ;
        RECT 11.395 127.675 11.725 128.005 ;
        RECT 11.395 126.315 11.725 126.645 ;
        RECT 11.395 124.955 11.725 125.285 ;
        RECT 11.395 123.595 11.725 123.925 ;
        RECT 11.4 123.595 11.72 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.395 -1.525 11.725 -1.195 ;
        RECT 11.395 -2.885 11.725 -2.555 ;
        RECT 11.4 -3.56 11.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.755 129.8 13.085 130.93 ;
        RECT 12.755 127.675 13.085 128.005 ;
        RECT 12.755 126.315 13.085 126.645 ;
        RECT 12.755 124.955 13.085 125.285 ;
        RECT 12.755 123.595 13.085 123.925 ;
        RECT 12.76 123.595 13.08 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.755 -1.525 13.085 -1.195 ;
        RECT 12.755 -2.885 13.085 -2.555 ;
        RECT 12.76 -3.56 13.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.755 -118.485 13.085 -118.155 ;
        RECT 12.755 -119.845 13.085 -119.515 ;
        RECT 12.755 -121.205 13.085 -120.875 ;
        RECT 12.755 -122.565 13.085 -122.235 ;
        RECT 12.755 -123.925 13.085 -123.595 ;
        RECT 12.755 -125.285 13.085 -124.955 ;
        RECT 12.755 -126.645 13.085 -126.315 ;
        RECT 12.755 -128.005 13.085 -127.675 ;
        RECT 12.755 -129.365 13.085 -129.035 ;
        RECT 12.755 -130.725 13.085 -130.395 ;
        RECT 12.755 -132.085 13.085 -131.755 ;
        RECT 12.755 -133.445 13.085 -133.115 ;
        RECT 12.755 -134.805 13.085 -134.475 ;
        RECT 12.755 -136.165 13.085 -135.835 ;
        RECT 12.755 -137.525 13.085 -137.195 ;
        RECT 12.755 -138.885 13.085 -138.555 ;
        RECT 12.755 -140.245 13.085 -139.915 ;
        RECT 12.755 -141.605 13.085 -141.275 ;
        RECT 12.755 -142.965 13.085 -142.635 ;
        RECT 12.755 -144.325 13.085 -143.995 ;
        RECT 12.755 -145.685 13.085 -145.355 ;
        RECT 12.755 -147.045 13.085 -146.715 ;
        RECT 12.755 -148.405 13.085 -148.075 ;
        RECT 12.755 -149.765 13.085 -149.435 ;
        RECT 12.755 -151.125 13.085 -150.795 ;
        RECT 12.755 -152.485 13.085 -152.155 ;
        RECT 12.755 -153.845 13.085 -153.515 ;
        RECT 12.755 -155.205 13.085 -154.875 ;
        RECT 12.755 -156.565 13.085 -156.235 ;
        RECT 12.755 -157.925 13.085 -157.595 ;
        RECT 12.755 -159.285 13.085 -158.955 ;
        RECT 12.755 -160.645 13.085 -160.315 ;
        RECT 12.755 -162.005 13.085 -161.675 ;
        RECT 12.755 -163.365 13.085 -163.035 ;
        RECT 12.755 -164.725 13.085 -164.395 ;
        RECT 12.755 -166.085 13.085 -165.755 ;
        RECT 12.755 -167.445 13.085 -167.115 ;
        RECT 12.755 -168.805 13.085 -168.475 ;
        RECT 12.755 -170.165 13.085 -169.835 ;
        RECT 12.755 -171.525 13.085 -171.195 ;
        RECT 12.755 -172.885 13.085 -172.555 ;
        RECT 12.755 -174.245 13.085 -173.915 ;
        RECT 12.755 -175.605 13.085 -175.275 ;
        RECT 12.755 -176.965 13.085 -176.635 ;
        RECT 12.755 -178.325 13.085 -177.995 ;
        RECT 12.755 -179.685 13.085 -179.355 ;
        RECT 12.755 -181.045 13.085 -180.715 ;
        RECT 12.755 -182.405 13.085 -182.075 ;
        RECT 12.755 -183.765 13.085 -183.435 ;
        RECT 12.755 -185.125 13.085 -184.795 ;
        RECT 12.755 -186.485 13.085 -186.155 ;
        RECT 12.755 -187.845 13.085 -187.515 ;
        RECT 12.755 -189.205 13.085 -188.875 ;
        RECT 12.755 -190.565 13.085 -190.235 ;
        RECT 12.755 -191.925 13.085 -191.595 ;
        RECT 12.755 -193.285 13.085 -192.955 ;
        RECT 12.755 -194.645 13.085 -194.315 ;
        RECT 12.755 -196.005 13.085 -195.675 ;
        RECT 12.755 -197.365 13.085 -197.035 ;
        RECT 12.755 -198.725 13.085 -198.395 ;
        RECT 12.755 -200.085 13.085 -199.755 ;
        RECT 12.755 -201.445 13.085 -201.115 ;
        RECT 12.755 -202.805 13.085 -202.475 ;
        RECT 12.755 -204.165 13.085 -203.835 ;
        RECT 12.755 -205.525 13.085 -205.195 ;
        RECT 12.755 -206.885 13.085 -206.555 ;
        RECT 12.755 -208.245 13.085 -207.915 ;
        RECT 12.755 -209.605 13.085 -209.275 ;
        RECT 12.755 -210.965 13.085 -210.635 ;
        RECT 12.755 -212.325 13.085 -211.995 ;
        RECT 12.755 -213.685 13.085 -213.355 ;
        RECT 12.755 -215.045 13.085 -214.715 ;
        RECT 12.755 -216.405 13.085 -216.075 ;
        RECT 12.755 -217.765 13.085 -217.435 ;
        RECT 12.755 -219.125 13.085 -218.795 ;
        RECT 12.755 -221.37 13.085 -220.24 ;
        RECT 12.76 -221.485 13.08 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.115 129.8 14.445 130.93 ;
        RECT 14.115 127.675 14.445 128.005 ;
        RECT 14.115 126.315 14.445 126.645 ;
        RECT 14.115 124.955 14.445 125.285 ;
        RECT 14.115 123.595 14.445 123.925 ;
        RECT 14.12 123.595 14.44 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.115 -1.525 14.445 -1.195 ;
        RECT 14.115 -2.885 14.445 -2.555 ;
        RECT 14.12 -3.56 14.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.115 -118.485 14.445 -118.155 ;
        RECT 14.115 -119.845 14.445 -119.515 ;
        RECT 14.115 -121.205 14.445 -120.875 ;
        RECT 14.115 -122.565 14.445 -122.235 ;
        RECT 14.115 -123.925 14.445 -123.595 ;
        RECT 14.115 -125.285 14.445 -124.955 ;
        RECT 14.115 -126.645 14.445 -126.315 ;
        RECT 14.115 -128.005 14.445 -127.675 ;
        RECT 14.115 -129.365 14.445 -129.035 ;
        RECT 14.115 -130.725 14.445 -130.395 ;
        RECT 14.115 -132.085 14.445 -131.755 ;
        RECT 14.115 -133.445 14.445 -133.115 ;
        RECT 14.115 -134.805 14.445 -134.475 ;
        RECT 14.115 -136.165 14.445 -135.835 ;
        RECT 14.115 -137.525 14.445 -137.195 ;
        RECT 14.115 -138.885 14.445 -138.555 ;
        RECT 14.115 -140.245 14.445 -139.915 ;
        RECT 14.115 -141.605 14.445 -141.275 ;
        RECT 14.115 -142.965 14.445 -142.635 ;
        RECT 14.115 -144.325 14.445 -143.995 ;
        RECT 14.115 -145.685 14.445 -145.355 ;
        RECT 14.115 -147.045 14.445 -146.715 ;
        RECT 14.115 -148.405 14.445 -148.075 ;
        RECT 14.115 -149.765 14.445 -149.435 ;
        RECT 14.115 -151.125 14.445 -150.795 ;
        RECT 14.115 -152.485 14.445 -152.155 ;
        RECT 14.115 -153.845 14.445 -153.515 ;
        RECT 14.115 -155.205 14.445 -154.875 ;
        RECT 14.115 -156.565 14.445 -156.235 ;
        RECT 14.115 -157.925 14.445 -157.595 ;
        RECT 14.115 -159.285 14.445 -158.955 ;
        RECT 14.115 -160.645 14.445 -160.315 ;
        RECT 14.115 -162.005 14.445 -161.675 ;
        RECT 14.115 -163.365 14.445 -163.035 ;
        RECT 14.115 -164.725 14.445 -164.395 ;
        RECT 14.115 -166.085 14.445 -165.755 ;
        RECT 14.115 -167.445 14.445 -167.115 ;
        RECT 14.115 -168.805 14.445 -168.475 ;
        RECT 14.115 -170.165 14.445 -169.835 ;
        RECT 14.115 -171.525 14.445 -171.195 ;
        RECT 14.115 -172.885 14.445 -172.555 ;
        RECT 14.115 -174.245 14.445 -173.915 ;
        RECT 14.115 -175.605 14.445 -175.275 ;
        RECT 14.115 -176.965 14.445 -176.635 ;
        RECT 14.115 -178.325 14.445 -177.995 ;
        RECT 14.115 -179.685 14.445 -179.355 ;
        RECT 14.115 -181.045 14.445 -180.715 ;
        RECT 14.115 -182.405 14.445 -182.075 ;
        RECT 14.115 -183.765 14.445 -183.435 ;
        RECT 14.115 -185.125 14.445 -184.795 ;
        RECT 14.115 -186.485 14.445 -186.155 ;
        RECT 14.115 -187.845 14.445 -187.515 ;
        RECT 14.115 -189.205 14.445 -188.875 ;
        RECT 14.115 -190.565 14.445 -190.235 ;
        RECT 14.115 -191.925 14.445 -191.595 ;
        RECT 14.115 -193.285 14.445 -192.955 ;
        RECT 14.115 -194.645 14.445 -194.315 ;
        RECT 14.115 -196.005 14.445 -195.675 ;
        RECT 14.115 -197.365 14.445 -197.035 ;
        RECT 14.115 -198.725 14.445 -198.395 ;
        RECT 14.115 -200.085 14.445 -199.755 ;
        RECT 14.115 -201.445 14.445 -201.115 ;
        RECT 14.115 -202.805 14.445 -202.475 ;
        RECT 14.115 -204.165 14.445 -203.835 ;
        RECT 14.115 -205.525 14.445 -205.195 ;
        RECT 14.115 -206.885 14.445 -206.555 ;
        RECT 14.115 -208.245 14.445 -207.915 ;
        RECT 14.115 -209.605 14.445 -209.275 ;
        RECT 14.115 -210.965 14.445 -210.635 ;
        RECT 14.115 -212.325 14.445 -211.995 ;
        RECT 14.115 -213.685 14.445 -213.355 ;
        RECT 14.115 -215.045 14.445 -214.715 ;
        RECT 14.115 -216.405 14.445 -216.075 ;
        RECT 14.115 -217.765 14.445 -217.435 ;
        RECT 14.115 -219.125 14.445 -218.795 ;
        RECT 14.115 -221.37 14.445 -220.24 ;
        RECT 14.12 -221.485 14.44 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.475 129.8 15.805 130.93 ;
        RECT 15.475 127.675 15.805 128.005 ;
        RECT 15.475 126.315 15.805 126.645 ;
        RECT 15.475 124.955 15.805 125.285 ;
        RECT 15.475 123.595 15.805 123.925 ;
        RECT 15.48 123.595 15.8 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.475 -122.565 15.805 -122.235 ;
        RECT 15.475 -123.925 15.805 -123.595 ;
        RECT 15.475 -125.285 15.805 -124.955 ;
        RECT 15.475 -126.645 15.805 -126.315 ;
        RECT 15.475 -128.005 15.805 -127.675 ;
        RECT 15.475 -129.365 15.805 -129.035 ;
        RECT 15.475 -130.725 15.805 -130.395 ;
        RECT 15.475 -132.085 15.805 -131.755 ;
        RECT 15.475 -133.445 15.805 -133.115 ;
        RECT 15.475 -134.805 15.805 -134.475 ;
        RECT 15.475 -136.165 15.805 -135.835 ;
        RECT 15.475 -137.525 15.805 -137.195 ;
        RECT 15.475 -138.885 15.805 -138.555 ;
        RECT 15.475 -140.245 15.805 -139.915 ;
        RECT 15.475 -141.605 15.805 -141.275 ;
        RECT 15.475 -142.965 15.805 -142.635 ;
        RECT 15.475 -144.325 15.805 -143.995 ;
        RECT 15.475 -145.685 15.805 -145.355 ;
        RECT 15.475 -147.045 15.805 -146.715 ;
        RECT 15.475 -148.405 15.805 -148.075 ;
        RECT 15.475 -149.765 15.805 -149.435 ;
        RECT 15.475 -151.125 15.805 -150.795 ;
        RECT 15.475 -152.485 15.805 -152.155 ;
        RECT 15.475 -153.845 15.805 -153.515 ;
        RECT 15.475 -155.205 15.805 -154.875 ;
        RECT 15.475 -156.565 15.805 -156.235 ;
        RECT 15.475 -157.925 15.805 -157.595 ;
        RECT 15.475 -159.285 15.805 -158.955 ;
        RECT 15.475 -160.645 15.805 -160.315 ;
        RECT 15.475 -162.005 15.805 -161.675 ;
        RECT 15.475 -163.365 15.805 -163.035 ;
        RECT 15.475 -164.725 15.805 -164.395 ;
        RECT 15.475 -166.085 15.805 -165.755 ;
        RECT 15.475 -167.445 15.805 -167.115 ;
        RECT 15.475 -168.805 15.805 -168.475 ;
        RECT 15.475 -170.165 15.805 -169.835 ;
        RECT 15.475 -171.525 15.805 -171.195 ;
        RECT 15.475 -172.885 15.805 -172.555 ;
        RECT 15.475 -174.245 15.805 -173.915 ;
        RECT 15.475 -175.605 15.805 -175.275 ;
        RECT 15.475 -176.965 15.805 -176.635 ;
        RECT 15.475 -178.325 15.805 -177.995 ;
        RECT 15.475 -179.685 15.805 -179.355 ;
        RECT 15.475 -181.045 15.805 -180.715 ;
        RECT 15.475 -182.405 15.805 -182.075 ;
        RECT 15.475 -183.765 15.805 -183.435 ;
        RECT 15.475 -185.125 15.805 -184.795 ;
        RECT 15.475 -186.485 15.805 -186.155 ;
        RECT 15.475 -187.845 15.805 -187.515 ;
        RECT 15.475 -189.205 15.805 -188.875 ;
        RECT 15.475 -190.565 15.805 -190.235 ;
        RECT 15.475 -191.925 15.805 -191.595 ;
        RECT 15.475 -193.285 15.805 -192.955 ;
        RECT 15.475 -194.645 15.805 -194.315 ;
        RECT 15.475 -196.005 15.805 -195.675 ;
        RECT 15.475 -197.365 15.805 -197.035 ;
        RECT 15.475 -198.725 15.805 -198.395 ;
        RECT 15.475 -200.085 15.805 -199.755 ;
        RECT 15.475 -201.445 15.805 -201.115 ;
        RECT 15.475 -202.805 15.805 -202.475 ;
        RECT 15.475 -204.165 15.805 -203.835 ;
        RECT 15.475 -205.525 15.805 -205.195 ;
        RECT 15.475 -206.885 15.805 -206.555 ;
        RECT 15.475 -208.245 15.805 -207.915 ;
        RECT 15.475 -209.605 15.805 -209.275 ;
        RECT 15.475 -210.965 15.805 -210.635 ;
        RECT 15.475 -212.325 15.805 -211.995 ;
        RECT 15.475 -213.685 15.805 -213.355 ;
        RECT 15.475 -215.045 15.805 -214.715 ;
        RECT 15.475 -216.405 15.805 -216.075 ;
        RECT 15.475 -217.765 15.805 -217.435 ;
        RECT 15.475 -219.125 15.805 -218.795 ;
        RECT 15.475 -221.37 15.805 -220.24 ;
        RECT 15.48 -221.485 15.8 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.51 -121.535 15.84 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.835 129.8 17.165 130.93 ;
        RECT 16.835 127.675 17.165 128.005 ;
        RECT 16.835 126.315 17.165 126.645 ;
        RECT 16.835 124.955 17.165 125.285 ;
        RECT 16.835 123.595 17.165 123.925 ;
        RECT 16.84 123.595 17.16 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.835 -1.525 17.165 -1.195 ;
        RECT 16.835 -2.885 17.165 -2.555 ;
        RECT 16.84 -3.56 17.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.195 129.8 18.525 130.93 ;
        RECT 18.195 127.675 18.525 128.005 ;
        RECT 18.195 126.315 18.525 126.645 ;
        RECT 18.195 124.955 18.525 125.285 ;
        RECT 18.195 123.595 18.525 123.925 ;
        RECT 18.2 123.595 18.52 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.195 -1.525 18.525 -1.195 ;
        RECT 18.195 -2.885 18.525 -2.555 ;
        RECT 18.2 -3.56 18.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.555 129.8 19.885 130.93 ;
        RECT 19.555 127.675 19.885 128.005 ;
        RECT 19.555 126.315 19.885 126.645 ;
        RECT 19.555 124.955 19.885 125.285 ;
        RECT 19.555 123.595 19.885 123.925 ;
        RECT 19.56 123.595 19.88 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.555 -1.525 19.885 -1.195 ;
        RECT 19.555 -2.885 19.885 -2.555 ;
        RECT 19.56 -3.56 19.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.555 -118.485 19.885 -118.155 ;
        RECT 19.555 -119.845 19.885 -119.515 ;
        RECT 19.555 -121.205 19.885 -120.875 ;
        RECT 19.555 -122.565 19.885 -122.235 ;
        RECT 19.555 -123.925 19.885 -123.595 ;
        RECT 19.555 -125.285 19.885 -124.955 ;
        RECT 19.555 -126.645 19.885 -126.315 ;
        RECT 19.555 -128.005 19.885 -127.675 ;
        RECT 19.555 -129.365 19.885 -129.035 ;
        RECT 19.555 -130.725 19.885 -130.395 ;
        RECT 19.555 -132.085 19.885 -131.755 ;
        RECT 19.555 -133.445 19.885 -133.115 ;
        RECT 19.555 -134.805 19.885 -134.475 ;
        RECT 19.555 -136.165 19.885 -135.835 ;
        RECT 19.555 -137.525 19.885 -137.195 ;
        RECT 19.555 -138.885 19.885 -138.555 ;
        RECT 19.555 -140.245 19.885 -139.915 ;
        RECT 19.555 -141.605 19.885 -141.275 ;
        RECT 19.555 -142.965 19.885 -142.635 ;
        RECT 19.555 -144.325 19.885 -143.995 ;
        RECT 19.555 -145.685 19.885 -145.355 ;
        RECT 19.555 -147.045 19.885 -146.715 ;
        RECT 19.555 -148.405 19.885 -148.075 ;
        RECT 19.555 -149.765 19.885 -149.435 ;
        RECT 19.555 -151.125 19.885 -150.795 ;
        RECT 19.555 -152.485 19.885 -152.155 ;
        RECT 19.555 -153.845 19.885 -153.515 ;
        RECT 19.555 -155.205 19.885 -154.875 ;
        RECT 19.555 -156.565 19.885 -156.235 ;
        RECT 19.555 -157.925 19.885 -157.595 ;
        RECT 19.555 -159.285 19.885 -158.955 ;
        RECT 19.555 -160.645 19.885 -160.315 ;
        RECT 19.555 -162.005 19.885 -161.675 ;
        RECT 19.555 -163.365 19.885 -163.035 ;
        RECT 19.555 -164.725 19.885 -164.395 ;
        RECT 19.555 -166.085 19.885 -165.755 ;
        RECT 19.555 -167.445 19.885 -167.115 ;
        RECT 19.555 -168.805 19.885 -168.475 ;
        RECT 19.555 -170.165 19.885 -169.835 ;
        RECT 19.555 -171.525 19.885 -171.195 ;
        RECT 19.555 -172.885 19.885 -172.555 ;
        RECT 19.555 -174.245 19.885 -173.915 ;
        RECT 19.555 -175.605 19.885 -175.275 ;
        RECT 19.555 -176.965 19.885 -176.635 ;
        RECT 19.555 -178.325 19.885 -177.995 ;
        RECT 19.555 -179.685 19.885 -179.355 ;
        RECT 19.555 -181.045 19.885 -180.715 ;
        RECT 19.555 -182.405 19.885 -182.075 ;
        RECT 19.555 -183.765 19.885 -183.435 ;
        RECT 19.555 -185.125 19.885 -184.795 ;
        RECT 19.555 -186.485 19.885 -186.155 ;
        RECT 19.555 -187.845 19.885 -187.515 ;
        RECT 19.555 -189.205 19.885 -188.875 ;
        RECT 19.555 -190.565 19.885 -190.235 ;
        RECT 19.555 -191.925 19.885 -191.595 ;
        RECT 19.555 -193.285 19.885 -192.955 ;
        RECT 19.555 -194.645 19.885 -194.315 ;
        RECT 19.555 -196.005 19.885 -195.675 ;
        RECT 19.555 -197.365 19.885 -197.035 ;
        RECT 19.555 -198.725 19.885 -198.395 ;
        RECT 19.555 -200.085 19.885 -199.755 ;
        RECT 19.555 -201.445 19.885 -201.115 ;
        RECT 19.555 -202.805 19.885 -202.475 ;
        RECT 19.555 -204.165 19.885 -203.835 ;
        RECT 19.555 -205.525 19.885 -205.195 ;
        RECT 19.555 -206.885 19.885 -206.555 ;
        RECT 19.555 -208.245 19.885 -207.915 ;
        RECT 19.555 -209.605 19.885 -209.275 ;
        RECT 19.555 -210.965 19.885 -210.635 ;
        RECT 19.555 -212.325 19.885 -211.995 ;
        RECT 19.555 -213.685 19.885 -213.355 ;
        RECT 19.555 -215.045 19.885 -214.715 ;
        RECT 19.555 -216.405 19.885 -216.075 ;
        RECT 19.555 -217.765 19.885 -217.435 ;
        RECT 19.555 -219.125 19.885 -218.795 ;
        RECT 19.555 -221.37 19.885 -220.24 ;
        RECT 19.56 -221.485 19.88 -118.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.915 129.8 21.245 130.93 ;
        RECT 20.915 127.675 21.245 128.005 ;
        RECT 20.915 126.315 21.245 126.645 ;
        RECT 20.915 124.955 21.245 125.285 ;
        RECT 20.915 123.595 21.245 123.925 ;
        RECT 20.92 123.595 21.24 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.915 -164.725 21.245 -164.395 ;
        RECT 20.915 -166.085 21.245 -165.755 ;
        RECT 20.915 -167.445 21.245 -167.115 ;
        RECT 20.915 -168.805 21.245 -168.475 ;
        RECT 20.915 -170.165 21.245 -169.835 ;
        RECT 20.915 -171.525 21.245 -171.195 ;
        RECT 20.915 -172.885 21.245 -172.555 ;
        RECT 20.915 -174.245 21.245 -173.915 ;
        RECT 20.915 -175.605 21.245 -175.275 ;
        RECT 20.915 -176.965 21.245 -176.635 ;
        RECT 20.915 -178.325 21.245 -177.995 ;
        RECT 20.915 -179.685 21.245 -179.355 ;
        RECT 20.915 -181.045 21.245 -180.715 ;
        RECT 20.915 -182.405 21.245 -182.075 ;
        RECT 20.915 -183.765 21.245 -183.435 ;
        RECT 20.915 -185.125 21.245 -184.795 ;
        RECT 20.915 -186.485 21.245 -186.155 ;
        RECT 20.915 -187.845 21.245 -187.515 ;
        RECT 20.915 -189.205 21.245 -188.875 ;
        RECT 20.915 -190.565 21.245 -190.235 ;
        RECT 20.915 -191.925 21.245 -191.595 ;
        RECT 20.915 -193.285 21.245 -192.955 ;
        RECT 20.915 -194.645 21.245 -194.315 ;
        RECT 20.915 -196.005 21.245 -195.675 ;
        RECT 20.915 -197.365 21.245 -197.035 ;
        RECT 20.915 -198.725 21.245 -198.395 ;
        RECT 20.915 -200.085 21.245 -199.755 ;
        RECT 20.915 -201.445 21.245 -201.115 ;
        RECT 20.915 -202.805 21.245 -202.475 ;
        RECT 20.915 -204.165 21.245 -203.835 ;
        RECT 20.915 -205.525 21.245 -205.195 ;
        RECT 20.915 -206.885 21.245 -206.555 ;
        RECT 20.915 -208.245 21.245 -207.915 ;
        RECT 20.915 -209.605 21.245 -209.275 ;
        RECT 20.915 -210.965 21.245 -210.635 ;
        RECT 20.915 -212.325 21.245 -211.995 ;
        RECT 20.915 -213.685 21.245 -213.355 ;
        RECT 20.915 -215.045 21.245 -214.715 ;
        RECT 20.915 -216.405 21.245 -216.075 ;
        RECT 20.915 -217.765 21.245 -217.435 ;
        RECT 20.915 -219.125 21.245 -218.795 ;
        RECT 20.915 -221.37 21.245 -220.24 ;
        RECT 20.92 -221.485 21.24 -122.235 ;
        RECT 20.915 -122.565 21.245 -122.235 ;
        RECT 20.915 -123.925 21.245 -123.595 ;
        RECT 20.915 -125.285 21.245 -124.955 ;
        RECT 20.915 -126.645 21.245 -126.315 ;
        RECT 20.915 -128.005 21.245 -127.675 ;
        RECT 20.915 -129.365 21.245 -129.035 ;
        RECT 20.915 -130.725 21.245 -130.395 ;
        RECT 20.915 -132.085 21.245 -131.755 ;
        RECT 20.915 -133.445 21.245 -133.115 ;
        RECT 20.915 -134.805 21.245 -134.475 ;
        RECT 20.915 -136.165 21.245 -135.835 ;
        RECT 20.915 -137.525 21.245 -137.195 ;
        RECT 20.915 -138.885 21.245 -138.555 ;
        RECT 20.915 -140.245 21.245 -139.915 ;
        RECT 20.915 -141.605 21.245 -141.275 ;
        RECT 20.915 -142.965 21.245 -142.635 ;
        RECT 20.915 -144.325 21.245 -143.995 ;
        RECT 20.915 -145.685 21.245 -145.355 ;
        RECT 20.915 -147.045 21.245 -146.715 ;
        RECT 20.915 -148.405 21.245 -148.075 ;
        RECT 20.915 -149.765 21.245 -149.435 ;
        RECT 20.915 -151.125 21.245 -150.795 ;
        RECT 20.915 -152.485 21.245 -152.155 ;
        RECT 20.915 -153.845 21.245 -153.515 ;
        RECT 20.915 -155.205 21.245 -154.875 ;
        RECT 20.915 -156.565 21.245 -156.235 ;
        RECT 20.915 -157.925 21.245 -157.595 ;
        RECT 20.915 -159.285 21.245 -158.955 ;
        RECT 20.915 -160.645 21.245 -160.315 ;
        RECT 20.915 -162.005 21.245 -161.675 ;
        RECT 20.915 -163.365 21.245 -163.035 ;
    END
    PORT
      LAYER met3 ;
        RECT -6.285 129.8 -5.955 130.93 ;
        RECT -6.285 127.675 -5.955 128.005 ;
        RECT -6.285 126.315 -5.955 126.645 ;
        RECT -6.285 124.955 -5.955 125.285 ;
        RECT -6.285 123.595 -5.955 123.925 ;
        RECT -6.285 -1.525 -5.955 -1.195 ;
        RECT -6.285 -2.885 -5.955 -2.555 ;
        RECT -6.285 -4.245 -5.955 -3.915 ;
        RECT -6.285 -5.605 -5.955 -5.275 ;
        RECT -6.285 -6.965 -5.955 -6.635 ;
        RECT -6.285 -8.325 -5.955 -7.995 ;
        RECT -6.285 -9.685 -5.955 -9.355 ;
        RECT -6.285 -12.405 -5.955 -12.075 ;
        RECT -6.285 -13.765 -5.955 -13.435 ;
        RECT -6.285 -15.125 -5.955 -14.795 ;
        RECT -6.285 -16.485 -5.955 -16.155 ;
        RECT -6.285 -17.845 -5.955 -17.515 ;
        RECT -6.285 -19.205 -5.955 -18.875 ;
        RECT -6.285 -20.565 -5.955 -20.235 ;
        RECT -6.285 -21.925 -5.955 -21.595 ;
        RECT -6.285 -23.285 -5.955 -22.955 ;
        RECT -6.285 -24.645 -5.955 -24.315 ;
        RECT -6.285 -26.005 -5.955 -25.675 ;
        RECT -6.285 -27.365 -5.955 -27.035 ;
        RECT -6.285 -28.725 -5.955 -28.395 ;
        RECT -6.285 -30.085 -5.955 -29.755 ;
        RECT -6.285 -31.445 -5.955 -31.115 ;
        RECT -6.285 -32.805 -5.955 -32.475 ;
        RECT -6.285 -34.165 -5.955 -33.835 ;
        RECT -6.285 -35.525 -5.955 -35.195 ;
        RECT -6.285 -36.885 -5.955 -36.555 ;
        RECT -6.285 -38.245 -5.955 -37.915 ;
        RECT -6.285 -39.605 -5.955 -39.275 ;
        RECT -6.285 -40.965 -5.955 -40.635 ;
        RECT -6.285 -42.325 -5.955 -41.995 ;
        RECT -6.285 -43.685 -5.955 -43.355 ;
        RECT -6.285 -45.045 -5.955 -44.715 ;
        RECT -6.285 -46.405 -5.955 -46.075 ;
        RECT -6.285 -47.765 -5.955 -47.435 ;
        RECT -6.285 -49.125 -5.955 -48.795 ;
        RECT -6.285 -50.485 -5.955 -50.155 ;
        RECT -6.285 -51.845 -5.955 -51.515 ;
        RECT -6.285 -53.205 -5.955 -52.875 ;
        RECT -6.285 -54.565 -5.955 -54.235 ;
        RECT -6.285 -55.925 -5.955 -55.595 ;
        RECT -6.285 -57.285 -5.955 -56.955 ;
        RECT -6.285 -58.645 -5.955 -58.315 ;
        RECT -6.285 -61.365 -5.955 -61.035 ;
        RECT -6.285 -65.445 -5.955 -65.115 ;
        RECT -6.285 -66.805 -5.955 -66.475 ;
        RECT -6.285 -68.165 -5.955 -67.835 ;
        RECT -6.285 -69.525 -5.955 -69.195 ;
        RECT -6.285 -70.885 -5.955 -70.555 ;
        RECT -6.285 -72.245 -5.955 -71.915 ;
        RECT -6.285 -73.605 -5.955 -73.275 ;
        RECT -6.285 -74.965 -5.955 -74.635 ;
        RECT -6.285 -76.325 -5.955 -75.995 ;
        RECT -6.285 -77.685 -5.955 -77.355 ;
        RECT -6.285 -79.045 -5.955 -78.715 ;
        RECT -6.285 -80.405 -5.955 -80.075 ;
        RECT -6.285 -81.765 -5.955 -81.435 ;
        RECT -6.285 -83.125 -5.955 -82.795 ;
        RECT -6.285 -84.485 -5.955 -84.155 ;
        RECT -6.285 -85.845 -5.955 -85.515 ;
        RECT -6.285 -87.205 -5.955 -86.875 ;
        RECT -6.285 -88.565 -5.955 -88.235 ;
        RECT -6.285 -89.925 -5.955 -89.595 ;
        RECT -6.285 -91.285 -5.955 -90.955 ;
        RECT -6.285 -92.645 -5.955 -92.315 ;
        RECT -6.285 -94.005 -5.955 -93.675 ;
        RECT -6.285 -95.365 -5.955 -95.035 ;
        RECT -6.285 -96.725 -5.955 -96.395 ;
        RECT -6.285 -98.085 -5.955 -97.755 ;
        RECT -6.285 -99.445 -5.955 -99.115 ;
        RECT -6.285 -100.805 -5.955 -100.475 ;
        RECT -6.285 -102.165 -5.955 -101.835 ;
        RECT -6.285 -103.525 -5.955 -103.195 ;
        RECT -6.285 -104.885 -5.955 -104.555 ;
        RECT -6.285 -106.245 -5.955 -105.915 ;
        RECT -6.285 -107.605 -5.955 -107.275 ;
        RECT -6.285 -108.965 -5.955 -108.635 ;
        RECT -6.285 -110.325 -5.955 -109.995 ;
        RECT -6.285 -111.685 -5.955 -111.355 ;
        RECT -6.285 -114.405 -5.955 -114.075 ;
        RECT -6.285 -115.765 -5.955 -115.435 ;
        RECT -6.285 -117.125 -5.955 -116.795 ;
        RECT -6.285 -118.485 -5.955 -118.155 ;
        RECT -6.285 -119.845 -5.955 -119.515 ;
        RECT -6.285 -121.205 -5.955 -120.875 ;
        RECT -6.285 -122.565 -5.955 -122.235 ;
        RECT -6.285 -123.925 -5.955 -123.595 ;
        RECT -6.285 -125.285 -5.955 -124.955 ;
        RECT -6.285 -126.645 -5.955 -126.315 ;
        RECT -6.285 -128.005 -5.955 -127.675 ;
        RECT -6.285 -129.365 -5.955 -129.035 ;
        RECT -6.285 -130.725 -5.955 -130.395 ;
        RECT -6.285 -132.085 -5.955 -131.755 ;
        RECT -6.285 -133.445 -5.955 -133.115 ;
        RECT -6.285 -134.805 -5.955 -134.475 ;
        RECT -6.285 -136.165 -5.955 -135.835 ;
        RECT -6.285 -137.525 -5.955 -137.195 ;
        RECT -6.285 -138.885 -5.955 -138.555 ;
        RECT -6.285 -140.245 -5.955 -139.915 ;
        RECT -6.285 -141.605 -5.955 -141.275 ;
        RECT -6.285 -142.965 -5.955 -142.635 ;
        RECT -6.285 -144.325 -5.955 -143.995 ;
        RECT -6.285 -145.685 -5.955 -145.355 ;
        RECT -6.285 -147.045 -5.955 -146.715 ;
        RECT -6.285 -148.405 -5.955 -148.075 ;
        RECT -6.285 -149.765 -5.955 -149.435 ;
        RECT -6.285 -151.125 -5.955 -150.795 ;
        RECT -6.285 -152.485 -5.955 -152.155 ;
        RECT -6.285 -153.845 -5.955 -153.515 ;
        RECT -6.285 -155.205 -5.955 -154.875 ;
        RECT -6.285 -156.565 -5.955 -156.235 ;
        RECT -6.285 -157.925 -5.955 -157.595 ;
        RECT -6.285 -159.285 -5.955 -158.955 ;
        RECT -6.285 -160.645 -5.955 -160.315 ;
        RECT -6.285 -162.005 -5.955 -161.675 ;
        RECT -6.285 -163.365 -5.955 -163.035 ;
        RECT -6.285 -164.725 -5.955 -164.395 ;
        RECT -6.285 -166.085 -5.955 -165.755 ;
        RECT -6.285 -167.445 -5.955 -167.115 ;
        RECT -6.285 -168.805 -5.955 -168.475 ;
        RECT -6.285 -170.165 -5.955 -169.835 ;
        RECT -6.285 -171.525 -5.955 -171.195 ;
        RECT -6.285 -172.885 -5.955 -172.555 ;
        RECT -6.285 -174.245 -5.955 -173.915 ;
        RECT -6.285 -175.605 -5.955 -175.275 ;
        RECT -6.285 -176.965 -5.955 -176.635 ;
        RECT -6.285 -178.325 -5.955 -177.995 ;
        RECT -6.285 -179.685 -5.955 -179.355 ;
        RECT -6.285 -181.045 -5.955 -180.715 ;
        RECT -6.285 -182.405 -5.955 -182.075 ;
        RECT -6.285 -183.765 -5.955 -183.435 ;
        RECT -6.285 -185.125 -5.955 -184.795 ;
        RECT -6.285 -186.485 -5.955 -186.155 ;
        RECT -6.285 -187.845 -5.955 -187.515 ;
        RECT -6.285 -189.205 -5.955 -188.875 ;
        RECT -6.285 -190.565 -5.955 -190.235 ;
        RECT -6.285 -191.925 -5.955 -191.595 ;
        RECT -6.285 -193.285 -5.955 -192.955 ;
        RECT -6.285 -194.645 -5.955 -194.315 ;
        RECT -6.285 -196.005 -5.955 -195.675 ;
        RECT -6.285 -197.365 -5.955 -197.035 ;
        RECT -6.285 -198.725 -5.955 -198.395 ;
        RECT -6.285 -200.085 -5.955 -199.755 ;
        RECT -6.285 -201.445 -5.955 -201.115 ;
        RECT -6.285 -202.805 -5.955 -202.475 ;
        RECT -6.285 -204.165 -5.955 -203.835 ;
        RECT -6.285 -205.525 -5.955 -205.195 ;
        RECT -6.285 -206.885 -5.955 -206.555 ;
        RECT -6.285 -208.245 -5.955 -207.915 ;
        RECT -6.285 -209.605 -5.955 -209.275 ;
        RECT -6.285 -210.965 -5.955 -210.635 ;
        RECT -6.285 -212.325 -5.955 -211.995 ;
        RECT -6.285 -213.685 -5.955 -213.355 ;
        RECT -6.285 -215.045 -5.955 -214.715 ;
        RECT -6.285 -216.405 -5.955 -216.075 ;
        RECT -6.285 -217.765 -5.955 -217.435 ;
        RECT -6.285 -219.125 -5.955 -218.795 ;
        RECT -6.285 -221.37 -5.955 -220.24 ;
        RECT -6.28 -221.485 -5.96 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -4.925 129.8 -4.595 130.93 ;
        RECT -4.925 127.675 -4.595 128.005 ;
        RECT -4.925 126.315 -4.595 126.645 ;
        RECT -4.925 124.955 -4.595 125.285 ;
        RECT -4.925 123.595 -4.595 123.925 ;
        RECT -4.925 122.215 -4.595 122.545 ;
        RECT -4.925 120.165 -4.595 120.495 ;
        RECT -4.925 118.235 -4.595 118.565 ;
        RECT -4.925 116.395 -4.595 116.725 ;
        RECT -4.925 114.905 -4.595 115.235 ;
        RECT -4.925 113.235 -4.595 113.565 ;
        RECT -4.925 111.745 -4.595 112.075 ;
        RECT -4.925 110.075 -4.595 110.405 ;
        RECT -4.925 108.585 -4.595 108.915 ;
        RECT -4.925 106.915 -4.595 107.245 ;
        RECT -4.925 105.425 -4.595 105.755 ;
        RECT -4.925 104.015 -4.595 104.345 ;
        RECT -4.925 102.175 -4.595 102.505 ;
        RECT -4.925 100.685 -4.595 101.015 ;
        RECT -4.925 99.015 -4.595 99.345 ;
        RECT -4.925 97.525 -4.595 97.855 ;
        RECT -4.925 95.855 -4.595 96.185 ;
        RECT -4.925 94.365 -4.595 94.695 ;
        RECT -4.925 92.695 -4.595 93.025 ;
        RECT -4.925 91.205 -4.595 91.535 ;
        RECT -4.925 89.795 -4.595 90.125 ;
        RECT -4.925 87.955 -4.595 88.285 ;
        RECT -4.925 86.465 -4.595 86.795 ;
        RECT -4.925 84.795 -4.595 85.125 ;
        RECT -4.925 83.305 -4.595 83.635 ;
        RECT -4.925 81.635 -4.595 81.965 ;
        RECT -4.925 80.145 -4.595 80.475 ;
        RECT -4.925 78.475 -4.595 78.805 ;
        RECT -4.925 76.985 -4.595 77.315 ;
        RECT -4.925 75.575 -4.595 75.905 ;
        RECT -4.925 73.735 -4.595 74.065 ;
        RECT -4.925 72.245 -4.595 72.575 ;
        RECT -4.925 70.575 -4.595 70.905 ;
        RECT -4.925 69.085 -4.595 69.415 ;
        RECT -4.925 67.415 -4.595 67.745 ;
        RECT -4.925 65.925 -4.595 66.255 ;
        RECT -4.925 64.255 -4.595 64.585 ;
        RECT -4.925 62.765 -4.595 63.095 ;
        RECT -4.925 61.355 -4.595 61.685 ;
        RECT -4.925 59.515 -4.595 59.845 ;
        RECT -4.925 58.025 -4.595 58.355 ;
        RECT -4.925 56.355 -4.595 56.685 ;
        RECT -4.925 54.865 -4.595 55.195 ;
        RECT -4.925 53.195 -4.595 53.525 ;
        RECT -4.925 51.705 -4.595 52.035 ;
        RECT -4.925 50.035 -4.595 50.365 ;
        RECT -4.925 48.545 -4.595 48.875 ;
        RECT -4.925 47.135 -4.595 47.465 ;
        RECT -4.925 45.295 -4.595 45.625 ;
        RECT -4.925 43.805 -4.595 44.135 ;
        RECT -4.925 42.135 -4.595 42.465 ;
        RECT -4.925 40.645 -4.595 40.975 ;
        RECT -4.925 38.975 -4.595 39.305 ;
        RECT -4.925 37.485 -4.595 37.815 ;
        RECT -4.925 35.815 -4.595 36.145 ;
        RECT -4.925 34.325 -4.595 34.655 ;
        RECT -4.925 32.915 -4.595 33.245 ;
        RECT -4.925 31.075 -4.595 31.405 ;
        RECT -4.925 29.585 -4.595 29.915 ;
        RECT -4.925 27.915 -4.595 28.245 ;
        RECT -4.925 26.425 -4.595 26.755 ;
        RECT -4.925 24.755 -4.595 25.085 ;
        RECT -4.925 23.265 -4.595 23.595 ;
        RECT -4.925 21.595 -4.595 21.925 ;
        RECT -4.925 20.105 -4.595 20.435 ;
        RECT -4.925 18.695 -4.595 19.025 ;
        RECT -4.925 16.855 -4.595 17.185 ;
        RECT -4.925 15.365 -4.595 15.695 ;
        RECT -4.925 13.695 -4.595 14.025 ;
        RECT -4.925 12.205 -4.595 12.535 ;
        RECT -4.925 10.535 -4.595 10.865 ;
        RECT -4.925 9.045 -4.595 9.375 ;
        RECT -4.925 7.375 -4.595 7.705 ;
        RECT -4.925 5.885 -4.595 6.215 ;
        RECT -4.925 4.475 -4.595 4.805 ;
        RECT -4.925 2.115 -4.595 2.445 ;
        RECT -4.925 0.06 -4.595 0.39 ;
        RECT -4.925 -1.525 -4.595 -1.195 ;
        RECT -4.925 -2.885 -4.595 -2.555 ;
        RECT -4.925 -4.245 -4.595 -3.915 ;
        RECT -4.925 -5.605 -4.595 -5.275 ;
        RECT -4.925 -6.965 -4.595 -6.635 ;
        RECT -4.925 -8.325 -4.595 -7.995 ;
        RECT -4.925 -9.685 -4.595 -9.355 ;
        RECT -4.925 -12.405 -4.595 -12.075 ;
        RECT -4.925 -13.765 -4.595 -13.435 ;
        RECT -4.925 -15.125 -4.595 -14.795 ;
        RECT -4.925 -16.485 -4.595 -16.155 ;
        RECT -4.925 -17.845 -4.595 -17.515 ;
        RECT -4.925 -19.205 -4.595 -18.875 ;
        RECT -4.925 -20.565 -4.595 -20.235 ;
        RECT -4.925 -21.925 -4.595 -21.595 ;
        RECT -4.925 -23.285 -4.595 -22.955 ;
        RECT -4.925 -24.645 -4.595 -24.315 ;
        RECT -4.925 -26.005 -4.595 -25.675 ;
        RECT -4.925 -27.365 -4.595 -27.035 ;
        RECT -4.925 -28.725 -4.595 -28.395 ;
        RECT -4.925 -30.085 -4.595 -29.755 ;
        RECT -4.925 -31.445 -4.595 -31.115 ;
        RECT -4.925 -32.805 -4.595 -32.475 ;
        RECT -4.925 -34.165 -4.595 -33.835 ;
        RECT -4.925 -35.525 -4.595 -35.195 ;
        RECT -4.925 -36.885 -4.595 -36.555 ;
        RECT -4.925 -38.245 -4.595 -37.915 ;
        RECT -4.925 -39.605 -4.595 -39.275 ;
        RECT -4.925 -40.965 -4.595 -40.635 ;
        RECT -4.925 -42.325 -4.595 -41.995 ;
        RECT -4.925 -43.685 -4.595 -43.355 ;
        RECT -4.925 -45.045 -4.595 -44.715 ;
        RECT -4.925 -46.405 -4.595 -46.075 ;
        RECT -4.925 -47.765 -4.595 -47.435 ;
        RECT -4.925 -49.125 -4.595 -48.795 ;
        RECT -4.925 -50.485 -4.595 -50.155 ;
        RECT -4.925 -51.845 -4.595 -51.515 ;
        RECT -4.925 -53.205 -4.595 -52.875 ;
        RECT -4.925 -54.565 -4.595 -54.235 ;
        RECT -4.925 -55.925 -4.595 -55.595 ;
        RECT -4.925 -57.285 -4.595 -56.955 ;
        RECT -4.925 -58.645 -4.595 -58.315 ;
        RECT -4.925 -61.365 -4.595 -61.035 ;
        RECT -4.925 -65.445 -4.595 -65.115 ;
        RECT -4.925 -66.805 -4.595 -66.475 ;
        RECT -4.925 -68.165 -4.595 -67.835 ;
        RECT -4.925 -69.525 -4.595 -69.195 ;
        RECT -4.925 -70.885 -4.595 -70.555 ;
        RECT -4.925 -72.245 -4.595 -71.915 ;
        RECT -4.925 -73.605 -4.595 -73.275 ;
        RECT -4.925 -74.965 -4.595 -74.635 ;
        RECT -4.925 -76.325 -4.595 -75.995 ;
        RECT -4.925 -77.685 -4.595 -77.355 ;
        RECT -4.925 -79.045 -4.595 -78.715 ;
        RECT -4.925 -80.405 -4.595 -80.075 ;
        RECT -4.925 -81.765 -4.595 -81.435 ;
        RECT -4.925 -83.125 -4.595 -82.795 ;
        RECT -4.925 -84.485 -4.595 -84.155 ;
        RECT -4.925 -85.845 -4.595 -85.515 ;
        RECT -4.925 -87.205 -4.595 -86.875 ;
        RECT -4.925 -88.565 -4.595 -88.235 ;
        RECT -4.925 -89.925 -4.595 -89.595 ;
        RECT -4.925 -91.285 -4.595 -90.955 ;
        RECT -4.925 -92.645 -4.595 -92.315 ;
        RECT -4.925 -94.005 -4.595 -93.675 ;
        RECT -4.925 -95.365 -4.595 -95.035 ;
        RECT -4.925 -96.725 -4.595 -96.395 ;
        RECT -4.925 -98.085 -4.595 -97.755 ;
        RECT -4.925 -99.445 -4.595 -99.115 ;
        RECT -4.925 -100.805 -4.595 -100.475 ;
        RECT -4.925 -102.165 -4.595 -101.835 ;
        RECT -4.925 -103.525 -4.595 -103.195 ;
        RECT -4.925 -104.885 -4.595 -104.555 ;
        RECT -4.925 -106.245 -4.595 -105.915 ;
        RECT -4.925 -107.605 -4.595 -107.275 ;
        RECT -4.925 -108.965 -4.595 -108.635 ;
        RECT -4.925 -110.325 -4.595 -109.995 ;
        RECT -4.925 -111.685 -4.595 -111.355 ;
        RECT -4.925 -114.405 -4.595 -114.075 ;
        RECT -4.925 -115.765 -4.595 -115.435 ;
        RECT -4.925 -117.125 -4.595 -116.795 ;
        RECT -4.925 -118.485 -4.595 -118.155 ;
        RECT -4.925 -119.845 -4.595 -119.515 ;
        RECT -4.925 -121.205 -4.595 -120.875 ;
        RECT -4.925 -122.565 -4.595 -122.235 ;
        RECT -4.925 -123.925 -4.595 -123.595 ;
        RECT -4.925 -125.285 -4.595 -124.955 ;
        RECT -4.925 -126.645 -4.595 -126.315 ;
        RECT -4.925 -128.005 -4.595 -127.675 ;
        RECT -4.925 -129.365 -4.595 -129.035 ;
        RECT -4.925 -130.725 -4.595 -130.395 ;
        RECT -4.925 -132.085 -4.595 -131.755 ;
        RECT -4.925 -133.445 -4.595 -133.115 ;
        RECT -4.925 -134.805 -4.595 -134.475 ;
        RECT -4.925 -136.165 -4.595 -135.835 ;
        RECT -4.925 -137.525 -4.595 -137.195 ;
        RECT -4.925 -138.885 -4.595 -138.555 ;
        RECT -4.925 -140.245 -4.595 -139.915 ;
        RECT -4.925 -141.605 -4.595 -141.275 ;
        RECT -4.925 -142.965 -4.595 -142.635 ;
        RECT -4.925 -144.325 -4.595 -143.995 ;
        RECT -4.925 -145.685 -4.595 -145.355 ;
        RECT -4.925 -147.045 -4.595 -146.715 ;
        RECT -4.925 -148.405 -4.595 -148.075 ;
        RECT -4.925 -149.765 -4.595 -149.435 ;
        RECT -4.925 -151.125 -4.595 -150.795 ;
        RECT -4.925 -152.485 -4.595 -152.155 ;
        RECT -4.925 -153.845 -4.595 -153.515 ;
        RECT -4.925 -155.205 -4.595 -154.875 ;
        RECT -4.925 -156.565 -4.595 -156.235 ;
        RECT -4.925 -157.925 -4.595 -157.595 ;
        RECT -4.925 -159.285 -4.595 -158.955 ;
        RECT -4.925 -160.645 -4.595 -160.315 ;
        RECT -4.925 -162.005 -4.595 -161.675 ;
        RECT -4.925 -163.365 -4.595 -163.035 ;
        RECT -4.925 -164.725 -4.595 -164.395 ;
        RECT -4.925 -166.085 -4.595 -165.755 ;
        RECT -4.925 -167.445 -4.595 -167.115 ;
        RECT -4.925 -168.805 -4.595 -168.475 ;
        RECT -4.925 -170.165 -4.595 -169.835 ;
        RECT -4.925 -171.525 -4.595 -171.195 ;
        RECT -4.925 -172.885 -4.595 -172.555 ;
        RECT -4.925 -174.245 -4.595 -173.915 ;
        RECT -4.925 -175.605 -4.595 -175.275 ;
        RECT -4.925 -176.965 -4.595 -176.635 ;
        RECT -4.925 -178.325 -4.595 -177.995 ;
        RECT -4.925 -179.685 -4.595 -179.355 ;
        RECT -4.925 -181.045 -4.595 -180.715 ;
        RECT -4.925 -182.405 -4.595 -182.075 ;
        RECT -4.925 -183.765 -4.595 -183.435 ;
        RECT -4.925 -185.125 -4.595 -184.795 ;
        RECT -4.925 -186.485 -4.595 -186.155 ;
        RECT -4.925 -187.845 -4.595 -187.515 ;
        RECT -4.925 -189.205 -4.595 -188.875 ;
        RECT -4.925 -190.565 -4.595 -190.235 ;
        RECT -4.925 -191.925 -4.595 -191.595 ;
        RECT -4.925 -193.285 -4.595 -192.955 ;
        RECT -4.925 -194.645 -4.595 -194.315 ;
        RECT -4.925 -196.005 -4.595 -195.675 ;
        RECT -4.925 -197.365 -4.595 -197.035 ;
        RECT -4.925 -198.725 -4.595 -198.395 ;
        RECT -4.925 -200.085 -4.595 -199.755 ;
        RECT -4.925 -201.445 -4.595 -201.115 ;
        RECT -4.925 -202.805 -4.595 -202.475 ;
        RECT -4.925 -204.165 -4.595 -203.835 ;
        RECT -4.925 -205.525 -4.595 -205.195 ;
        RECT -4.925 -206.885 -4.595 -206.555 ;
        RECT -4.925 -208.245 -4.595 -207.915 ;
        RECT -4.925 -209.605 -4.595 -209.275 ;
        RECT -4.925 -210.965 -4.595 -210.635 ;
        RECT -4.925 -212.325 -4.595 -211.995 ;
        RECT -4.925 -213.685 -4.595 -213.355 ;
        RECT -4.925 -215.045 -4.595 -214.715 ;
        RECT -4.925 -216.405 -4.595 -216.075 ;
        RECT -4.925 -217.765 -4.595 -217.435 ;
        RECT -4.925 -219.125 -4.595 -218.795 ;
        RECT -4.925 -221.37 -4.595 -220.24 ;
        RECT -4.92 -221.485 -4.6 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -3.565 129.8 -3.235 130.93 ;
        RECT -3.565 127.675 -3.235 128.005 ;
        RECT -3.565 126.315 -3.235 126.645 ;
        RECT -3.565 124.955 -3.235 125.285 ;
        RECT -3.565 123.595 -3.235 123.925 ;
        RECT -3.565 122.215 -3.235 122.545 ;
        RECT -3.565 120.165 -3.235 120.495 ;
        RECT -3.565 118.235 -3.235 118.565 ;
        RECT -3.565 116.395 -3.235 116.725 ;
        RECT -3.565 114.905 -3.235 115.235 ;
        RECT -3.565 113.235 -3.235 113.565 ;
        RECT -3.565 111.745 -3.235 112.075 ;
        RECT -3.565 110.075 -3.235 110.405 ;
        RECT -3.565 108.585 -3.235 108.915 ;
        RECT -3.565 106.915 -3.235 107.245 ;
        RECT -3.565 105.425 -3.235 105.755 ;
        RECT -3.565 104.015 -3.235 104.345 ;
        RECT -3.565 102.175 -3.235 102.505 ;
        RECT -3.565 100.685 -3.235 101.015 ;
        RECT -3.565 99.015 -3.235 99.345 ;
        RECT -3.565 97.525 -3.235 97.855 ;
        RECT -3.565 95.855 -3.235 96.185 ;
        RECT -3.565 94.365 -3.235 94.695 ;
        RECT -3.565 92.695 -3.235 93.025 ;
        RECT -3.565 91.205 -3.235 91.535 ;
        RECT -3.565 89.795 -3.235 90.125 ;
        RECT -3.565 87.955 -3.235 88.285 ;
        RECT -3.565 86.465 -3.235 86.795 ;
        RECT -3.565 84.795 -3.235 85.125 ;
        RECT -3.565 83.305 -3.235 83.635 ;
        RECT -3.565 81.635 -3.235 81.965 ;
        RECT -3.565 80.145 -3.235 80.475 ;
        RECT -3.565 78.475 -3.235 78.805 ;
        RECT -3.565 76.985 -3.235 77.315 ;
        RECT -3.565 75.575 -3.235 75.905 ;
        RECT -3.565 73.735 -3.235 74.065 ;
        RECT -3.565 72.245 -3.235 72.575 ;
        RECT -3.565 70.575 -3.235 70.905 ;
        RECT -3.565 69.085 -3.235 69.415 ;
        RECT -3.565 67.415 -3.235 67.745 ;
        RECT -3.565 65.925 -3.235 66.255 ;
        RECT -3.565 64.255 -3.235 64.585 ;
        RECT -3.565 62.765 -3.235 63.095 ;
        RECT -3.565 61.355 -3.235 61.685 ;
        RECT -3.565 59.515 -3.235 59.845 ;
        RECT -3.565 58.025 -3.235 58.355 ;
        RECT -3.565 56.355 -3.235 56.685 ;
        RECT -3.565 54.865 -3.235 55.195 ;
        RECT -3.565 53.195 -3.235 53.525 ;
        RECT -3.565 51.705 -3.235 52.035 ;
        RECT -3.565 50.035 -3.235 50.365 ;
        RECT -3.565 48.545 -3.235 48.875 ;
        RECT -3.565 47.135 -3.235 47.465 ;
        RECT -3.565 45.295 -3.235 45.625 ;
        RECT -3.565 43.805 -3.235 44.135 ;
        RECT -3.565 42.135 -3.235 42.465 ;
        RECT -3.565 40.645 -3.235 40.975 ;
        RECT -3.565 38.975 -3.235 39.305 ;
        RECT -3.565 37.485 -3.235 37.815 ;
        RECT -3.565 35.815 -3.235 36.145 ;
        RECT -3.565 34.325 -3.235 34.655 ;
        RECT -3.565 32.915 -3.235 33.245 ;
        RECT -3.565 31.075 -3.235 31.405 ;
        RECT -3.565 29.585 -3.235 29.915 ;
        RECT -3.565 27.915 -3.235 28.245 ;
        RECT -3.565 26.425 -3.235 26.755 ;
        RECT -3.565 24.755 -3.235 25.085 ;
        RECT -3.565 23.265 -3.235 23.595 ;
        RECT -3.565 21.595 -3.235 21.925 ;
        RECT -3.565 20.105 -3.235 20.435 ;
        RECT -3.565 18.695 -3.235 19.025 ;
        RECT -3.565 16.855 -3.235 17.185 ;
        RECT -3.565 15.365 -3.235 15.695 ;
        RECT -3.565 13.695 -3.235 14.025 ;
        RECT -3.565 12.205 -3.235 12.535 ;
        RECT -3.565 10.535 -3.235 10.865 ;
        RECT -3.565 9.045 -3.235 9.375 ;
        RECT -3.565 7.375 -3.235 7.705 ;
        RECT -3.565 5.885 -3.235 6.215 ;
        RECT -3.565 4.475 -3.235 4.805 ;
        RECT -3.565 2.115 -3.235 2.445 ;
        RECT -3.565 0.06 -3.235 0.39 ;
        RECT -3.565 -1.525 -3.235 -1.195 ;
        RECT -3.565 -2.885 -3.235 -2.555 ;
        RECT -3.565 -4.245 -3.235 -3.915 ;
        RECT -3.565 -5.605 -3.235 -5.275 ;
        RECT -3.565 -6.965 -3.235 -6.635 ;
        RECT -3.565 -8.325 -3.235 -7.995 ;
        RECT -3.565 -9.685 -3.235 -9.355 ;
        RECT -3.565 -12.405 -3.235 -12.075 ;
        RECT -3.565 -13.765 -3.235 -13.435 ;
        RECT -3.565 -15.125 -3.235 -14.795 ;
        RECT -3.565 -16.485 -3.235 -16.155 ;
        RECT -3.565 -17.845 -3.235 -17.515 ;
        RECT -3.565 -19.205 -3.235 -18.875 ;
        RECT -3.565 -20.565 -3.235 -20.235 ;
        RECT -3.565 -21.925 -3.235 -21.595 ;
        RECT -3.565 -23.285 -3.235 -22.955 ;
        RECT -3.565 -24.645 -3.235 -24.315 ;
        RECT -3.565 -26.005 -3.235 -25.675 ;
        RECT -3.565 -27.365 -3.235 -27.035 ;
        RECT -3.565 -28.725 -3.235 -28.395 ;
        RECT -3.565 -30.085 -3.235 -29.755 ;
        RECT -3.565 -31.445 -3.235 -31.115 ;
        RECT -3.565 -32.805 -3.235 -32.475 ;
        RECT -3.565 -34.165 -3.235 -33.835 ;
        RECT -3.565 -35.525 -3.235 -35.195 ;
        RECT -3.565 -36.885 -3.235 -36.555 ;
        RECT -3.565 -38.245 -3.235 -37.915 ;
        RECT -3.565 -39.605 -3.235 -39.275 ;
        RECT -3.565 -40.965 -3.235 -40.635 ;
        RECT -3.565 -42.325 -3.235 -41.995 ;
        RECT -3.565 -43.685 -3.235 -43.355 ;
        RECT -3.565 -45.045 -3.235 -44.715 ;
        RECT -3.565 -46.405 -3.235 -46.075 ;
        RECT -3.565 -47.765 -3.235 -47.435 ;
        RECT -3.565 -49.125 -3.235 -48.795 ;
        RECT -3.565 -50.485 -3.235 -50.155 ;
        RECT -3.565 -51.845 -3.235 -51.515 ;
        RECT -3.565 -53.205 -3.235 -52.875 ;
        RECT -3.565 -54.565 -3.235 -54.235 ;
        RECT -3.565 -55.925 -3.235 -55.595 ;
        RECT -3.565 -57.285 -3.235 -56.955 ;
        RECT -3.565 -58.645 -3.235 -58.315 ;
        RECT -3.565 -61.365 -3.235 -61.035 ;
        RECT -3.565 -65.445 -3.235 -65.115 ;
        RECT -3.565 -66.805 -3.235 -66.475 ;
        RECT -3.565 -68.165 -3.235 -67.835 ;
        RECT -3.565 -69.525 -3.235 -69.195 ;
        RECT -3.565 -70.885 -3.235 -70.555 ;
        RECT -3.565 -72.245 -3.235 -71.915 ;
        RECT -3.565 -73.605 -3.235 -73.275 ;
        RECT -3.565 -74.965 -3.235 -74.635 ;
        RECT -3.565 -76.325 -3.235 -75.995 ;
        RECT -3.565 -77.685 -3.235 -77.355 ;
        RECT -3.565 -79.045 -3.235 -78.715 ;
        RECT -3.565 -80.405 -3.235 -80.075 ;
        RECT -3.565 -81.765 -3.235 -81.435 ;
        RECT -3.565 -83.125 -3.235 -82.795 ;
        RECT -3.565 -84.485 -3.235 -84.155 ;
        RECT -3.565 -85.845 -3.235 -85.515 ;
        RECT -3.565 -87.205 -3.235 -86.875 ;
        RECT -3.565 -88.565 -3.235 -88.235 ;
        RECT -3.565 -89.925 -3.235 -89.595 ;
        RECT -3.565 -91.285 -3.235 -90.955 ;
        RECT -3.565 -92.645 -3.235 -92.315 ;
        RECT -3.565 -94.005 -3.235 -93.675 ;
        RECT -3.565 -95.365 -3.235 -95.035 ;
        RECT -3.565 -96.725 -3.235 -96.395 ;
        RECT -3.565 -98.085 -3.235 -97.755 ;
        RECT -3.565 -99.445 -3.235 -99.115 ;
        RECT -3.565 -100.805 -3.235 -100.475 ;
        RECT -3.565 -102.165 -3.235 -101.835 ;
        RECT -3.565 -103.525 -3.235 -103.195 ;
        RECT -3.565 -104.885 -3.235 -104.555 ;
        RECT -3.565 -106.245 -3.235 -105.915 ;
        RECT -3.565 -107.605 -3.235 -107.275 ;
        RECT -3.565 -108.965 -3.235 -108.635 ;
        RECT -3.565 -110.325 -3.235 -109.995 ;
        RECT -3.565 -111.685 -3.235 -111.355 ;
        RECT -3.565 -114.405 -3.235 -114.075 ;
        RECT -3.565 -115.765 -3.235 -115.435 ;
        RECT -3.565 -117.125 -3.235 -116.795 ;
        RECT -3.565 -118.485 -3.235 -118.155 ;
        RECT -3.565 -119.845 -3.235 -119.515 ;
        RECT -3.565 -121.205 -3.235 -120.875 ;
        RECT -3.565 -122.565 -3.235 -122.235 ;
        RECT -3.565 -123.925 -3.235 -123.595 ;
        RECT -3.565 -125.285 -3.235 -124.955 ;
        RECT -3.565 -126.645 -3.235 -126.315 ;
        RECT -3.565 -128.005 -3.235 -127.675 ;
        RECT -3.565 -129.365 -3.235 -129.035 ;
        RECT -3.565 -130.725 -3.235 -130.395 ;
        RECT -3.565 -132.085 -3.235 -131.755 ;
        RECT -3.565 -133.445 -3.235 -133.115 ;
        RECT -3.565 -134.805 -3.235 -134.475 ;
        RECT -3.565 -136.165 -3.235 -135.835 ;
        RECT -3.565 -137.525 -3.235 -137.195 ;
        RECT -3.565 -138.885 -3.235 -138.555 ;
        RECT -3.565 -140.245 -3.235 -139.915 ;
        RECT -3.565 -141.605 -3.235 -141.275 ;
        RECT -3.565 -142.965 -3.235 -142.635 ;
        RECT -3.565 -144.325 -3.235 -143.995 ;
        RECT -3.565 -145.685 -3.235 -145.355 ;
        RECT -3.565 -147.045 -3.235 -146.715 ;
        RECT -3.565 -148.405 -3.235 -148.075 ;
        RECT -3.565 -149.765 -3.235 -149.435 ;
        RECT -3.565 -151.125 -3.235 -150.795 ;
        RECT -3.565 -152.485 -3.235 -152.155 ;
        RECT -3.565 -153.845 -3.235 -153.515 ;
        RECT -3.565 -155.205 -3.235 -154.875 ;
        RECT -3.565 -156.565 -3.235 -156.235 ;
        RECT -3.565 -157.925 -3.235 -157.595 ;
        RECT -3.565 -159.285 -3.235 -158.955 ;
        RECT -3.565 -160.645 -3.235 -160.315 ;
        RECT -3.565 -162.005 -3.235 -161.675 ;
        RECT -3.565 -163.365 -3.235 -163.035 ;
        RECT -3.565 -164.725 -3.235 -164.395 ;
        RECT -3.565 -166.085 -3.235 -165.755 ;
        RECT -3.565 -167.445 -3.235 -167.115 ;
        RECT -3.565 -168.805 -3.235 -168.475 ;
        RECT -3.565 -170.165 -3.235 -169.835 ;
        RECT -3.565 -171.525 -3.235 -171.195 ;
        RECT -3.565 -172.885 -3.235 -172.555 ;
        RECT -3.565 -174.245 -3.235 -173.915 ;
        RECT -3.565 -175.605 -3.235 -175.275 ;
        RECT -3.565 -176.965 -3.235 -176.635 ;
        RECT -3.565 -178.325 -3.235 -177.995 ;
        RECT -3.565 -179.685 -3.235 -179.355 ;
        RECT -3.565 -181.045 -3.235 -180.715 ;
        RECT -3.565 -182.405 -3.235 -182.075 ;
        RECT -3.565 -183.765 -3.235 -183.435 ;
        RECT -3.565 -185.125 -3.235 -184.795 ;
        RECT -3.565 -186.485 -3.235 -186.155 ;
        RECT -3.565 -187.845 -3.235 -187.515 ;
        RECT -3.565 -189.205 -3.235 -188.875 ;
        RECT -3.565 -190.565 -3.235 -190.235 ;
        RECT -3.565 -191.925 -3.235 -191.595 ;
        RECT -3.565 -193.285 -3.235 -192.955 ;
        RECT -3.565 -194.645 -3.235 -194.315 ;
        RECT -3.565 -196.005 -3.235 -195.675 ;
        RECT -3.565 -197.365 -3.235 -197.035 ;
        RECT -3.565 -198.725 -3.235 -198.395 ;
        RECT -3.565 -200.085 -3.235 -199.755 ;
        RECT -3.565 -201.445 -3.235 -201.115 ;
        RECT -3.565 -202.805 -3.235 -202.475 ;
        RECT -3.565 -204.165 -3.235 -203.835 ;
        RECT -3.565 -205.525 -3.235 -205.195 ;
        RECT -3.565 -206.885 -3.235 -206.555 ;
        RECT -3.565 -208.245 -3.235 -207.915 ;
        RECT -3.565 -209.605 -3.235 -209.275 ;
        RECT -3.565 -210.965 -3.235 -210.635 ;
        RECT -3.565 -212.325 -3.235 -211.995 ;
        RECT -3.565 -213.685 -3.235 -213.355 ;
        RECT -3.565 -215.045 -3.235 -214.715 ;
        RECT -3.565 -216.405 -3.235 -216.075 ;
        RECT -3.565 -217.765 -3.235 -217.435 ;
        RECT -3.565 -219.125 -3.235 -218.795 ;
        RECT -3.565 -221.37 -3.235 -220.24 ;
        RECT -3.56 -221.485 -3.24 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -2.205 129.8 -1.875 130.93 ;
        RECT -2.205 127.675 -1.875 128.005 ;
        RECT -2.205 126.315 -1.875 126.645 ;
        RECT -2.205 124.955 -1.875 125.285 ;
        RECT -2.205 123.595 -1.875 123.925 ;
        RECT -2.205 122.215 -1.875 122.545 ;
        RECT -2.205 120.165 -1.875 120.495 ;
        RECT -2.205 118.235 -1.875 118.565 ;
        RECT -2.205 116.395 -1.875 116.725 ;
        RECT -2.205 114.905 -1.875 115.235 ;
        RECT -2.205 113.235 -1.875 113.565 ;
        RECT -2.205 111.745 -1.875 112.075 ;
        RECT -2.205 110.075 -1.875 110.405 ;
        RECT -2.205 108.585 -1.875 108.915 ;
        RECT -2.205 106.915 -1.875 107.245 ;
        RECT -2.205 105.425 -1.875 105.755 ;
        RECT -2.205 104.015 -1.875 104.345 ;
        RECT -2.205 102.175 -1.875 102.505 ;
        RECT -2.205 100.685 -1.875 101.015 ;
        RECT -2.205 99.015 -1.875 99.345 ;
        RECT -2.205 97.525 -1.875 97.855 ;
        RECT -2.205 95.855 -1.875 96.185 ;
        RECT -2.205 94.365 -1.875 94.695 ;
        RECT -2.205 92.695 -1.875 93.025 ;
        RECT -2.205 91.205 -1.875 91.535 ;
        RECT -2.205 89.795 -1.875 90.125 ;
        RECT -2.205 87.955 -1.875 88.285 ;
        RECT -2.205 86.465 -1.875 86.795 ;
        RECT -2.205 84.795 -1.875 85.125 ;
        RECT -2.205 83.305 -1.875 83.635 ;
        RECT -2.205 81.635 -1.875 81.965 ;
        RECT -2.205 80.145 -1.875 80.475 ;
        RECT -2.205 78.475 -1.875 78.805 ;
        RECT -2.205 76.985 -1.875 77.315 ;
        RECT -2.205 75.575 -1.875 75.905 ;
        RECT -2.205 73.735 -1.875 74.065 ;
        RECT -2.205 72.245 -1.875 72.575 ;
        RECT -2.205 70.575 -1.875 70.905 ;
        RECT -2.205 69.085 -1.875 69.415 ;
        RECT -2.205 67.415 -1.875 67.745 ;
        RECT -2.205 65.925 -1.875 66.255 ;
        RECT -2.205 64.255 -1.875 64.585 ;
        RECT -2.205 62.765 -1.875 63.095 ;
        RECT -2.205 61.355 -1.875 61.685 ;
        RECT -2.205 59.515 -1.875 59.845 ;
        RECT -2.205 58.025 -1.875 58.355 ;
        RECT -2.205 56.355 -1.875 56.685 ;
        RECT -2.205 54.865 -1.875 55.195 ;
        RECT -2.205 53.195 -1.875 53.525 ;
        RECT -2.205 51.705 -1.875 52.035 ;
        RECT -2.205 50.035 -1.875 50.365 ;
        RECT -2.205 48.545 -1.875 48.875 ;
        RECT -2.205 47.135 -1.875 47.465 ;
        RECT -2.205 45.295 -1.875 45.625 ;
        RECT -2.205 43.805 -1.875 44.135 ;
        RECT -2.205 42.135 -1.875 42.465 ;
        RECT -2.205 40.645 -1.875 40.975 ;
        RECT -2.205 38.975 -1.875 39.305 ;
        RECT -2.205 37.485 -1.875 37.815 ;
        RECT -2.205 35.815 -1.875 36.145 ;
        RECT -2.205 34.325 -1.875 34.655 ;
        RECT -2.205 32.915 -1.875 33.245 ;
        RECT -2.205 31.075 -1.875 31.405 ;
        RECT -2.205 29.585 -1.875 29.915 ;
        RECT -2.205 27.915 -1.875 28.245 ;
        RECT -2.205 26.425 -1.875 26.755 ;
        RECT -2.205 24.755 -1.875 25.085 ;
        RECT -2.205 23.265 -1.875 23.595 ;
        RECT -2.205 21.595 -1.875 21.925 ;
        RECT -2.205 20.105 -1.875 20.435 ;
        RECT -2.205 18.695 -1.875 19.025 ;
        RECT -2.205 16.855 -1.875 17.185 ;
        RECT -2.205 15.365 -1.875 15.695 ;
        RECT -2.205 13.695 -1.875 14.025 ;
        RECT -2.205 12.205 -1.875 12.535 ;
        RECT -2.205 10.535 -1.875 10.865 ;
        RECT -2.205 9.045 -1.875 9.375 ;
        RECT -2.205 7.375 -1.875 7.705 ;
        RECT -2.205 5.885 -1.875 6.215 ;
        RECT -2.205 4.475 -1.875 4.805 ;
        RECT -2.205 2.115 -1.875 2.445 ;
        RECT -2.205 0.06 -1.875 0.39 ;
        RECT -2.205 -1.525 -1.875 -1.195 ;
        RECT -2.205 -2.885 -1.875 -2.555 ;
        RECT -2.205 -4.245 -1.875 -3.915 ;
        RECT -2.205 -5.605 -1.875 -5.275 ;
        RECT -2.205 -6.965 -1.875 -6.635 ;
        RECT -2.205 -8.325 -1.875 -7.995 ;
        RECT -2.205 -9.685 -1.875 -9.355 ;
        RECT -2.205 -12.405 -1.875 -12.075 ;
        RECT -2.205 -13.765 -1.875 -13.435 ;
        RECT -2.205 -15.125 -1.875 -14.795 ;
        RECT -2.205 -16.485 -1.875 -16.155 ;
        RECT -2.205 -17.845 -1.875 -17.515 ;
        RECT -2.205 -19.205 -1.875 -18.875 ;
        RECT -2.205 -20.565 -1.875 -20.235 ;
        RECT -2.205 -21.925 -1.875 -21.595 ;
        RECT -2.205 -23.285 -1.875 -22.955 ;
        RECT -2.205 -24.645 -1.875 -24.315 ;
        RECT -2.205 -26.005 -1.875 -25.675 ;
        RECT -2.205 -27.365 -1.875 -27.035 ;
        RECT -2.205 -28.725 -1.875 -28.395 ;
        RECT -2.205 -30.085 -1.875 -29.755 ;
        RECT -2.205 -31.445 -1.875 -31.115 ;
        RECT -2.205 -32.805 -1.875 -32.475 ;
        RECT -2.205 -34.165 -1.875 -33.835 ;
        RECT -2.205 -35.525 -1.875 -35.195 ;
        RECT -2.205 -36.885 -1.875 -36.555 ;
        RECT -2.205 -38.245 -1.875 -37.915 ;
        RECT -2.205 -39.605 -1.875 -39.275 ;
        RECT -2.205 -40.965 -1.875 -40.635 ;
        RECT -2.205 -42.325 -1.875 -41.995 ;
        RECT -2.205 -43.685 -1.875 -43.355 ;
        RECT -2.205 -45.045 -1.875 -44.715 ;
        RECT -2.205 -46.405 -1.875 -46.075 ;
        RECT -2.205 -47.765 -1.875 -47.435 ;
        RECT -2.205 -49.125 -1.875 -48.795 ;
        RECT -2.205 -50.485 -1.875 -50.155 ;
        RECT -2.205 -51.845 -1.875 -51.515 ;
        RECT -2.205 -53.205 -1.875 -52.875 ;
        RECT -2.205 -54.565 -1.875 -54.235 ;
        RECT -2.205 -55.925 -1.875 -55.595 ;
        RECT -2.205 -57.285 -1.875 -56.955 ;
        RECT -2.205 -58.645 -1.875 -58.315 ;
        RECT -2.205 -61.365 -1.875 -61.035 ;
        RECT -2.205 -65.445 -1.875 -65.115 ;
        RECT -2.205 -66.805 -1.875 -66.475 ;
        RECT -2.205 -68.165 -1.875 -67.835 ;
        RECT -2.205 -69.525 -1.875 -69.195 ;
        RECT -2.205 -70.885 -1.875 -70.555 ;
        RECT -2.205 -72.245 -1.875 -71.915 ;
        RECT -2.205 -73.605 -1.875 -73.275 ;
        RECT -2.205 -74.965 -1.875 -74.635 ;
        RECT -2.205 -76.325 -1.875 -75.995 ;
        RECT -2.205 -77.685 -1.875 -77.355 ;
        RECT -2.205 -79.045 -1.875 -78.715 ;
        RECT -2.205 -80.405 -1.875 -80.075 ;
        RECT -2.205 -81.765 -1.875 -81.435 ;
        RECT -2.205 -83.125 -1.875 -82.795 ;
        RECT -2.205 -84.485 -1.875 -84.155 ;
        RECT -2.205 -85.845 -1.875 -85.515 ;
        RECT -2.205 -87.205 -1.875 -86.875 ;
        RECT -2.205 -88.565 -1.875 -88.235 ;
        RECT -2.205 -89.925 -1.875 -89.595 ;
        RECT -2.205 -91.285 -1.875 -90.955 ;
        RECT -2.205 -92.645 -1.875 -92.315 ;
        RECT -2.205 -94.005 -1.875 -93.675 ;
        RECT -2.205 -95.365 -1.875 -95.035 ;
        RECT -2.205 -96.725 -1.875 -96.395 ;
        RECT -2.205 -98.085 -1.875 -97.755 ;
        RECT -2.205 -99.445 -1.875 -99.115 ;
        RECT -2.205 -100.805 -1.875 -100.475 ;
        RECT -2.205 -102.165 -1.875 -101.835 ;
        RECT -2.205 -103.525 -1.875 -103.195 ;
        RECT -2.205 -104.885 -1.875 -104.555 ;
        RECT -2.205 -106.245 -1.875 -105.915 ;
        RECT -2.205 -107.605 -1.875 -107.275 ;
        RECT -2.205 -108.965 -1.875 -108.635 ;
        RECT -2.205 -110.325 -1.875 -109.995 ;
        RECT -2.205 -111.685 -1.875 -111.355 ;
        RECT -2.205 -114.405 -1.875 -114.075 ;
        RECT -2.205 -115.765 -1.875 -115.435 ;
        RECT -2.205 -117.125 -1.875 -116.795 ;
        RECT -2.205 -118.485 -1.875 -118.155 ;
        RECT -2.205 -119.845 -1.875 -119.515 ;
        RECT -2.205 -121.205 -1.875 -120.875 ;
        RECT -2.205 -122.565 -1.875 -122.235 ;
        RECT -2.205 -123.925 -1.875 -123.595 ;
        RECT -2.205 -125.285 -1.875 -124.955 ;
        RECT -2.205 -126.645 -1.875 -126.315 ;
        RECT -2.205 -128.005 -1.875 -127.675 ;
        RECT -2.205 -129.365 -1.875 -129.035 ;
        RECT -2.205 -130.725 -1.875 -130.395 ;
        RECT -2.205 -132.085 -1.875 -131.755 ;
        RECT -2.205 -133.445 -1.875 -133.115 ;
        RECT -2.205 -134.805 -1.875 -134.475 ;
        RECT -2.205 -136.165 -1.875 -135.835 ;
        RECT -2.205 -137.525 -1.875 -137.195 ;
        RECT -2.205 -138.885 -1.875 -138.555 ;
        RECT -2.205 -140.245 -1.875 -139.915 ;
        RECT -2.205 -141.605 -1.875 -141.275 ;
        RECT -2.205 -142.965 -1.875 -142.635 ;
        RECT -2.205 -144.325 -1.875 -143.995 ;
        RECT -2.205 -145.685 -1.875 -145.355 ;
        RECT -2.205 -147.045 -1.875 -146.715 ;
        RECT -2.205 -148.405 -1.875 -148.075 ;
        RECT -2.205 -149.765 -1.875 -149.435 ;
        RECT -2.205 -151.125 -1.875 -150.795 ;
        RECT -2.205 -152.485 -1.875 -152.155 ;
        RECT -2.205 -153.845 -1.875 -153.515 ;
        RECT -2.205 -155.205 -1.875 -154.875 ;
        RECT -2.205 -156.565 -1.875 -156.235 ;
        RECT -2.205 -157.925 -1.875 -157.595 ;
        RECT -2.205 -159.285 -1.875 -158.955 ;
        RECT -2.205 -160.645 -1.875 -160.315 ;
        RECT -2.205 -162.005 -1.875 -161.675 ;
        RECT -2.205 -163.365 -1.875 -163.035 ;
        RECT -2.205 -164.725 -1.875 -164.395 ;
        RECT -2.205 -166.085 -1.875 -165.755 ;
        RECT -2.205 -167.445 -1.875 -167.115 ;
        RECT -2.205 -168.805 -1.875 -168.475 ;
        RECT -2.205 -170.165 -1.875 -169.835 ;
        RECT -2.205 -171.525 -1.875 -171.195 ;
        RECT -2.205 -172.885 -1.875 -172.555 ;
        RECT -2.205 -174.245 -1.875 -173.915 ;
        RECT -2.205 -175.605 -1.875 -175.275 ;
        RECT -2.205 -176.965 -1.875 -176.635 ;
        RECT -2.205 -178.325 -1.875 -177.995 ;
        RECT -2.205 -179.685 -1.875 -179.355 ;
        RECT -2.205 -181.045 -1.875 -180.715 ;
        RECT -2.205 -182.405 -1.875 -182.075 ;
        RECT -2.205 -183.765 -1.875 -183.435 ;
        RECT -2.205 -185.125 -1.875 -184.795 ;
        RECT -2.205 -186.485 -1.875 -186.155 ;
        RECT -2.205 -187.845 -1.875 -187.515 ;
        RECT -2.205 -189.205 -1.875 -188.875 ;
        RECT -2.205 -190.565 -1.875 -190.235 ;
        RECT -2.205 -191.925 -1.875 -191.595 ;
        RECT -2.205 -193.285 -1.875 -192.955 ;
        RECT -2.205 -194.645 -1.875 -194.315 ;
        RECT -2.205 -196.005 -1.875 -195.675 ;
        RECT -2.205 -197.365 -1.875 -197.035 ;
        RECT -2.205 -198.725 -1.875 -198.395 ;
        RECT -2.205 -200.085 -1.875 -199.755 ;
        RECT -2.205 -201.445 -1.875 -201.115 ;
        RECT -2.205 -202.805 -1.875 -202.475 ;
        RECT -2.205 -204.165 -1.875 -203.835 ;
        RECT -2.205 -205.525 -1.875 -205.195 ;
        RECT -2.205 -206.885 -1.875 -206.555 ;
        RECT -2.205 -208.245 -1.875 -207.915 ;
        RECT -2.205 -209.605 -1.875 -209.275 ;
        RECT -2.205 -210.965 -1.875 -210.635 ;
        RECT -2.205 -212.325 -1.875 -211.995 ;
        RECT -2.205 -213.685 -1.875 -213.355 ;
        RECT -2.205 -215.045 -1.875 -214.715 ;
        RECT -2.205 -216.405 -1.875 -216.075 ;
        RECT -2.205 -217.765 -1.875 -217.435 ;
        RECT -2.205 -219.125 -1.875 -218.795 ;
        RECT -2.205 -221.37 -1.875 -220.24 ;
        RECT -2.2 -221.485 -1.88 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.845 -87.205 -0.515 -86.875 ;
        RECT -0.845 -88.565 -0.515 -88.235 ;
        RECT -0.845 -89.925 -0.515 -89.595 ;
        RECT -0.845 -91.285 -0.515 -90.955 ;
        RECT -0.845 -92.645 -0.515 -92.315 ;
        RECT -0.845 -94.005 -0.515 -93.675 ;
        RECT -0.845 -95.365 -0.515 -95.035 ;
        RECT -0.845 -96.725 -0.515 -96.395 ;
        RECT -0.845 -98.085 -0.515 -97.755 ;
        RECT -0.845 -99.445 -0.515 -99.115 ;
        RECT -0.845 -100.805 -0.515 -100.475 ;
        RECT -0.845 -102.165 -0.515 -101.835 ;
        RECT -0.845 -103.525 -0.515 -103.195 ;
        RECT -0.845 -104.885 -0.515 -104.555 ;
        RECT -0.845 -106.245 -0.515 -105.915 ;
        RECT -0.845 -107.605 -0.515 -107.275 ;
        RECT -0.845 -108.965 -0.515 -108.635 ;
        RECT -0.845 -110.325 -0.515 -109.995 ;
        RECT -0.845 -111.685 -0.515 -111.355 ;
        RECT -0.845 -114.405 -0.515 -114.075 ;
        RECT -0.845 -115.765 -0.515 -115.435 ;
        RECT -0.845 -117.125 -0.515 -116.795 ;
        RECT -0.845 -118.485 -0.515 -118.155 ;
        RECT -0.845 -119.845 -0.515 -119.515 ;
        RECT -0.845 -121.205 -0.515 -120.875 ;
        RECT -0.845 -122.565 -0.515 -122.235 ;
        RECT -0.845 -123.925 -0.515 -123.595 ;
        RECT -0.845 -125.285 -0.515 -124.955 ;
        RECT -0.845 -126.645 -0.515 -126.315 ;
        RECT -0.845 -128.005 -0.515 -127.675 ;
        RECT -0.845 -129.365 -0.515 -129.035 ;
        RECT -0.845 -130.725 -0.515 -130.395 ;
        RECT -0.845 -132.085 -0.515 -131.755 ;
        RECT -0.845 -133.445 -0.515 -133.115 ;
        RECT -0.845 -134.805 -0.515 -134.475 ;
        RECT -0.845 -136.165 -0.515 -135.835 ;
        RECT -0.845 -137.525 -0.515 -137.195 ;
        RECT -0.845 -138.885 -0.515 -138.555 ;
        RECT -0.845 -140.245 -0.515 -139.915 ;
        RECT -0.845 -141.605 -0.515 -141.275 ;
        RECT -0.845 -142.965 -0.515 -142.635 ;
        RECT -0.845 -144.325 -0.515 -143.995 ;
        RECT -0.845 -145.685 -0.515 -145.355 ;
        RECT -0.845 -147.045 -0.515 -146.715 ;
        RECT -0.845 -148.405 -0.515 -148.075 ;
        RECT -0.845 -149.765 -0.515 -149.435 ;
        RECT -0.845 -151.125 -0.515 -150.795 ;
        RECT -0.845 -152.485 -0.515 -152.155 ;
        RECT -0.845 -153.845 -0.515 -153.515 ;
        RECT -0.845 -155.205 -0.515 -154.875 ;
        RECT -0.845 -156.565 -0.515 -156.235 ;
        RECT -0.845 -157.925 -0.515 -157.595 ;
        RECT -0.845 -159.285 -0.515 -158.955 ;
        RECT -0.845 -160.645 -0.515 -160.315 ;
        RECT -0.845 -162.005 -0.515 -161.675 ;
        RECT -0.845 -163.365 -0.515 -163.035 ;
        RECT -0.845 -164.725 -0.515 -164.395 ;
        RECT -0.845 -166.085 -0.515 -165.755 ;
        RECT -0.845 -167.445 -0.515 -167.115 ;
        RECT -0.845 -168.805 -0.515 -168.475 ;
        RECT -0.845 -170.165 -0.515 -169.835 ;
        RECT -0.845 -171.525 -0.515 -171.195 ;
        RECT -0.845 -172.885 -0.515 -172.555 ;
        RECT -0.845 -174.245 -0.515 -173.915 ;
        RECT -0.845 -175.605 -0.515 -175.275 ;
        RECT -0.845 -176.965 -0.515 -176.635 ;
        RECT -0.845 -178.325 -0.515 -177.995 ;
        RECT -0.845 -179.685 -0.515 -179.355 ;
        RECT -0.845 -181.045 -0.515 -180.715 ;
        RECT -0.845 -182.405 -0.515 -182.075 ;
        RECT -0.845 -183.765 -0.515 -183.435 ;
        RECT -0.845 -185.125 -0.515 -184.795 ;
        RECT -0.845 -186.485 -0.515 -186.155 ;
        RECT -0.845 -187.845 -0.515 -187.515 ;
        RECT -0.845 -189.205 -0.515 -188.875 ;
        RECT -0.845 -190.565 -0.515 -190.235 ;
        RECT -0.845 -191.925 -0.515 -191.595 ;
        RECT -0.845 -193.285 -0.515 -192.955 ;
        RECT -0.845 -194.645 -0.515 -194.315 ;
        RECT -0.845 -196.005 -0.515 -195.675 ;
        RECT -0.845 -197.365 -0.515 -197.035 ;
        RECT -0.845 -198.725 -0.515 -198.395 ;
        RECT -0.845 -200.085 -0.515 -199.755 ;
        RECT -0.845 -201.445 -0.515 -201.115 ;
        RECT -0.845 -202.805 -0.515 -202.475 ;
        RECT -0.845 -204.165 -0.515 -203.835 ;
        RECT -0.845 -205.525 -0.515 -205.195 ;
        RECT -0.845 -206.885 -0.515 -206.555 ;
        RECT -0.845 -208.245 -0.515 -207.915 ;
        RECT -0.845 -209.605 -0.515 -209.275 ;
        RECT -0.845 -210.965 -0.515 -210.635 ;
        RECT -0.845 -212.325 -0.515 -211.995 ;
        RECT -0.845 -213.685 -0.515 -213.355 ;
        RECT -0.845 -215.045 -0.515 -214.715 ;
        RECT -0.845 -216.405 -0.515 -216.075 ;
        RECT -0.845 -217.765 -0.515 -217.435 ;
        RECT -0.845 -219.125 -0.515 -218.795 ;
        RECT -0.845 -221.37 -0.515 -220.24 ;
        RECT -0.84 -221.485 -0.52 131.045 ;
        RECT -0.845 129.8 -0.515 130.93 ;
        RECT -0.845 127.675 -0.515 128.005 ;
        RECT -0.845 126.315 -0.515 126.645 ;
        RECT -0.845 124.955 -0.515 125.285 ;
        RECT -0.845 123.595 -0.515 123.925 ;
        RECT -0.845 122.215 -0.515 122.545 ;
        RECT -0.845 120.165 -0.515 120.495 ;
        RECT -0.845 118.235 -0.515 118.565 ;
        RECT -0.845 116.395 -0.515 116.725 ;
        RECT -0.845 114.905 -0.515 115.235 ;
        RECT -0.845 113.235 -0.515 113.565 ;
        RECT -0.845 111.745 -0.515 112.075 ;
        RECT -0.845 110.075 -0.515 110.405 ;
        RECT -0.845 108.585 -0.515 108.915 ;
        RECT -0.845 106.915 -0.515 107.245 ;
        RECT -0.845 105.425 -0.515 105.755 ;
        RECT -0.845 104.015 -0.515 104.345 ;
        RECT -0.845 102.175 -0.515 102.505 ;
        RECT -0.845 100.685 -0.515 101.015 ;
        RECT -0.845 99.015 -0.515 99.345 ;
        RECT -0.845 97.525 -0.515 97.855 ;
        RECT -0.845 95.855 -0.515 96.185 ;
        RECT -0.845 94.365 -0.515 94.695 ;
        RECT -0.845 92.695 -0.515 93.025 ;
        RECT -0.845 91.205 -0.515 91.535 ;
        RECT -0.845 89.795 -0.515 90.125 ;
        RECT -0.845 87.955 -0.515 88.285 ;
        RECT -0.845 86.465 -0.515 86.795 ;
        RECT -0.845 84.795 -0.515 85.125 ;
        RECT -0.845 83.305 -0.515 83.635 ;
        RECT -0.845 81.635 -0.515 81.965 ;
        RECT -0.845 80.145 -0.515 80.475 ;
        RECT -0.845 78.475 -0.515 78.805 ;
        RECT -0.845 76.985 -0.515 77.315 ;
        RECT -0.845 75.575 -0.515 75.905 ;
        RECT -0.845 73.735 -0.515 74.065 ;
        RECT -0.845 72.245 -0.515 72.575 ;
        RECT -0.845 70.575 -0.515 70.905 ;
        RECT -0.845 69.085 -0.515 69.415 ;
        RECT -0.845 67.415 -0.515 67.745 ;
        RECT -0.845 65.925 -0.515 66.255 ;
        RECT -0.845 64.255 -0.515 64.585 ;
        RECT -0.845 62.765 -0.515 63.095 ;
        RECT -0.845 61.355 -0.515 61.685 ;
        RECT -0.845 59.515 -0.515 59.845 ;
        RECT -0.845 58.025 -0.515 58.355 ;
        RECT -0.845 56.355 -0.515 56.685 ;
        RECT -0.845 54.865 -0.515 55.195 ;
        RECT -0.845 53.195 -0.515 53.525 ;
        RECT -0.845 51.705 -0.515 52.035 ;
        RECT -0.845 50.035 -0.515 50.365 ;
        RECT -0.845 48.545 -0.515 48.875 ;
        RECT -0.845 47.135 -0.515 47.465 ;
        RECT -0.845 45.295 -0.515 45.625 ;
        RECT -0.845 43.805 -0.515 44.135 ;
        RECT -0.845 42.135 -0.515 42.465 ;
        RECT -0.845 40.645 -0.515 40.975 ;
        RECT -0.845 38.975 -0.515 39.305 ;
        RECT -0.845 37.485 -0.515 37.815 ;
        RECT -0.845 35.815 -0.515 36.145 ;
        RECT -0.845 34.325 -0.515 34.655 ;
        RECT -0.845 32.915 -0.515 33.245 ;
        RECT -0.845 31.075 -0.515 31.405 ;
        RECT -0.845 29.585 -0.515 29.915 ;
        RECT -0.845 27.915 -0.515 28.245 ;
        RECT -0.845 26.425 -0.515 26.755 ;
        RECT -0.845 24.755 -0.515 25.085 ;
        RECT -0.845 23.265 -0.515 23.595 ;
        RECT -0.845 21.595 -0.515 21.925 ;
        RECT -0.845 20.105 -0.515 20.435 ;
        RECT -0.845 18.695 -0.515 19.025 ;
        RECT -0.845 16.855 -0.515 17.185 ;
        RECT -0.845 15.365 -0.515 15.695 ;
        RECT -0.845 13.695 -0.515 14.025 ;
        RECT -0.845 12.205 -0.515 12.535 ;
        RECT -0.845 10.535 -0.515 10.865 ;
        RECT -0.845 9.045 -0.515 9.375 ;
        RECT -0.845 7.375 -0.515 7.705 ;
        RECT -0.845 5.885 -0.515 6.215 ;
        RECT -0.845 4.475 -0.515 4.805 ;
        RECT -0.845 2.115 -0.515 2.445 ;
        RECT -0.845 0.06 -0.515 0.39 ;
        RECT -0.845 -1.525 -0.515 -1.195 ;
        RECT -0.845 -2.885 -0.515 -2.555 ;
        RECT -0.845 -4.245 -0.515 -3.915 ;
        RECT -0.845 -5.605 -0.515 -5.275 ;
        RECT -0.845 -6.965 -0.515 -6.635 ;
        RECT -0.845 -8.325 -0.515 -7.995 ;
        RECT -0.845 -9.685 -0.515 -9.355 ;
        RECT -0.845 -12.405 -0.515 -12.075 ;
        RECT -0.845 -13.765 -0.515 -13.435 ;
        RECT -0.845 -15.125 -0.515 -14.795 ;
        RECT -0.845 -16.485 -0.515 -16.155 ;
        RECT -0.845 -17.845 -0.515 -17.515 ;
        RECT -0.845 -19.205 -0.515 -18.875 ;
        RECT -0.845 -20.565 -0.515 -20.235 ;
        RECT -0.845 -21.925 -0.515 -21.595 ;
        RECT -0.845 -23.285 -0.515 -22.955 ;
        RECT -0.845 -24.645 -0.515 -24.315 ;
        RECT -0.845 -26.005 -0.515 -25.675 ;
        RECT -0.845 -27.365 -0.515 -27.035 ;
        RECT -0.845 -28.725 -0.515 -28.395 ;
        RECT -0.845 -30.085 -0.515 -29.755 ;
        RECT -0.845 -31.445 -0.515 -31.115 ;
        RECT -0.845 -32.805 -0.515 -32.475 ;
        RECT -0.845 -34.165 -0.515 -33.835 ;
        RECT -0.845 -35.525 -0.515 -35.195 ;
        RECT -0.845 -36.885 -0.515 -36.555 ;
        RECT -0.845 -38.245 -0.515 -37.915 ;
        RECT -0.845 -39.605 -0.515 -39.275 ;
        RECT -0.845 -40.965 -0.515 -40.635 ;
        RECT -0.845 -42.325 -0.515 -41.995 ;
        RECT -0.845 -43.685 -0.515 -43.355 ;
        RECT -0.845 -45.045 -0.515 -44.715 ;
        RECT -0.845 -46.405 -0.515 -46.075 ;
        RECT -0.845 -47.765 -0.515 -47.435 ;
        RECT -0.845 -49.125 -0.515 -48.795 ;
        RECT -0.845 -50.485 -0.515 -50.155 ;
        RECT -0.845 -51.845 -0.515 -51.515 ;
        RECT -0.845 -53.205 -0.515 -52.875 ;
        RECT -0.845 -54.565 -0.515 -54.235 ;
        RECT -0.845 -55.925 -0.515 -55.595 ;
        RECT -0.845 -57.285 -0.515 -56.955 ;
        RECT -0.845 -58.645 -0.515 -58.315 ;
        RECT -0.845 -61.365 -0.515 -61.035 ;
        RECT -0.845 -65.445 -0.515 -65.115 ;
        RECT -0.845 -66.805 -0.515 -66.475 ;
        RECT -0.845 -68.165 -0.515 -67.835 ;
        RECT -0.845 -69.525 -0.515 -69.195 ;
        RECT -0.845 -70.885 -0.515 -70.555 ;
        RECT -0.845 -72.245 -0.515 -71.915 ;
        RECT -0.845 -73.605 -0.515 -73.275 ;
        RECT -0.845 -74.965 -0.515 -74.635 ;
        RECT -0.845 -76.325 -0.515 -75.995 ;
        RECT -0.845 -77.685 -0.515 -77.355 ;
        RECT -0.845 -79.045 -0.515 -78.715 ;
        RECT -0.845 -80.405 -0.515 -80.075 ;
        RECT -0.845 -81.765 -0.515 -81.435 ;
        RECT -0.845 -83.125 -0.515 -82.795 ;
        RECT -0.845 -84.485 -0.515 -84.155 ;
        RECT -0.845 -85.845 -0.515 -85.515 ;
    END
    PORT
      LAYER met3 ;
        RECT -14.445 -210.965 -14.115 -210.635 ;
        RECT -14.445 -212.325 -14.115 -211.995 ;
        RECT -14.445 -213.625 -14.115 -213.295 ;
        RECT -14.445 -215.045 -14.115 -214.715 ;
        RECT -14.445 -216.405 -14.115 -216.075 ;
        RECT -14.445 -217.765 -14.115 -217.435 ;
        RECT -14.445 -219.125 -14.115 -218.795 ;
        RECT -14.445 -221.37 -14.115 -220.24 ;
        RECT -14.44 -221.485 -14.12 -209.28 ;
    END
    PORT
      LAYER met3 ;
        RECT -13.085 129.8 -12.755 130.93 ;
        RECT -13.085 127.675 -12.755 128.005 ;
        RECT -13.085 126.315 -12.755 126.645 ;
        RECT -13.085 124.955 -12.755 125.285 ;
        RECT -13.085 123.595 -12.755 123.925 ;
        RECT -13.085 122.235 -12.755 122.565 ;
        RECT -13.085 120.875 -12.755 121.205 ;
        RECT -13.085 119.515 -12.755 119.845 ;
        RECT -13.085 118.155 -12.755 118.485 ;
        RECT -13.085 116.795 -12.755 117.125 ;
        RECT -13.085 115.435 -12.755 115.765 ;
        RECT -13.085 114.075 -12.755 114.405 ;
        RECT -13.085 112.715 -12.755 113.045 ;
        RECT -13.085 111.355 -12.755 111.685 ;
        RECT -13.085 109.995 -12.755 110.325 ;
        RECT -13.085 108.635 -12.755 108.965 ;
        RECT -13.085 107.275 -12.755 107.605 ;
        RECT -13.085 105.915 -12.755 106.245 ;
        RECT -13.085 104.555 -12.755 104.885 ;
        RECT -13.085 103.195 -12.755 103.525 ;
        RECT -13.085 101.835 -12.755 102.165 ;
        RECT -13.085 100.475 -12.755 100.805 ;
        RECT -13.085 99.115 -12.755 99.445 ;
        RECT -13.085 97.755 -12.755 98.085 ;
        RECT -13.085 96.395 -12.755 96.725 ;
        RECT -13.085 95.035 -12.755 95.365 ;
        RECT -13.085 93.675 -12.755 94.005 ;
        RECT -13.085 92.315 -12.755 92.645 ;
        RECT -13.085 90.955 -12.755 91.285 ;
        RECT -13.085 89.595 -12.755 89.925 ;
        RECT -13.085 88.235 -12.755 88.565 ;
        RECT -13.085 86.875 -12.755 87.205 ;
        RECT -13.085 85.515 -12.755 85.845 ;
        RECT -13.085 84.155 -12.755 84.485 ;
        RECT -13.085 82.795 -12.755 83.125 ;
        RECT -13.085 81.435 -12.755 81.765 ;
        RECT -13.085 80.075 -12.755 80.405 ;
        RECT -13.085 78.715 -12.755 79.045 ;
        RECT -13.085 77.355 -12.755 77.685 ;
        RECT -13.085 75.995 -12.755 76.325 ;
        RECT -13.085 74.635 -12.755 74.965 ;
        RECT -13.085 73.275 -12.755 73.605 ;
        RECT -13.085 71.915 -12.755 72.245 ;
        RECT -13.085 70.555 -12.755 70.885 ;
        RECT -13.085 69.195 -12.755 69.525 ;
        RECT -13.085 67.835 -12.755 68.165 ;
        RECT -13.085 66.475 -12.755 66.805 ;
        RECT -13.085 65.115 -12.755 65.445 ;
        RECT -13.085 63.755 -12.755 64.085 ;
        RECT -13.085 62.395 -12.755 62.725 ;
        RECT -13.085 61.035 -12.755 61.365 ;
        RECT -13.085 59.675 -12.755 60.005 ;
        RECT -13.085 58.315 -12.755 58.645 ;
        RECT -13.085 56.955 -12.755 57.285 ;
        RECT -13.085 55.595 -12.755 55.925 ;
        RECT -13.085 54.235 -12.755 54.565 ;
        RECT -13.085 52.875 -12.755 53.205 ;
        RECT -13.085 51.515 -12.755 51.845 ;
        RECT -13.085 50.155 -12.755 50.485 ;
        RECT -13.085 48.795 -12.755 49.125 ;
        RECT -13.085 47.435 -12.755 47.765 ;
        RECT -13.085 46.075 -12.755 46.405 ;
        RECT -13.085 44.715 -12.755 45.045 ;
        RECT -13.085 43.355 -12.755 43.685 ;
        RECT -13.085 41.995 -12.755 42.325 ;
        RECT -13.085 40.635 -12.755 40.965 ;
        RECT -13.085 39.275 -12.755 39.605 ;
        RECT -13.085 37.915 -12.755 38.245 ;
        RECT -13.085 36.555 -12.755 36.885 ;
        RECT -13.085 35.195 -12.755 35.525 ;
        RECT -13.085 33.835 -12.755 34.165 ;
        RECT -13.085 32.475 -12.755 32.805 ;
        RECT -13.085 31.115 -12.755 31.445 ;
        RECT -13.085 29.755 -12.755 30.085 ;
        RECT -13.085 28.395 -12.755 28.725 ;
        RECT -13.085 27.035 -12.755 27.365 ;
        RECT -13.085 25.675 -12.755 26.005 ;
        RECT -13.085 24.315 -12.755 24.645 ;
        RECT -13.085 22.955 -12.755 23.285 ;
        RECT -13.085 21.595 -12.755 21.925 ;
        RECT -13.085 20.235 -12.755 20.565 ;
        RECT -13.085 18.875 -12.755 19.205 ;
        RECT -13.085 17.515 -12.755 17.845 ;
        RECT -13.085 16.155 -12.755 16.485 ;
        RECT -13.085 14.795 -12.755 15.125 ;
        RECT -13.085 13.435 -12.755 13.765 ;
        RECT -13.085 12.075 -12.755 12.405 ;
        RECT -13.085 10.715 -12.755 11.045 ;
        RECT -13.085 9.355 -12.755 9.685 ;
        RECT -13.085 7.995 -12.755 8.325 ;
        RECT -13.085 6.635 -12.755 6.965 ;
        RECT -13.085 5.275 -12.755 5.605 ;
        RECT -13.085 3.915 -12.755 4.245 ;
        RECT -13.085 2.555 -12.755 2.885 ;
        RECT -13.085 1.195 -12.755 1.525 ;
        RECT -13.085 -0.165 -12.755 0.165 ;
        RECT -13.085 -1.525 -12.755 -1.195 ;
        RECT -13.085 -2.885 -12.755 -2.555 ;
        RECT -13.085 -4.245 -12.755 -3.915 ;
        RECT -13.085 -8.325 -12.755 -7.995 ;
        RECT -13.085 -9.685 -12.755 -9.355 ;
        RECT -13.085 -11.16 -12.755 -10.83 ;
        RECT -13.085 -12.405 -12.755 -12.075 ;
        RECT -13.085 -15.125 -12.755 -14.795 ;
        RECT -13.085 -16.25 -12.755 -15.92 ;
        RECT -13.085 -21.925 -12.755 -21.595 ;
        RECT -13.085 -23.285 -12.755 -22.955 ;
        RECT -13.085 -24.645 -12.755 -24.315 ;
        RECT -13.085 -27.365 -12.755 -27.035 ;
        RECT -13.085 -30.085 -12.755 -29.755 ;
        RECT -13.085 -31.445 -12.755 -31.115 ;
        RECT -13.085 -32.34 -12.755 -32.01 ;
        RECT -13.085 -34.165 -12.755 -33.835 ;
        RECT -13.085 -37.43 -12.755 -37.1 ;
        RECT -13.085 -38.245 -12.755 -37.915 ;
        RECT -13.085 -43.685 -12.755 -43.355 ;
        RECT -13.085 -45.045 -12.755 -44.715 ;
        RECT -13.085 -46.405 -12.755 -46.075 ;
        RECT -13.085 -47.765 -12.755 -47.435 ;
        RECT -13.085 -49.125 -12.755 -48.795 ;
        RECT -13.085 -50.485 -12.755 -50.155 ;
        RECT -13.085 -53.205 -12.755 -52.875 ;
        RECT -13.085 -54.565 -12.755 -54.235 ;
        RECT -13.085 -55.925 -12.755 -55.595 ;
        RECT -13.085 -57.285 -12.755 -56.955 ;
        RECT -13.085 -58.645 -12.755 -58.315 ;
        RECT -13.085 -60.005 -12.755 -59.675 ;
        RECT -13.085 -61.67 -12.755 -61.34 ;
        RECT -13.085 -65.445 -12.755 -65.115 ;
        RECT -13.085 -66.805 -12.755 -66.475 ;
        RECT -13.085 -68.165 -12.755 -67.835 ;
        RECT -13.085 -69.525 -12.755 -69.195 ;
        RECT -13.085 -72.245 -12.755 -71.915 ;
        RECT -13.085 -73.605 -12.755 -73.275 ;
        RECT -13.085 -74.965 -12.755 -74.635 ;
        RECT -13.085 -76.325 -12.755 -75.995 ;
        RECT -13.085 -77.685 -12.755 -77.355 ;
        RECT -13.085 -79.045 -12.755 -78.715 ;
        RECT -13.085 -80.21 -12.755 -79.88 ;
        RECT -13.085 -81.765 -12.755 -81.435 ;
        RECT -13.085 -83.125 -12.755 -82.795 ;
        RECT -13.085 -84.485 -12.755 -84.155 ;
        RECT -13.085 -87.205 -12.755 -86.875 ;
        RECT -13.085 -88.565 -12.755 -88.235 ;
        RECT -13.085 -89.925 -12.755 -89.595 ;
        RECT -13.085 -91.285 -12.755 -90.955 ;
        RECT -13.085 -92.645 -12.755 -92.315 ;
        RECT -13.085 -94.005 -12.755 -93.675 ;
        RECT -13.085 -95.365 -12.755 -95.035 ;
        RECT -13.085 -98.085 -12.755 -97.755 ;
        RECT -13.085 -99.445 -12.755 -99.115 ;
        RECT -13.085 -100.805 -12.755 -100.475 ;
        RECT -13.085 -102.165 -12.755 -101.835 ;
        RECT -13.085 -103.525 -12.755 -103.195 ;
        RECT -13.085 -104.885 -12.755 -104.555 ;
        RECT -13.085 -105.85 -12.755 -105.52 ;
        RECT -13.085 -107.605 -12.755 -107.275 ;
        RECT -13.085 -108.965 -12.755 -108.635 ;
        RECT -13.085 -110.325 -12.755 -109.995 ;
        RECT -13.085 -111.685 -12.755 -111.355 ;
        RECT -13.085 -115.765 -12.755 -115.435 ;
        RECT -13.085 -117.125 -12.755 -116.795 ;
        RECT -13.085 -118.485 -12.755 -118.155 ;
        RECT -13.085 -119.845 -12.755 -119.515 ;
        RECT -13.085 -121.205 -12.755 -120.875 ;
        RECT -13.085 -122.565 -12.755 -122.235 ;
        RECT -13.085 -124.39 -12.755 -124.06 ;
        RECT -13.085 -125.285 -12.755 -124.955 ;
        RECT -13.085 -126.645 -12.755 -126.315 ;
        RECT -13.085 -128.005 -12.755 -127.675 ;
        RECT -13.085 -129.365 -12.755 -129.035 ;
        RECT -13.085 -133.445 -12.755 -133.115 ;
        RECT -13.085 -134.805 -12.755 -134.475 ;
        RECT -13.085 -136.165 -12.755 -135.835 ;
        RECT -13.085 -137.525 -12.755 -137.195 ;
        RECT -13.085 -138.885 -12.755 -138.555 ;
        RECT -13.085 -140.245 -12.755 -139.915 ;
        RECT -13.085 -144.325 -12.755 -143.995 ;
        RECT -13.085 -148.405 -12.755 -148.075 ;
        RECT -13.085 -152.485 -12.755 -152.155 ;
        RECT -13.085 -155.205 -12.755 -154.875 ;
        RECT -13.085 -156.565 -12.755 -156.235 ;
        RECT -13.085 -157.925 -12.755 -157.595 ;
        RECT -13.085 -159.285 -12.755 -158.955 ;
        RECT -13.085 -160.645 -12.755 -160.315 ;
        RECT -13.085 -162.005 -12.755 -161.675 ;
        RECT -13.085 -163.365 -12.755 -163.035 ;
        RECT -13.085 -166.085 -12.755 -165.755 ;
        RECT -13.085 -168.805 -12.755 -168.475 ;
        RECT -13.085 -170.165 -12.755 -169.835 ;
        RECT -13.085 -171.525 -12.755 -171.195 ;
        RECT -13.085 -174.245 -12.755 -173.915 ;
        RECT -13.085 -175.605 -12.755 -175.275 ;
        RECT -13.085 -176.965 -12.755 -176.635 ;
        RECT -13.085 -178.325 -12.755 -177.995 ;
        RECT -13.085 -179.685 -12.755 -179.355 ;
        RECT -13.085 -183.765 -12.755 -183.435 ;
        RECT -13.085 -185.125 -12.755 -184.795 ;
        RECT -13.085 -187.845 -12.755 -187.515 ;
        RECT -13.085 -191.925 -12.755 -191.595 ;
        RECT -13.085 -194.645 -12.755 -194.315 ;
        RECT -13.085 -196.005 -12.755 -195.675 ;
        RECT -13.085 -197.365 -12.755 -197.035 ;
        RECT -13.085 -198.725 -12.755 -198.395 ;
        RECT -13.085 -200.085 -12.755 -199.755 ;
        RECT -13.085 -201.445 -12.755 -201.115 ;
        RECT -13.085 -202.805 -12.755 -202.475 ;
        RECT -13.085 -204.165 -12.755 -203.835 ;
        RECT -13.085 -208.245 -12.755 -207.915 ;
        RECT -13.085 -210.965 -12.755 -210.635 ;
        RECT -13.085 -212.325 -12.755 -211.995 ;
        RECT -13.085 -213.625 -12.755 -213.295 ;
        RECT -13.085 -215.045 -12.755 -214.715 ;
        RECT -13.085 -216.405 -12.755 -216.075 ;
        RECT -13.085 -217.765 -12.755 -217.435 ;
        RECT -13.085 -219.125 -12.755 -218.795 ;
        RECT -13.085 -221.37 -12.755 -220.24 ;
        RECT -13.08 -221.485 -12.76 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.725 129.8 -11.395 130.93 ;
        RECT -11.725 127.675 -11.395 128.005 ;
        RECT -11.725 126.315 -11.395 126.645 ;
        RECT -11.725 124.955 -11.395 125.285 ;
        RECT -11.725 123.595 -11.395 123.925 ;
        RECT -11.725 122.235 -11.395 122.565 ;
        RECT -11.725 120.875 -11.395 121.205 ;
        RECT -11.725 119.515 -11.395 119.845 ;
        RECT -11.725 118.155 -11.395 118.485 ;
        RECT -11.725 116.795 -11.395 117.125 ;
        RECT -11.725 115.435 -11.395 115.765 ;
        RECT -11.725 114.075 -11.395 114.405 ;
        RECT -11.725 112.715 -11.395 113.045 ;
        RECT -11.725 111.355 -11.395 111.685 ;
        RECT -11.725 109.995 -11.395 110.325 ;
        RECT -11.725 108.635 -11.395 108.965 ;
        RECT -11.725 107.275 -11.395 107.605 ;
        RECT -11.725 105.915 -11.395 106.245 ;
        RECT -11.725 104.555 -11.395 104.885 ;
        RECT -11.725 103.195 -11.395 103.525 ;
        RECT -11.725 101.835 -11.395 102.165 ;
        RECT -11.725 100.475 -11.395 100.805 ;
        RECT -11.725 99.115 -11.395 99.445 ;
        RECT -11.725 97.755 -11.395 98.085 ;
        RECT -11.725 96.395 -11.395 96.725 ;
        RECT -11.725 95.035 -11.395 95.365 ;
        RECT -11.725 93.675 -11.395 94.005 ;
        RECT -11.725 92.315 -11.395 92.645 ;
        RECT -11.725 90.955 -11.395 91.285 ;
        RECT -11.725 89.595 -11.395 89.925 ;
        RECT -11.725 88.235 -11.395 88.565 ;
        RECT -11.725 86.875 -11.395 87.205 ;
        RECT -11.725 85.515 -11.395 85.845 ;
        RECT -11.725 84.155 -11.395 84.485 ;
        RECT -11.725 82.795 -11.395 83.125 ;
        RECT -11.725 81.435 -11.395 81.765 ;
        RECT -11.725 80.075 -11.395 80.405 ;
        RECT -11.725 78.715 -11.395 79.045 ;
        RECT -11.725 77.355 -11.395 77.685 ;
        RECT -11.725 75.995 -11.395 76.325 ;
        RECT -11.725 74.635 -11.395 74.965 ;
        RECT -11.725 73.275 -11.395 73.605 ;
        RECT -11.725 71.915 -11.395 72.245 ;
        RECT -11.725 70.555 -11.395 70.885 ;
        RECT -11.725 69.195 -11.395 69.525 ;
        RECT -11.725 67.835 -11.395 68.165 ;
        RECT -11.725 66.475 -11.395 66.805 ;
        RECT -11.725 65.115 -11.395 65.445 ;
        RECT -11.725 63.755 -11.395 64.085 ;
        RECT -11.725 62.395 -11.395 62.725 ;
        RECT -11.725 61.035 -11.395 61.365 ;
        RECT -11.725 59.675 -11.395 60.005 ;
        RECT -11.725 58.315 -11.395 58.645 ;
        RECT -11.725 56.955 -11.395 57.285 ;
        RECT -11.725 55.595 -11.395 55.925 ;
        RECT -11.725 54.235 -11.395 54.565 ;
        RECT -11.725 52.875 -11.395 53.205 ;
        RECT -11.725 51.515 -11.395 51.845 ;
        RECT -11.725 50.155 -11.395 50.485 ;
        RECT -11.725 48.795 -11.395 49.125 ;
        RECT -11.725 47.435 -11.395 47.765 ;
        RECT -11.725 46.075 -11.395 46.405 ;
        RECT -11.725 44.715 -11.395 45.045 ;
        RECT -11.725 43.355 -11.395 43.685 ;
        RECT -11.725 41.995 -11.395 42.325 ;
        RECT -11.725 40.635 -11.395 40.965 ;
        RECT -11.725 39.275 -11.395 39.605 ;
        RECT -11.725 37.915 -11.395 38.245 ;
        RECT -11.725 36.555 -11.395 36.885 ;
        RECT -11.725 35.195 -11.395 35.525 ;
        RECT -11.725 33.835 -11.395 34.165 ;
        RECT -11.725 32.475 -11.395 32.805 ;
        RECT -11.725 31.115 -11.395 31.445 ;
        RECT -11.725 29.755 -11.395 30.085 ;
        RECT -11.725 28.395 -11.395 28.725 ;
        RECT -11.725 27.035 -11.395 27.365 ;
        RECT -11.725 25.675 -11.395 26.005 ;
        RECT -11.725 24.315 -11.395 24.645 ;
        RECT -11.725 22.955 -11.395 23.285 ;
        RECT -11.725 21.595 -11.395 21.925 ;
        RECT -11.725 20.235 -11.395 20.565 ;
        RECT -11.725 18.875 -11.395 19.205 ;
        RECT -11.725 17.515 -11.395 17.845 ;
        RECT -11.725 16.155 -11.395 16.485 ;
        RECT -11.725 14.795 -11.395 15.125 ;
        RECT -11.725 13.435 -11.395 13.765 ;
        RECT -11.725 12.075 -11.395 12.405 ;
        RECT -11.725 10.715 -11.395 11.045 ;
        RECT -11.725 9.355 -11.395 9.685 ;
        RECT -11.725 7.995 -11.395 8.325 ;
        RECT -11.725 6.635 -11.395 6.965 ;
        RECT -11.725 5.275 -11.395 5.605 ;
        RECT -11.725 3.915 -11.395 4.245 ;
        RECT -11.725 2.555 -11.395 2.885 ;
        RECT -11.725 1.195 -11.395 1.525 ;
        RECT -11.725 -0.165 -11.395 0.165 ;
        RECT -11.725 -1.525 -11.395 -1.195 ;
        RECT -11.725 -2.885 -11.395 -2.555 ;
        RECT -11.725 -4.245 -11.395 -3.915 ;
        RECT -11.725 -5.605 -11.395 -5.275 ;
        RECT -11.725 -8.325 -11.395 -7.995 ;
        RECT -11.725 -9.685 -11.395 -9.355 ;
        RECT -11.725 -11.16 -11.395 -10.83 ;
        RECT -11.725 -12.405 -11.395 -12.075 ;
        RECT -11.725 -15.125 -11.395 -14.795 ;
        RECT -11.725 -16.25 -11.395 -15.92 ;
        RECT -11.725 -21.925 -11.395 -21.595 ;
        RECT -11.725 -23.285 -11.395 -22.955 ;
        RECT -11.725 -24.645 -11.395 -24.315 ;
        RECT -11.725 -26.005 -11.395 -25.675 ;
        RECT -11.725 -27.365 -11.395 -27.035 ;
        RECT -11.725 -30.085 -11.395 -29.755 ;
        RECT -11.725 -31.445 -11.395 -31.115 ;
        RECT -11.725 -32.34 -11.395 -32.01 ;
        RECT -11.725 -34.165 -11.395 -33.835 ;
        RECT -11.725 -37.43 -11.395 -37.1 ;
        RECT -11.725 -38.245 -11.395 -37.915 ;
        RECT -11.725 -43.685 -11.395 -43.355 ;
        RECT -11.725 -45.045 -11.395 -44.715 ;
        RECT -11.725 -46.405 -11.395 -46.075 ;
        RECT -11.725 -47.765 -11.395 -47.435 ;
        RECT -11.725 -49.125 -11.395 -48.795 ;
        RECT -11.725 -50.485 -11.395 -50.155 ;
        RECT -11.725 -53.205 -11.395 -52.875 ;
        RECT -11.725 -54.565 -11.395 -54.235 ;
        RECT -11.725 -55.925 -11.395 -55.595 ;
        RECT -11.725 -57.285 -11.395 -56.955 ;
        RECT -11.725 -58.645 -11.395 -58.315 ;
        RECT -11.725 -61.67 -11.395 -61.34 ;
        RECT -11.725 -65.445 -11.395 -65.115 ;
        RECT -11.725 -66.805 -11.395 -66.475 ;
        RECT -11.725 -68.165 -11.395 -67.835 ;
        RECT -11.725 -69.525 -11.395 -69.195 ;
        RECT -11.725 -72.245 -11.395 -71.915 ;
        RECT -11.725 -73.605 -11.395 -73.275 ;
        RECT -11.725 -74.965 -11.395 -74.635 ;
        RECT -11.725 -76.325 -11.395 -75.995 ;
        RECT -11.725 -77.685 -11.395 -77.355 ;
        RECT -11.725 -79.045 -11.395 -78.715 ;
        RECT -11.725 -80.21 -11.395 -79.88 ;
        RECT -11.725 -81.765 -11.395 -81.435 ;
        RECT -11.725 -83.125 -11.395 -82.795 ;
        RECT -11.725 -84.485 -11.395 -84.155 ;
        RECT -11.725 -87.205 -11.395 -86.875 ;
        RECT -11.725 -88.565 -11.395 -88.235 ;
        RECT -11.725 -89.925 -11.395 -89.595 ;
        RECT -11.725 -91.285 -11.395 -90.955 ;
        RECT -11.725 -92.645 -11.395 -92.315 ;
        RECT -11.725 -94.005 -11.395 -93.675 ;
        RECT -11.725 -95.365 -11.395 -95.035 ;
        RECT -11.725 -98.085 -11.395 -97.755 ;
        RECT -11.725 -99.445 -11.395 -99.115 ;
        RECT -11.725 -100.805 -11.395 -100.475 ;
        RECT -11.725 -102.165 -11.395 -101.835 ;
        RECT -11.725 -103.525 -11.395 -103.195 ;
        RECT -11.725 -104.885 -11.395 -104.555 ;
        RECT -11.725 -105.85 -11.395 -105.52 ;
        RECT -11.725 -107.605 -11.395 -107.275 ;
        RECT -11.725 -108.965 -11.395 -108.635 ;
        RECT -11.725 -110.325 -11.395 -109.995 ;
        RECT -11.725 -111.685 -11.395 -111.355 ;
        RECT -11.725 -115.765 -11.395 -115.435 ;
        RECT -11.725 -117.125 -11.395 -116.795 ;
        RECT -11.725 -118.485 -11.395 -118.155 ;
        RECT -11.725 -119.845 -11.395 -119.515 ;
        RECT -11.725 -121.205 -11.395 -120.875 ;
        RECT -11.725 -122.565 -11.395 -122.235 ;
        RECT -11.725 -124.39 -11.395 -124.06 ;
        RECT -11.725 -125.285 -11.395 -124.955 ;
        RECT -11.725 -126.645 -11.395 -126.315 ;
        RECT -11.725 -128.005 -11.395 -127.675 ;
        RECT -11.725 -129.365 -11.395 -129.035 ;
        RECT -11.725 -133.445 -11.395 -133.115 ;
        RECT -11.725 -134.805 -11.395 -134.475 ;
        RECT -11.725 -136.165 -11.395 -135.835 ;
        RECT -11.725 -137.525 -11.395 -137.195 ;
        RECT -11.725 -138.885 -11.395 -138.555 ;
        RECT -11.725 -140.245 -11.395 -139.915 ;
        RECT -11.725 -144.325 -11.395 -143.995 ;
        RECT -11.725 -148.405 -11.395 -148.075 ;
        RECT -11.725 -152.485 -11.395 -152.155 ;
        RECT -11.725 -153.845 -11.395 -153.515 ;
        RECT -11.725 -155.205 -11.395 -154.875 ;
        RECT -11.725 -156.565 -11.395 -156.235 ;
        RECT -11.725 -157.925 -11.395 -157.595 ;
        RECT -11.725 -159.285 -11.395 -158.955 ;
        RECT -11.725 -160.645 -11.395 -160.315 ;
        RECT -11.725 -162.005 -11.395 -161.675 ;
        RECT -11.725 -163.365 -11.395 -163.035 ;
        RECT -11.725 -164.725 -11.395 -164.395 ;
        RECT -11.725 -166.085 -11.395 -165.755 ;
        RECT -11.725 -168.805 -11.395 -168.475 ;
        RECT -11.725 -170.165 -11.395 -169.835 ;
        RECT -11.725 -171.525 -11.395 -171.195 ;
        RECT -11.725 -172.885 -11.395 -172.555 ;
        RECT -11.725 -174.245 -11.395 -173.915 ;
        RECT -11.725 -175.605 -11.395 -175.275 ;
        RECT -11.725 -176.965 -11.395 -176.635 ;
        RECT -11.725 -178.325 -11.395 -177.995 ;
        RECT -11.725 -179.685 -11.395 -179.355 ;
        RECT -11.725 -183.765 -11.395 -183.435 ;
        RECT -11.725 -185.125 -11.395 -184.795 ;
        RECT -11.725 -186.485 -11.395 -186.155 ;
        RECT -11.725 -187.845 -11.395 -187.515 ;
        RECT -11.725 -189.205 -11.395 -188.875 ;
        RECT -11.725 -190.565 -11.395 -190.235 ;
        RECT -11.725 -191.925 -11.395 -191.595 ;
        RECT -11.725 -193.285 -11.395 -192.955 ;
        RECT -11.725 -194.645 -11.395 -194.315 ;
        RECT -11.725 -196.005 -11.395 -195.675 ;
        RECT -11.725 -197.365 -11.395 -197.035 ;
        RECT -11.725 -198.725 -11.395 -198.395 ;
        RECT -11.725 -200.085 -11.395 -199.755 ;
        RECT -11.725 -201.445 -11.395 -201.115 ;
        RECT -11.725 -202.805 -11.395 -202.475 ;
        RECT -11.725 -204.165 -11.395 -203.835 ;
        RECT -11.725 -208.245 -11.395 -207.915 ;
        RECT -11.725 -210.965 -11.395 -210.635 ;
        RECT -11.725 -212.325 -11.395 -211.995 ;
        RECT -11.725 -213.625 -11.395 -213.295 ;
        RECT -11.725 -215.045 -11.395 -214.715 ;
        RECT -11.725 -216.405 -11.395 -216.075 ;
        RECT -11.725 -217.765 -11.395 -217.435 ;
        RECT -11.725 -219.125 -11.395 -218.795 ;
        RECT -11.725 -221.37 -11.395 -220.24 ;
        RECT -11.72 -221.485 -11.4 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -10.365 129.8 -10.035 130.93 ;
        RECT -10.365 127.675 -10.035 128.005 ;
        RECT -10.365 126.315 -10.035 126.645 ;
        RECT -10.365 124.955 -10.035 125.285 ;
        RECT -10.365 123.595 -10.035 123.925 ;
        RECT -10.365 122.235 -10.035 122.565 ;
        RECT -10.365 120.875 -10.035 121.205 ;
        RECT -10.365 119.515 -10.035 119.845 ;
        RECT -10.365 118.155 -10.035 118.485 ;
        RECT -10.365 114.075 -10.035 114.405 ;
        RECT -10.365 104.555 -10.035 104.885 ;
        RECT -10.365 103.195 -10.035 103.525 ;
        RECT -10.365 96.395 -10.035 96.725 ;
        RECT -10.365 93.675 -10.035 94.005 ;
        RECT -10.365 89.595 -10.035 89.925 ;
        RECT -10.365 85.515 -10.035 85.845 ;
        RECT -10.365 82.795 -10.035 83.125 ;
        RECT -10.365 75.995 -10.035 76.325 ;
        RECT -10.365 74.635 -10.035 74.965 ;
        RECT -10.365 65.115 -10.035 65.445 ;
        RECT -10.365 61.035 -10.035 61.365 ;
        RECT -10.365 56.955 -10.035 57.285 ;
        RECT -10.365 54.235 -10.035 54.565 ;
        RECT -10.365 47.435 -10.035 47.765 ;
        RECT -10.365 46.075 -10.035 46.405 ;
        RECT -10.365 43.355 -10.035 43.685 ;
        RECT -10.365 36.555 -10.035 36.885 ;
        RECT -10.365 33.835 -10.035 34.165 ;
        RECT -10.365 32.475 -10.035 32.805 ;
        RECT -10.365 28.395 -10.035 28.725 ;
        RECT -10.365 25.675 -10.035 26.005 ;
        RECT -10.365 18.875 -10.035 19.205 ;
        RECT -10.365 17.515 -10.035 17.845 ;
        RECT -10.365 14.795 -10.035 15.125 ;
        RECT -10.365 7.995 -10.035 8.325 ;
        RECT -10.365 5.275 -10.035 5.605 ;
        RECT -10.365 3.915 -10.035 4.245 ;
        RECT -10.365 2.555 -10.035 2.885 ;
        RECT -10.365 1.195 -10.035 1.525 ;
        RECT -10.365 -0.165 -10.035 0.165 ;
        RECT -10.365 -1.525 -10.035 -1.195 ;
        RECT -10.365 -2.885 -10.035 -2.555 ;
        RECT -10.365 -4.245 -10.035 -3.915 ;
        RECT -10.365 -5.605 -10.035 -5.275 ;
        RECT -10.365 -8.325 -10.035 -7.995 ;
        RECT -10.365 -9.685 -10.035 -9.355 ;
        RECT -10.365 -11.16 -10.035 -10.83 ;
        RECT -10.365 -12.405 -10.035 -12.075 ;
        RECT -10.365 -15.125 -10.035 -14.795 ;
        RECT -10.365 -16.25 -10.035 -15.92 ;
        RECT -10.365 -21.925 -10.035 -21.595 ;
        RECT -10.365 -23.285 -10.035 -22.955 ;
        RECT -10.365 -24.645 -10.035 -24.315 ;
        RECT -10.365 -26.005 -10.035 -25.675 ;
        RECT -10.365 -27.365 -10.035 -27.035 ;
        RECT -10.365 -30.085 -10.035 -29.755 ;
        RECT -10.365 -31.445 -10.035 -31.115 ;
        RECT -10.365 -32.34 -10.035 -32.01 ;
        RECT -10.365 -34.165 -10.035 -33.835 ;
        RECT -10.365 -37.43 -10.035 -37.1 ;
        RECT -10.365 -38.245 -10.035 -37.915 ;
        RECT -10.365 -43.685 -10.035 -43.355 ;
        RECT -10.365 -45.045 -10.035 -44.715 ;
        RECT -10.365 -46.405 -10.035 -46.075 ;
        RECT -10.365 -47.765 -10.035 -47.435 ;
        RECT -10.365 -49.125 -10.035 -48.795 ;
        RECT -10.365 -50.485 -10.035 -50.155 ;
        RECT -10.365 -53.205 -10.035 -52.875 ;
        RECT -10.365 -54.565 -10.035 -54.235 ;
        RECT -10.365 -55.925 -10.035 -55.595 ;
        RECT -10.365 -57.285 -10.035 -56.955 ;
        RECT -10.365 -58.645 -10.035 -58.315 ;
        RECT -10.365 -61.67 -10.035 -61.34 ;
        RECT -10.365 -65.445 -10.035 -65.115 ;
        RECT -10.365 -66.805 -10.035 -66.475 ;
        RECT -10.365 -68.165 -10.035 -67.835 ;
        RECT -10.365 -69.525 -10.035 -69.195 ;
        RECT -10.365 -72.245 -10.035 -71.915 ;
        RECT -10.365 -73.605 -10.035 -73.275 ;
        RECT -10.365 -74.965 -10.035 -74.635 ;
        RECT -10.365 -76.325 -10.035 -75.995 ;
        RECT -10.365 -77.685 -10.035 -77.355 ;
        RECT -10.365 -79.045 -10.035 -78.715 ;
        RECT -10.365 -80.21 -10.035 -79.88 ;
        RECT -10.365 -81.765 -10.035 -81.435 ;
        RECT -10.365 -83.125 -10.035 -82.795 ;
        RECT -10.365 -84.485 -10.035 -84.155 ;
        RECT -10.365 -87.205 -10.035 -86.875 ;
        RECT -10.365 -88.565 -10.035 -88.235 ;
        RECT -10.365 -89.925 -10.035 -89.595 ;
        RECT -10.365 -91.285 -10.035 -90.955 ;
        RECT -10.365 -92.645 -10.035 -92.315 ;
        RECT -10.365 -94.005 -10.035 -93.675 ;
        RECT -10.365 -95.365 -10.035 -95.035 ;
        RECT -10.365 -98.085 -10.035 -97.755 ;
        RECT -10.365 -99.445 -10.035 -99.115 ;
        RECT -10.365 -100.805 -10.035 -100.475 ;
        RECT -10.365 -102.165 -10.035 -101.835 ;
        RECT -10.365 -103.525 -10.035 -103.195 ;
        RECT -10.365 -104.885 -10.035 -104.555 ;
        RECT -10.365 -105.85 -10.035 -105.52 ;
        RECT -10.365 -107.605 -10.035 -107.275 ;
        RECT -10.365 -108.965 -10.035 -108.635 ;
        RECT -10.365 -110.325 -10.035 -109.995 ;
        RECT -10.365 -111.685 -10.035 -111.355 ;
        RECT -10.365 -115.765 -10.035 -115.435 ;
        RECT -10.365 -117.125 -10.035 -116.795 ;
        RECT -10.365 -118.485 -10.035 -118.155 ;
        RECT -10.365 -119.845 -10.035 -119.515 ;
        RECT -10.365 -121.205 -10.035 -120.875 ;
        RECT -10.365 -122.565 -10.035 -122.235 ;
        RECT -10.365 -124.39 -10.035 -124.06 ;
        RECT -10.365 -125.285 -10.035 -124.955 ;
        RECT -10.365 -126.645 -10.035 -126.315 ;
        RECT -10.365 -128.005 -10.035 -127.675 ;
        RECT -10.365 -129.365 -10.035 -129.035 ;
        RECT -10.365 -133.445 -10.035 -133.115 ;
        RECT -10.365 -134.805 -10.035 -134.475 ;
        RECT -10.365 -136.165 -10.035 -135.835 ;
        RECT -10.365 -137.525 -10.035 -137.195 ;
        RECT -10.365 -138.885 -10.035 -138.555 ;
        RECT -10.365 -140.245 -10.035 -139.915 ;
        RECT -10.365 -144.325 -10.035 -143.995 ;
        RECT -10.365 -145.685 -10.035 -145.355 ;
        RECT -10.365 -147.045 -10.035 -146.715 ;
        RECT -10.365 -148.405 -10.035 -148.075 ;
        RECT -10.365 -151.125 -10.035 -150.795 ;
        RECT -10.365 -152.485 -10.035 -152.155 ;
        RECT -10.365 -153.845 -10.035 -153.515 ;
        RECT -10.365 -155.205 -10.035 -154.875 ;
        RECT -10.365 -156.565 -10.035 -156.235 ;
        RECT -10.365 -157.925 -10.035 -157.595 ;
        RECT -10.365 -159.285 -10.035 -158.955 ;
        RECT -10.365 -160.645 -10.035 -160.315 ;
        RECT -10.365 -162.005 -10.035 -161.675 ;
        RECT -10.365 -163.365 -10.035 -163.035 ;
        RECT -10.365 -164.725 -10.035 -164.395 ;
        RECT -10.365 -166.085 -10.035 -165.755 ;
        RECT -10.365 -167.445 -10.035 -167.115 ;
        RECT -10.365 -168.805 -10.035 -168.475 ;
        RECT -10.365 -170.165 -10.035 -169.835 ;
        RECT -10.365 -171.525 -10.035 -171.195 ;
        RECT -10.365 -172.885 -10.035 -172.555 ;
        RECT -10.365 -174.245 -10.035 -173.915 ;
        RECT -10.365 -175.605 -10.035 -175.275 ;
        RECT -10.365 -176.965 -10.035 -176.635 ;
        RECT -10.365 -178.325 -10.035 -177.995 ;
        RECT -10.365 -179.685 -10.035 -179.355 ;
        RECT -10.365 -183.765 -10.035 -183.435 ;
        RECT -10.365 -185.125 -10.035 -184.795 ;
        RECT -10.365 -186.485 -10.035 -186.155 ;
        RECT -10.365 -187.845 -10.035 -187.515 ;
        RECT -10.365 -189.205 -10.035 -188.875 ;
        RECT -10.365 -190.565 -10.035 -190.235 ;
        RECT -10.365 -191.925 -10.035 -191.595 ;
        RECT -10.365 -193.285 -10.035 -192.955 ;
        RECT -10.365 -194.645 -10.035 -194.315 ;
        RECT -10.365 -196.005 -10.035 -195.675 ;
        RECT -10.365 -197.365 -10.035 -197.035 ;
        RECT -10.365 -198.725 -10.035 -198.395 ;
        RECT -10.365 -200.085 -10.035 -199.755 ;
        RECT -10.365 -201.445 -10.035 -201.115 ;
        RECT -10.365 -202.805 -10.035 -202.475 ;
        RECT -10.365 -204.165 -10.035 -203.835 ;
        RECT -10.36 -204.84 -10.04 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -10.365 -212.325 -10.035 -211.995 ;
        RECT -10.365 -215.045 -10.035 -214.715 ;
        RECT -10.365 -216.405 -10.035 -216.075 ;
        RECT -10.365 -217.765 -10.035 -217.435 ;
        RECT -10.365 -219.125 -10.035 -218.795 ;
        RECT -10.365 -221.37 -10.035 -220.24 ;
        RECT -10.36 -221.485 -10.04 -210.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.005 129.8 -8.675 130.93 ;
        RECT -9.005 127.675 -8.675 128.005 ;
        RECT -9.005 126.315 -8.675 126.645 ;
        RECT -9.005 124.955 -8.675 125.285 ;
        RECT -9.005 123.595 -8.675 123.925 ;
        RECT -9.005 122.235 -8.675 122.565 ;
        RECT -9.005 120.875 -8.675 121.205 ;
        RECT -9.005 119.515 -8.675 119.845 ;
        RECT -9.005 118.155 -8.675 118.485 ;
        RECT -9.005 114.075 -8.675 114.405 ;
        RECT -9.005 104.555 -8.675 104.885 ;
        RECT -9.005 103.195 -8.675 103.525 ;
        RECT -9.005 96.395 -8.675 96.725 ;
        RECT -9.005 93.675 -8.675 94.005 ;
        RECT -9.005 89.595 -8.675 89.925 ;
        RECT -9.005 85.515 -8.675 85.845 ;
        RECT -9.005 82.795 -8.675 83.125 ;
        RECT -9.005 75.995 -8.675 76.325 ;
        RECT -9.005 74.635 -8.675 74.965 ;
        RECT -9.005 65.115 -8.675 65.445 ;
        RECT -9.005 61.035 -8.675 61.365 ;
        RECT -9.005 56.955 -8.675 57.285 ;
        RECT -9.005 54.235 -8.675 54.565 ;
        RECT -9.005 47.435 -8.675 47.765 ;
        RECT -9.005 46.075 -8.675 46.405 ;
        RECT -9.005 43.355 -8.675 43.685 ;
        RECT -9.005 36.555 -8.675 36.885 ;
        RECT -9.005 33.835 -8.675 34.165 ;
        RECT -9.005 32.475 -8.675 32.805 ;
        RECT -9.005 28.395 -8.675 28.725 ;
        RECT -9.005 25.675 -8.675 26.005 ;
        RECT -9.005 18.875 -8.675 19.205 ;
        RECT -9.005 17.515 -8.675 17.845 ;
        RECT -9.005 14.795 -8.675 15.125 ;
        RECT -9.005 7.995 -8.675 8.325 ;
        RECT -9.005 5.275 -8.675 5.605 ;
        RECT -9.005 3.915 -8.675 4.245 ;
        RECT -9.005 2.555 -8.675 2.885 ;
        RECT -9.005 1.195 -8.675 1.525 ;
        RECT -9.005 -0.165 -8.675 0.165 ;
        RECT -9.005 -1.525 -8.675 -1.195 ;
        RECT -9.005 -2.885 -8.675 -2.555 ;
        RECT -9.005 -4.245 -8.675 -3.915 ;
        RECT -9.005 -5.605 -8.675 -5.275 ;
        RECT -9.005 -6.965 -8.675 -6.635 ;
        RECT -9.005 -8.325 -8.675 -7.995 ;
        RECT -9.005 -9.685 -8.675 -9.355 ;
        RECT -9 -9.685 -8.68 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.005 -142.965 -8.675 -142.635 ;
        RECT -9.005 -144.325 -8.675 -143.995 ;
        RECT -9.005 -145.685 -8.675 -145.355 ;
        RECT -9.005 -147.045 -8.675 -146.715 ;
        RECT -9.005 -148.405 -8.675 -148.075 ;
        RECT -9.005 -149.765 -8.675 -149.435 ;
        RECT -9.005 -151.125 -8.675 -150.795 ;
        RECT -9.005 -152.485 -8.675 -152.155 ;
        RECT -9.005 -153.845 -8.675 -153.515 ;
        RECT -9.005 -155.205 -8.675 -154.875 ;
        RECT -9.005 -156.565 -8.675 -156.235 ;
        RECT -9.005 -157.925 -8.675 -157.595 ;
        RECT -9.005 -159.285 -8.675 -158.955 ;
        RECT -9.005 -160.645 -8.675 -160.315 ;
        RECT -9.005 -162.005 -8.675 -161.675 ;
        RECT -9.005 -163.365 -8.675 -163.035 ;
        RECT -9.005 -164.725 -8.675 -164.395 ;
        RECT -9.005 -166.085 -8.675 -165.755 ;
        RECT -9.005 -167.445 -8.675 -167.115 ;
        RECT -9.005 -168.805 -8.675 -168.475 ;
        RECT -9.005 -170.165 -8.675 -169.835 ;
        RECT -9.005 -171.525 -8.675 -171.195 ;
        RECT -9.005 -172.885 -8.675 -172.555 ;
        RECT -9.005 -174.245 -8.675 -173.915 ;
        RECT -9.005 -175.605 -8.675 -175.275 ;
        RECT -9.005 -176.965 -8.675 -176.635 ;
        RECT -9.005 -178.325 -8.675 -177.995 ;
        RECT -9.005 -179.685 -8.675 -179.355 ;
        RECT -9.005 -181.045 -8.675 -180.715 ;
        RECT -9.005 -182.405 -8.675 -182.075 ;
        RECT -9.005 -183.765 -8.675 -183.435 ;
        RECT -9.005 -185.125 -8.675 -184.795 ;
        RECT -9.005 -186.485 -8.675 -186.155 ;
        RECT -9.005 -187.845 -8.675 -187.515 ;
        RECT -9.005 -189.205 -8.675 -188.875 ;
        RECT -9.005 -190.565 -8.675 -190.235 ;
        RECT -9.005 -191.925 -8.675 -191.595 ;
        RECT -9.005 -193.285 -8.675 -192.955 ;
        RECT -9.005 -194.645 -8.675 -194.315 ;
        RECT -9.005 -196.005 -8.675 -195.675 ;
        RECT -9.005 -197.365 -8.675 -197.035 ;
        RECT -9.005 -198.725 -8.675 -198.395 ;
        RECT -9.005 -200.085 -8.675 -199.755 ;
        RECT -9.005 -201.445 -8.675 -201.115 ;
        RECT -9.005 -202.805 -8.675 -202.475 ;
        RECT -9.005 -204.165 -8.675 -203.835 ;
        RECT -9.005 -205.525 -8.675 -205.195 ;
        RECT -9.005 -206.885 -8.675 -206.555 ;
        RECT -9.005 -208.245 -8.675 -207.915 ;
        RECT -9.005 -209.605 -8.675 -209.275 ;
        RECT -9.005 -210.965 -8.675 -210.635 ;
        RECT -9.005 -212.325 -8.675 -211.995 ;
        RECT -9.005 -213.685 -8.675 -213.355 ;
        RECT -9.005 -215.045 -8.675 -214.715 ;
        RECT -9.005 -216.405 -8.675 -216.075 ;
        RECT -9.005 -217.765 -8.675 -217.435 ;
        RECT -9.005 -219.125 -8.675 -218.795 ;
        RECT -9.005 -221.37 -8.675 -220.24 ;
        RECT -9 -221.485 -8.68 -141.96 ;
    END
    PORT
      LAYER met3 ;
        RECT -7.645 74.635 -7.315 74.965 ;
        RECT -7.645 65.115 -7.315 65.445 ;
        RECT -7.645 61.035 -7.315 61.365 ;
        RECT -7.645 56.955 -7.315 57.285 ;
        RECT -7.645 54.235 -7.315 54.565 ;
        RECT -7.645 47.435 -7.315 47.765 ;
        RECT -7.645 46.075 -7.315 46.405 ;
        RECT -7.645 43.355 -7.315 43.685 ;
        RECT -7.645 36.555 -7.315 36.885 ;
        RECT -7.645 33.835 -7.315 34.165 ;
        RECT -7.645 32.475 -7.315 32.805 ;
        RECT -7.645 28.395 -7.315 28.725 ;
        RECT -7.645 25.675 -7.315 26.005 ;
        RECT -7.645 18.875 -7.315 19.205 ;
        RECT -7.645 17.515 -7.315 17.845 ;
        RECT -7.645 14.795 -7.315 15.125 ;
        RECT -7.645 7.995 -7.315 8.325 ;
        RECT -7.645 5.275 -7.315 5.605 ;
        RECT -7.645 3.915 -7.315 4.245 ;
        RECT -7.645 2.555 -7.315 2.885 ;
        RECT -7.645 1.195 -7.315 1.525 ;
        RECT -7.645 -0.165 -7.315 0.165 ;
        RECT -7.645 -1.525 -7.315 -1.195 ;
        RECT -7.645 -2.885 -7.315 -2.555 ;
        RECT -7.645 -4.245 -7.315 -3.915 ;
        RECT -7.645 -5.605 -7.315 -5.275 ;
        RECT -7.645 -6.965 -7.315 -6.635 ;
        RECT -7.645 -8.325 -7.315 -7.995 ;
        RECT -7.645 -9.685 -7.315 -9.355 ;
        RECT -7.645 -12.405 -7.315 -12.075 ;
        RECT -7.645 -13.765 -7.315 -13.435 ;
        RECT -7.645 -15.125 -7.315 -14.795 ;
        RECT -7.645 -16.485 -7.315 -16.155 ;
        RECT -7.645 -17.845 -7.315 -17.515 ;
        RECT -7.645 -19.205 -7.315 -18.875 ;
        RECT -7.645 -20.565 -7.315 -20.235 ;
        RECT -7.645 -21.925 -7.315 -21.595 ;
        RECT -7.645 -23.285 -7.315 -22.955 ;
        RECT -7.645 -24.645 -7.315 -24.315 ;
        RECT -7.645 -26.005 -7.315 -25.675 ;
        RECT -7.645 -27.365 -7.315 -27.035 ;
        RECT -7.645 -28.725 -7.315 -28.395 ;
        RECT -7.645 -30.085 -7.315 -29.755 ;
        RECT -7.645 -31.445 -7.315 -31.115 ;
        RECT -7.645 -32.805 -7.315 -32.475 ;
        RECT -7.645 -34.165 -7.315 -33.835 ;
        RECT -7.645 -35.525 -7.315 -35.195 ;
        RECT -7.645 -36.885 -7.315 -36.555 ;
        RECT -7.645 -38.245 -7.315 -37.915 ;
        RECT -7.645 -39.605 -7.315 -39.275 ;
        RECT -7.645 -40.965 -7.315 -40.635 ;
        RECT -7.645 -42.325 -7.315 -41.995 ;
        RECT -7.645 -43.685 -7.315 -43.355 ;
        RECT -7.645 -45.045 -7.315 -44.715 ;
        RECT -7.645 -46.405 -7.315 -46.075 ;
        RECT -7.645 -47.765 -7.315 -47.435 ;
        RECT -7.645 -49.125 -7.315 -48.795 ;
        RECT -7.645 -50.485 -7.315 -50.155 ;
        RECT -7.645 -51.845 -7.315 -51.515 ;
        RECT -7.645 -53.205 -7.315 -52.875 ;
        RECT -7.645 -54.565 -7.315 -54.235 ;
        RECT -7.645 -55.925 -7.315 -55.595 ;
        RECT -7.645 -57.285 -7.315 -56.955 ;
        RECT -7.645 -58.645 -7.315 -58.315 ;
        RECT -7.645 -61.365 -7.315 -61.035 ;
        RECT -7.645 -65.445 -7.315 -65.115 ;
        RECT -7.645 -66.805 -7.315 -66.475 ;
        RECT -7.645 -68.165 -7.315 -67.835 ;
        RECT -7.645 -69.525 -7.315 -69.195 ;
        RECT -7.645 -70.885 -7.315 -70.555 ;
        RECT -7.645 -72.245 -7.315 -71.915 ;
        RECT -7.645 -73.605 -7.315 -73.275 ;
        RECT -7.645 -74.965 -7.315 -74.635 ;
        RECT -7.645 -76.325 -7.315 -75.995 ;
        RECT -7.645 -77.685 -7.315 -77.355 ;
        RECT -7.645 -79.045 -7.315 -78.715 ;
        RECT -7.645 -80.405 -7.315 -80.075 ;
        RECT -7.645 -81.765 -7.315 -81.435 ;
        RECT -7.645 -83.125 -7.315 -82.795 ;
        RECT -7.645 -84.485 -7.315 -84.155 ;
        RECT -7.645 -85.845 -7.315 -85.515 ;
        RECT -7.645 -87.205 -7.315 -86.875 ;
        RECT -7.645 -88.565 -7.315 -88.235 ;
        RECT -7.645 -89.925 -7.315 -89.595 ;
        RECT -7.645 -91.285 -7.315 -90.955 ;
        RECT -7.645 -92.645 -7.315 -92.315 ;
        RECT -7.645 -94.005 -7.315 -93.675 ;
        RECT -7.645 -95.365 -7.315 -95.035 ;
        RECT -7.645 -96.725 -7.315 -96.395 ;
        RECT -7.645 -98.085 -7.315 -97.755 ;
        RECT -7.645 -99.445 -7.315 -99.115 ;
        RECT -7.645 -100.805 -7.315 -100.475 ;
        RECT -7.645 -102.165 -7.315 -101.835 ;
        RECT -7.645 -103.525 -7.315 -103.195 ;
        RECT -7.645 -104.885 -7.315 -104.555 ;
        RECT -7.645 -106.245 -7.315 -105.915 ;
        RECT -7.645 -107.605 -7.315 -107.275 ;
        RECT -7.645 -108.965 -7.315 -108.635 ;
        RECT -7.645 -110.325 -7.315 -109.995 ;
        RECT -7.645 -111.685 -7.315 -111.355 ;
        RECT -7.645 -114.405 -7.315 -114.075 ;
        RECT -7.645 -115.765 -7.315 -115.435 ;
        RECT -7.645 -117.125 -7.315 -116.795 ;
        RECT -7.645 -118.485 -7.315 -118.155 ;
        RECT -7.645 -119.845 -7.315 -119.515 ;
        RECT -7.645 -121.205 -7.315 -120.875 ;
        RECT -7.645 -122.565 -7.315 -122.235 ;
        RECT -7.645 -123.925 -7.315 -123.595 ;
        RECT -7.645 -125.285 -7.315 -124.955 ;
        RECT -7.645 -126.645 -7.315 -126.315 ;
        RECT -7.645 -128.005 -7.315 -127.675 ;
        RECT -7.645 -129.365 -7.315 -129.035 ;
        RECT -7.645 -130.725 -7.315 -130.395 ;
        RECT -7.645 -132.085 -7.315 -131.755 ;
        RECT -7.645 -133.445 -7.315 -133.115 ;
        RECT -7.645 -134.805 -7.315 -134.475 ;
        RECT -7.645 -136.165 -7.315 -135.835 ;
        RECT -7.645 -137.525 -7.315 -137.195 ;
        RECT -7.645 -138.885 -7.315 -138.555 ;
        RECT -7.645 -140.245 -7.315 -139.915 ;
        RECT -7.645 -141.605 -7.315 -141.275 ;
        RECT -7.645 -142.965 -7.315 -142.635 ;
        RECT -7.645 -144.325 -7.315 -143.995 ;
        RECT -7.645 -145.685 -7.315 -145.355 ;
        RECT -7.645 -147.045 -7.315 -146.715 ;
        RECT -7.645 -148.405 -7.315 -148.075 ;
        RECT -7.645 -149.765 -7.315 -149.435 ;
        RECT -7.645 -151.125 -7.315 -150.795 ;
        RECT -7.645 -152.485 -7.315 -152.155 ;
        RECT -7.645 -153.845 -7.315 -153.515 ;
        RECT -7.645 -155.205 -7.315 -154.875 ;
        RECT -7.645 -156.565 -7.315 -156.235 ;
        RECT -7.645 -157.925 -7.315 -157.595 ;
        RECT -7.645 -159.285 -7.315 -158.955 ;
        RECT -7.645 -160.645 -7.315 -160.315 ;
        RECT -7.645 -162.005 -7.315 -161.675 ;
        RECT -7.645 -163.365 -7.315 -163.035 ;
        RECT -7.645 -164.725 -7.315 -164.395 ;
        RECT -7.645 -166.085 -7.315 -165.755 ;
        RECT -7.645 -167.445 -7.315 -167.115 ;
        RECT -7.645 -168.805 -7.315 -168.475 ;
        RECT -7.645 -170.165 -7.315 -169.835 ;
        RECT -7.645 -171.525 -7.315 -171.195 ;
        RECT -7.645 -172.885 -7.315 -172.555 ;
        RECT -7.645 -174.245 -7.315 -173.915 ;
        RECT -7.645 -175.605 -7.315 -175.275 ;
        RECT -7.645 -176.965 -7.315 -176.635 ;
        RECT -7.645 -178.325 -7.315 -177.995 ;
        RECT -7.645 -179.685 -7.315 -179.355 ;
        RECT -7.645 -181.045 -7.315 -180.715 ;
        RECT -7.645 -182.405 -7.315 -182.075 ;
        RECT -7.645 -183.765 -7.315 -183.435 ;
        RECT -7.645 -185.125 -7.315 -184.795 ;
        RECT -7.645 -186.485 -7.315 -186.155 ;
        RECT -7.645 -187.845 -7.315 -187.515 ;
        RECT -7.645 -189.205 -7.315 -188.875 ;
        RECT -7.645 -190.565 -7.315 -190.235 ;
        RECT -7.645 -191.925 -7.315 -191.595 ;
        RECT -7.645 -193.285 -7.315 -192.955 ;
        RECT -7.645 -194.645 -7.315 -194.315 ;
        RECT -7.645 -196.005 -7.315 -195.675 ;
        RECT -7.645 -197.365 -7.315 -197.035 ;
        RECT -7.645 -198.725 -7.315 -198.395 ;
        RECT -7.645 -200.085 -7.315 -199.755 ;
        RECT -7.645 -201.445 -7.315 -201.115 ;
        RECT -7.645 -202.805 -7.315 -202.475 ;
        RECT -7.645 -204.165 -7.315 -203.835 ;
        RECT -7.645 -205.525 -7.315 -205.195 ;
        RECT -7.645 -206.885 -7.315 -206.555 ;
        RECT -7.645 -208.245 -7.315 -207.915 ;
        RECT -7.645 -209.605 -7.315 -209.275 ;
        RECT -7.645 -210.965 -7.315 -210.635 ;
        RECT -7.645 -212.325 -7.315 -211.995 ;
        RECT -7.645 -213.685 -7.315 -213.355 ;
        RECT -7.645 -215.045 -7.315 -214.715 ;
        RECT -7.645 -216.405 -7.315 -216.075 ;
        RECT -7.645 -217.765 -7.315 -217.435 ;
        RECT -7.645 -219.125 -7.315 -218.795 ;
        RECT -7.645 -221.37 -7.315 -220.24 ;
        RECT -7.64 -221.485 -7.32 131.045 ;
        RECT -7.645 129.8 -7.315 130.93 ;
        RECT -7.645 127.675 -7.315 128.005 ;
        RECT -7.645 126.315 -7.315 126.645 ;
        RECT -7.645 124.955 -7.315 125.285 ;
        RECT -7.645 123.595 -7.315 123.925 ;
        RECT -7.645 122.235 -7.315 122.565 ;
        RECT -7.645 120.875 -7.315 121.205 ;
        RECT -7.645 119.515 -7.315 119.845 ;
        RECT -7.645 118.155 -7.315 118.485 ;
        RECT -7.645 114.075 -7.315 114.405 ;
        RECT -7.645 104.555 -7.315 104.885 ;
        RECT -7.645 103.195 -7.315 103.525 ;
        RECT -7.645 96.395 -7.315 96.725 ;
        RECT -7.645 93.675 -7.315 94.005 ;
        RECT -7.645 89.595 -7.315 89.925 ;
        RECT -7.645 85.515 -7.315 85.845 ;
        RECT -7.645 82.795 -7.315 83.125 ;
        RECT -7.645 75.995 -7.315 76.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.245 129.8 -20.915 130.93 ;
        RECT -21.245 127.675 -20.915 128.005 ;
        RECT -21.245 126.315 -20.915 126.645 ;
        RECT -21.245 124.955 -20.915 125.285 ;
        RECT -21.245 123.595 -20.915 123.925 ;
        RECT -21.245 122.235 -20.915 122.565 ;
        RECT -21.245 120.875 -20.915 121.205 ;
        RECT -21.245 119.515 -20.915 119.845 ;
        RECT -21.245 118.155 -20.915 118.485 ;
        RECT -21.245 116.795 -20.915 117.125 ;
        RECT -21.245 115.435 -20.915 115.765 ;
        RECT -21.245 114.075 -20.915 114.405 ;
        RECT -21.245 112.715 -20.915 113.045 ;
        RECT -21.245 111.355 -20.915 111.685 ;
        RECT -21.245 109.995 -20.915 110.325 ;
        RECT -21.245 108.635 -20.915 108.965 ;
        RECT -21.245 107.275 -20.915 107.605 ;
        RECT -21.245 105.915 -20.915 106.245 ;
        RECT -21.245 104.555 -20.915 104.885 ;
        RECT -21.245 103.195 -20.915 103.525 ;
        RECT -21.245 101.835 -20.915 102.165 ;
        RECT -21.245 100.475 -20.915 100.805 ;
        RECT -21.245 99.115 -20.915 99.445 ;
        RECT -21.245 97.755 -20.915 98.085 ;
        RECT -21.245 96.395 -20.915 96.725 ;
        RECT -21.245 95.035 -20.915 95.365 ;
        RECT -21.245 93.675 -20.915 94.005 ;
        RECT -21.245 92.315 -20.915 92.645 ;
        RECT -21.245 90.955 -20.915 91.285 ;
        RECT -21.245 89.595 -20.915 89.925 ;
        RECT -21.245 88.235 -20.915 88.565 ;
        RECT -21.245 86.875 -20.915 87.205 ;
        RECT -21.245 85.515 -20.915 85.845 ;
        RECT -21.245 84.155 -20.915 84.485 ;
        RECT -21.245 82.795 -20.915 83.125 ;
        RECT -21.245 81.435 -20.915 81.765 ;
        RECT -21.245 80.075 -20.915 80.405 ;
        RECT -21.245 78.715 -20.915 79.045 ;
        RECT -21.245 77.355 -20.915 77.685 ;
        RECT -21.245 75.995 -20.915 76.325 ;
        RECT -21.245 74.635 -20.915 74.965 ;
        RECT -21.245 73.275 -20.915 73.605 ;
        RECT -21.245 71.915 -20.915 72.245 ;
        RECT -21.245 70.555 -20.915 70.885 ;
        RECT -21.245 69.195 -20.915 69.525 ;
        RECT -21.245 67.835 -20.915 68.165 ;
        RECT -21.245 66.475 -20.915 66.805 ;
        RECT -21.245 65.115 -20.915 65.445 ;
        RECT -21.245 63.755 -20.915 64.085 ;
        RECT -21.245 62.395 -20.915 62.725 ;
        RECT -21.245 61.035 -20.915 61.365 ;
        RECT -21.245 59.675 -20.915 60.005 ;
        RECT -21.245 58.315 -20.915 58.645 ;
        RECT -21.245 56.955 -20.915 57.285 ;
        RECT -21.245 55.595 -20.915 55.925 ;
        RECT -21.245 54.235 -20.915 54.565 ;
        RECT -21.245 52.875 -20.915 53.205 ;
        RECT -21.245 51.515 -20.915 51.845 ;
        RECT -21.245 50.155 -20.915 50.485 ;
        RECT -21.245 48.795 -20.915 49.125 ;
        RECT -21.245 47.435 -20.915 47.765 ;
        RECT -21.245 46.075 -20.915 46.405 ;
        RECT -21.245 44.715 -20.915 45.045 ;
        RECT -21.245 43.355 -20.915 43.685 ;
        RECT -21.245 41.995 -20.915 42.325 ;
        RECT -21.245 40.635 -20.915 40.965 ;
        RECT -21.245 39.275 -20.915 39.605 ;
        RECT -21.245 37.915 -20.915 38.245 ;
        RECT -21.245 36.555 -20.915 36.885 ;
        RECT -21.245 35.195 -20.915 35.525 ;
        RECT -21.245 33.835 -20.915 34.165 ;
        RECT -21.245 32.475 -20.915 32.805 ;
        RECT -21.245 31.115 -20.915 31.445 ;
        RECT -21.245 29.755 -20.915 30.085 ;
        RECT -21.245 28.395 -20.915 28.725 ;
        RECT -21.245 27.035 -20.915 27.365 ;
        RECT -21.245 25.675 -20.915 26.005 ;
        RECT -21.245 24.315 -20.915 24.645 ;
        RECT -21.245 22.955 -20.915 23.285 ;
        RECT -21.245 21.595 -20.915 21.925 ;
        RECT -21.245 20.235 -20.915 20.565 ;
        RECT -21.245 18.875 -20.915 19.205 ;
        RECT -21.245 17.515 -20.915 17.845 ;
        RECT -21.245 16.155 -20.915 16.485 ;
        RECT -21.245 14.795 -20.915 15.125 ;
        RECT -21.245 13.435 -20.915 13.765 ;
        RECT -21.245 12.075 -20.915 12.405 ;
        RECT -21.245 10.715 -20.915 11.045 ;
        RECT -21.245 9.355 -20.915 9.685 ;
        RECT -21.245 7.995 -20.915 8.325 ;
        RECT -21.245 6.635 -20.915 6.965 ;
        RECT -21.245 5.275 -20.915 5.605 ;
        RECT -21.245 3.915 -20.915 4.245 ;
        RECT -21.245 2.555 -20.915 2.885 ;
        RECT -21.245 1.195 -20.915 1.525 ;
        RECT -21.245 -0.165 -20.915 0.165 ;
        RECT -21.245 -1.525 -20.915 -1.195 ;
        RECT -21.245 -2.885 -20.915 -2.555 ;
        RECT -21.245 -8.325 -20.915 -7.995 ;
        RECT -21.245 -9.685 -20.915 -9.355 ;
        RECT -21.245 -11.16 -20.915 -10.83 ;
        RECT -21.245 -12.405 -20.915 -12.075 ;
        RECT -21.245 -15.125 -20.915 -14.795 ;
        RECT -21.245 -16.25 -20.915 -15.92 ;
        RECT -21.24 -19.2 -20.92 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.245 -32.34 -20.915 -32.01 ;
        RECT -21.245 -37.43 -20.915 -37.1 ;
        RECT -21.24 -40.28 -20.92 -31.8 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.245 -108.965 -20.915 -108.635 ;
        RECT -21.245 -110.325 -20.915 -109.995 ;
        RECT -21.245 -111.685 -20.915 -111.355 ;
        RECT -21.245 -113.045 -20.915 -112.715 ;
        RECT -21.245 -114.405 -20.915 -114.075 ;
        RECT -21.245 -115.765 -20.915 -115.435 ;
        RECT -21.245 -117.125 -20.915 -116.795 ;
        RECT -21.245 -118.485 -20.915 -118.155 ;
        RECT -21.245 -119.845 -20.915 -119.515 ;
        RECT -21.245 -121.205 -20.915 -120.875 ;
        RECT -21.245 -122.565 -20.915 -122.235 ;
        RECT -21.245 -123.925 -20.915 -123.595 ;
        RECT -21.245 -125.285 -20.915 -124.955 ;
        RECT -21.245 -126.645 -20.915 -126.315 ;
        RECT -21.245 -128.005 -20.915 -127.675 ;
        RECT -21.245 -129.365 -20.915 -129.035 ;
        RECT -21.245 -130.725 -20.915 -130.395 ;
        RECT -21.245 -132.085 -20.915 -131.755 ;
        RECT -21.245 -133.445 -20.915 -133.115 ;
        RECT -21.245 -134.805 -20.915 -134.475 ;
        RECT -21.245 -136.165 -20.915 -135.835 ;
        RECT -21.245 -137.525 -20.915 -137.195 ;
        RECT -21.245 -142.965 -20.915 -142.635 ;
        RECT -21.245 -144.325 -20.915 -143.995 ;
        RECT -21.245 -145.685 -20.915 -145.355 ;
        RECT -21.245 -147.045 -20.915 -146.715 ;
        RECT -21.245 -148.405 -20.915 -148.075 ;
        RECT -21.245 -149.765 -20.915 -149.435 ;
        RECT -21.245 -151.125 -20.915 -150.795 ;
        RECT -21.245 -152.485 -20.915 -152.155 ;
        RECT -21.245 -155.205 -20.915 -154.875 ;
        RECT -21.245 -156.565 -20.915 -156.235 ;
        RECT -21.245 -157.925 -20.915 -157.595 ;
        RECT -21.245 -159.285 -20.915 -158.955 ;
        RECT -21.245 -160.645 -20.915 -160.315 ;
        RECT -21.245 -162.005 -20.915 -161.675 ;
        RECT -21.245 -163.365 -20.915 -163.035 ;
        RECT -21.245 -172.885 -20.915 -172.555 ;
        RECT -21.245 -175.605 -20.915 -175.275 ;
        RECT -21.245 -176.965 -20.915 -176.635 ;
        RECT -21.245 -179.685 -20.915 -179.355 ;
        RECT -21.245 -181.045 -20.915 -180.715 ;
        RECT -21.245 -183.765 -20.915 -183.435 ;
        RECT -21.245 -185.125 -20.915 -184.795 ;
        RECT -21.245 -189.205 -20.915 -188.875 ;
        RECT -21.245 -190.565 -20.915 -190.235 ;
        RECT -21.245 -194.645 -20.915 -194.315 ;
        RECT -21.245 -196.005 -20.915 -195.675 ;
        RECT -21.245 -197.365 -20.915 -197.035 ;
        RECT -21.245 -198.725 -20.915 -198.395 ;
        RECT -21.245 -200.085 -20.915 -199.755 ;
        RECT -21.245 -201.445 -20.915 -201.115 ;
        RECT -21.245 -202.805 -20.915 -202.475 ;
        RECT -21.245 -204.165 -20.915 -203.835 ;
        RECT -21.245 -205.525 -20.915 -205.195 ;
        RECT -21.245 -208.245 -20.915 -207.915 ;
        RECT -21.24 -209.6 -20.92 -106.6 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.885 129.8 -19.555 130.93 ;
        RECT -19.885 127.675 -19.555 128.005 ;
        RECT -19.885 126.315 -19.555 126.645 ;
        RECT -19.885 124.955 -19.555 125.285 ;
        RECT -19.885 123.595 -19.555 123.925 ;
        RECT -19.885 122.235 -19.555 122.565 ;
        RECT -19.885 120.875 -19.555 121.205 ;
        RECT -19.885 119.515 -19.555 119.845 ;
        RECT -19.885 118.155 -19.555 118.485 ;
        RECT -19.885 116.795 -19.555 117.125 ;
        RECT -19.885 115.435 -19.555 115.765 ;
        RECT -19.885 114.075 -19.555 114.405 ;
        RECT -19.885 112.715 -19.555 113.045 ;
        RECT -19.885 111.355 -19.555 111.685 ;
        RECT -19.885 109.995 -19.555 110.325 ;
        RECT -19.885 108.635 -19.555 108.965 ;
        RECT -19.885 107.275 -19.555 107.605 ;
        RECT -19.885 105.915 -19.555 106.245 ;
        RECT -19.885 104.555 -19.555 104.885 ;
        RECT -19.885 103.195 -19.555 103.525 ;
        RECT -19.885 101.835 -19.555 102.165 ;
        RECT -19.885 100.475 -19.555 100.805 ;
        RECT -19.885 99.115 -19.555 99.445 ;
        RECT -19.885 97.755 -19.555 98.085 ;
        RECT -19.885 96.395 -19.555 96.725 ;
        RECT -19.885 95.035 -19.555 95.365 ;
        RECT -19.885 93.675 -19.555 94.005 ;
        RECT -19.885 92.315 -19.555 92.645 ;
        RECT -19.885 90.955 -19.555 91.285 ;
        RECT -19.885 89.595 -19.555 89.925 ;
        RECT -19.885 88.235 -19.555 88.565 ;
        RECT -19.885 86.875 -19.555 87.205 ;
        RECT -19.885 85.515 -19.555 85.845 ;
        RECT -19.885 84.155 -19.555 84.485 ;
        RECT -19.885 82.795 -19.555 83.125 ;
        RECT -19.885 81.435 -19.555 81.765 ;
        RECT -19.885 80.075 -19.555 80.405 ;
        RECT -19.885 78.715 -19.555 79.045 ;
        RECT -19.885 77.355 -19.555 77.685 ;
        RECT -19.885 75.995 -19.555 76.325 ;
        RECT -19.885 74.635 -19.555 74.965 ;
        RECT -19.885 73.275 -19.555 73.605 ;
        RECT -19.885 71.915 -19.555 72.245 ;
        RECT -19.885 70.555 -19.555 70.885 ;
        RECT -19.885 69.195 -19.555 69.525 ;
        RECT -19.885 67.835 -19.555 68.165 ;
        RECT -19.885 66.475 -19.555 66.805 ;
        RECT -19.885 65.115 -19.555 65.445 ;
        RECT -19.885 63.755 -19.555 64.085 ;
        RECT -19.885 62.395 -19.555 62.725 ;
        RECT -19.885 61.035 -19.555 61.365 ;
        RECT -19.885 59.675 -19.555 60.005 ;
        RECT -19.885 58.315 -19.555 58.645 ;
        RECT -19.885 56.955 -19.555 57.285 ;
        RECT -19.885 55.595 -19.555 55.925 ;
        RECT -19.885 54.235 -19.555 54.565 ;
        RECT -19.885 52.875 -19.555 53.205 ;
        RECT -19.885 51.515 -19.555 51.845 ;
        RECT -19.885 50.155 -19.555 50.485 ;
        RECT -19.885 48.795 -19.555 49.125 ;
        RECT -19.885 47.435 -19.555 47.765 ;
        RECT -19.885 46.075 -19.555 46.405 ;
        RECT -19.885 44.715 -19.555 45.045 ;
        RECT -19.885 43.355 -19.555 43.685 ;
        RECT -19.885 41.995 -19.555 42.325 ;
        RECT -19.885 40.635 -19.555 40.965 ;
        RECT -19.885 39.275 -19.555 39.605 ;
        RECT -19.885 37.915 -19.555 38.245 ;
        RECT -19.885 36.555 -19.555 36.885 ;
        RECT -19.885 35.195 -19.555 35.525 ;
        RECT -19.885 33.835 -19.555 34.165 ;
        RECT -19.885 32.475 -19.555 32.805 ;
        RECT -19.885 31.115 -19.555 31.445 ;
        RECT -19.885 29.755 -19.555 30.085 ;
        RECT -19.885 28.395 -19.555 28.725 ;
        RECT -19.885 27.035 -19.555 27.365 ;
        RECT -19.885 25.675 -19.555 26.005 ;
        RECT -19.885 24.315 -19.555 24.645 ;
        RECT -19.885 22.955 -19.555 23.285 ;
        RECT -19.885 21.595 -19.555 21.925 ;
        RECT -19.885 20.235 -19.555 20.565 ;
        RECT -19.885 18.875 -19.555 19.205 ;
        RECT -19.885 17.515 -19.555 17.845 ;
        RECT -19.885 16.155 -19.555 16.485 ;
        RECT -19.885 14.795 -19.555 15.125 ;
        RECT -19.885 13.435 -19.555 13.765 ;
        RECT -19.885 12.075 -19.555 12.405 ;
        RECT -19.885 10.715 -19.555 11.045 ;
        RECT -19.885 9.355 -19.555 9.685 ;
        RECT -19.885 7.995 -19.555 8.325 ;
        RECT -19.885 6.635 -19.555 6.965 ;
        RECT -19.885 5.275 -19.555 5.605 ;
        RECT -19.885 3.915 -19.555 4.245 ;
        RECT -19.885 2.555 -19.555 2.885 ;
        RECT -19.885 1.195 -19.555 1.525 ;
        RECT -19.885 -0.165 -19.555 0.165 ;
        RECT -19.885 -1.525 -19.555 -1.195 ;
        RECT -19.885 -2.885 -19.555 -2.555 ;
        RECT -19.885 -8.325 -19.555 -7.995 ;
        RECT -19.885 -9.685 -19.555 -9.355 ;
        RECT -19.885 -11.16 -19.555 -10.83 ;
        RECT -19.885 -12.405 -19.555 -12.075 ;
        RECT -19.885 -15.125 -19.555 -14.795 ;
        RECT -19.885 -16.25 -19.555 -15.92 ;
        RECT -19.88 -17.84 -19.56 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.885 -37.43 -19.555 -37.1 ;
        RECT -19.88 -39.6 -19.56 -34.52 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.885 -108.965 -19.555 -108.635 ;
        RECT -19.885 -110.325 -19.555 -109.995 ;
        RECT -19.885 -111.685 -19.555 -111.355 ;
        RECT -19.885 -113.045 -19.555 -112.715 ;
        RECT -19.885 -115.765 -19.555 -115.435 ;
        RECT -19.885 -117.125 -19.555 -116.795 ;
        RECT -19.885 -118.485 -19.555 -118.155 ;
        RECT -19.885 -119.845 -19.555 -119.515 ;
        RECT -19.885 -121.205 -19.555 -120.875 ;
        RECT -19.885 -122.565 -19.555 -122.235 ;
        RECT -19.885 -124.39 -19.555 -124.06 ;
        RECT -19.885 -125.285 -19.555 -124.955 ;
        RECT -19.885 -126.645 -19.555 -126.315 ;
        RECT -19.885 -128.005 -19.555 -127.675 ;
        RECT -19.885 -129.365 -19.555 -129.035 ;
        RECT -19.885 -133.445 -19.555 -133.115 ;
        RECT -19.885 -134.805 -19.555 -134.475 ;
        RECT -19.885 -136.165 -19.555 -135.835 ;
        RECT -19.885 -137.525 -19.555 -137.195 ;
        RECT -19.885 -144.325 -19.555 -143.995 ;
        RECT -19.885 -147.045 -19.555 -146.715 ;
        RECT -19.885 -148.405 -19.555 -148.075 ;
        RECT -19.885 -149.765 -19.555 -149.435 ;
        RECT -19.885 -151.125 -19.555 -150.795 ;
        RECT -19.885 -152.485 -19.555 -152.155 ;
        RECT -19.885 -155.205 -19.555 -154.875 ;
        RECT -19.885 -156.565 -19.555 -156.235 ;
        RECT -19.885 -157.925 -19.555 -157.595 ;
        RECT -19.885 -159.285 -19.555 -158.955 ;
        RECT -19.885 -160.645 -19.555 -160.315 ;
        RECT -19.885 -162.005 -19.555 -161.675 ;
        RECT -19.885 -163.365 -19.555 -163.035 ;
        RECT -19.885 -172.885 -19.555 -172.555 ;
        RECT -19.885 -175.605 -19.555 -175.275 ;
        RECT -19.885 -176.965 -19.555 -176.635 ;
        RECT -19.885 -179.685 -19.555 -179.355 ;
        RECT -19.885 -182.405 -19.555 -182.075 ;
        RECT -19.885 -185.125 -19.555 -184.795 ;
        RECT -19.885 -189.205 -19.555 -188.875 ;
        RECT -19.885 -190.565 -19.555 -190.235 ;
        RECT -19.885 -194.645 -19.555 -194.315 ;
        RECT -19.885 -196.005 -19.555 -195.675 ;
        RECT -19.885 -197.365 -19.555 -197.035 ;
        RECT -19.885 -198.725 -19.555 -198.395 ;
        RECT -19.885 -200.085 -19.555 -199.755 ;
        RECT -19.885 -201.445 -19.555 -201.115 ;
        RECT -19.885 -202.805 -19.555 -202.475 ;
        RECT -19.885 -204.165 -19.555 -203.835 ;
        RECT -19.88 -204.165 -19.56 -107.28 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.885 -210.965 -19.555 -210.635 ;
        RECT -19.885 -212.325 -19.555 -211.995 ;
        RECT -19.885 -213.625 -19.555 -213.295 ;
        RECT -19.885 -215.045 -19.555 -214.715 ;
        RECT -19.885 -216.405 -19.555 -216.075 ;
        RECT -19.885 -217.765 -19.555 -217.435 ;
        RECT -19.885 -219.125 -19.555 -218.795 ;
        RECT -19.885 -221.37 -19.555 -220.24 ;
        RECT -19.88 -221.485 -19.56 -209.96 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.525 129.8 -18.195 130.93 ;
        RECT -18.525 127.675 -18.195 128.005 ;
        RECT -18.525 126.315 -18.195 126.645 ;
        RECT -18.525 124.955 -18.195 125.285 ;
        RECT -18.525 123.595 -18.195 123.925 ;
        RECT -18.525 122.235 -18.195 122.565 ;
        RECT -18.525 120.875 -18.195 121.205 ;
        RECT -18.525 119.515 -18.195 119.845 ;
        RECT -18.525 118.155 -18.195 118.485 ;
        RECT -18.525 116.795 -18.195 117.125 ;
        RECT -18.525 115.435 -18.195 115.765 ;
        RECT -18.525 114.075 -18.195 114.405 ;
        RECT -18.525 112.715 -18.195 113.045 ;
        RECT -18.525 111.355 -18.195 111.685 ;
        RECT -18.525 109.995 -18.195 110.325 ;
        RECT -18.525 108.635 -18.195 108.965 ;
        RECT -18.525 107.275 -18.195 107.605 ;
        RECT -18.525 105.915 -18.195 106.245 ;
        RECT -18.525 104.555 -18.195 104.885 ;
        RECT -18.525 103.195 -18.195 103.525 ;
        RECT -18.525 101.835 -18.195 102.165 ;
        RECT -18.525 100.475 -18.195 100.805 ;
        RECT -18.525 99.115 -18.195 99.445 ;
        RECT -18.525 97.755 -18.195 98.085 ;
        RECT -18.525 96.395 -18.195 96.725 ;
        RECT -18.525 95.035 -18.195 95.365 ;
        RECT -18.525 93.675 -18.195 94.005 ;
        RECT -18.525 92.315 -18.195 92.645 ;
        RECT -18.525 90.955 -18.195 91.285 ;
        RECT -18.525 89.595 -18.195 89.925 ;
        RECT -18.525 88.235 -18.195 88.565 ;
        RECT -18.525 86.875 -18.195 87.205 ;
        RECT -18.525 85.515 -18.195 85.845 ;
        RECT -18.525 84.155 -18.195 84.485 ;
        RECT -18.525 82.795 -18.195 83.125 ;
        RECT -18.525 81.435 -18.195 81.765 ;
        RECT -18.525 80.075 -18.195 80.405 ;
        RECT -18.525 78.715 -18.195 79.045 ;
        RECT -18.525 77.355 -18.195 77.685 ;
        RECT -18.525 75.995 -18.195 76.325 ;
        RECT -18.525 74.635 -18.195 74.965 ;
        RECT -18.525 73.275 -18.195 73.605 ;
        RECT -18.525 71.915 -18.195 72.245 ;
        RECT -18.525 70.555 -18.195 70.885 ;
        RECT -18.525 69.195 -18.195 69.525 ;
        RECT -18.525 67.835 -18.195 68.165 ;
        RECT -18.525 66.475 -18.195 66.805 ;
        RECT -18.525 65.115 -18.195 65.445 ;
        RECT -18.525 63.755 -18.195 64.085 ;
        RECT -18.525 62.395 -18.195 62.725 ;
        RECT -18.525 61.035 -18.195 61.365 ;
        RECT -18.525 59.675 -18.195 60.005 ;
        RECT -18.525 58.315 -18.195 58.645 ;
        RECT -18.525 56.955 -18.195 57.285 ;
        RECT -18.525 55.595 -18.195 55.925 ;
        RECT -18.525 54.235 -18.195 54.565 ;
        RECT -18.525 52.875 -18.195 53.205 ;
        RECT -18.525 51.515 -18.195 51.845 ;
        RECT -18.525 50.155 -18.195 50.485 ;
        RECT -18.525 48.795 -18.195 49.125 ;
        RECT -18.525 47.435 -18.195 47.765 ;
        RECT -18.525 46.075 -18.195 46.405 ;
        RECT -18.525 44.715 -18.195 45.045 ;
        RECT -18.525 43.355 -18.195 43.685 ;
        RECT -18.525 41.995 -18.195 42.325 ;
        RECT -18.525 40.635 -18.195 40.965 ;
        RECT -18.525 39.275 -18.195 39.605 ;
        RECT -18.525 37.915 -18.195 38.245 ;
        RECT -18.525 36.555 -18.195 36.885 ;
        RECT -18.525 35.195 -18.195 35.525 ;
        RECT -18.525 33.835 -18.195 34.165 ;
        RECT -18.525 32.475 -18.195 32.805 ;
        RECT -18.525 31.115 -18.195 31.445 ;
        RECT -18.525 29.755 -18.195 30.085 ;
        RECT -18.525 28.395 -18.195 28.725 ;
        RECT -18.525 27.035 -18.195 27.365 ;
        RECT -18.525 25.675 -18.195 26.005 ;
        RECT -18.525 24.315 -18.195 24.645 ;
        RECT -18.525 22.955 -18.195 23.285 ;
        RECT -18.525 21.595 -18.195 21.925 ;
        RECT -18.525 20.235 -18.195 20.565 ;
        RECT -18.525 18.875 -18.195 19.205 ;
        RECT -18.525 17.515 -18.195 17.845 ;
        RECT -18.525 16.155 -18.195 16.485 ;
        RECT -18.525 14.795 -18.195 15.125 ;
        RECT -18.525 13.435 -18.195 13.765 ;
        RECT -18.525 12.075 -18.195 12.405 ;
        RECT -18.525 10.715 -18.195 11.045 ;
        RECT -18.525 9.355 -18.195 9.685 ;
        RECT -18.525 7.995 -18.195 8.325 ;
        RECT -18.525 6.635 -18.195 6.965 ;
        RECT -18.525 5.275 -18.195 5.605 ;
        RECT -18.525 3.915 -18.195 4.245 ;
        RECT -18.525 2.555 -18.195 2.885 ;
        RECT -18.525 1.195 -18.195 1.525 ;
        RECT -18.525 -0.165 -18.195 0.165 ;
        RECT -18.525 -1.525 -18.195 -1.195 ;
        RECT -18.525 -2.885 -18.195 -2.555 ;
        RECT -18.525 -8.325 -18.195 -7.995 ;
        RECT -18.525 -9.685 -18.195 -9.355 ;
        RECT -18.525 -11.16 -18.195 -10.83 ;
        RECT -18.525 -12.405 -18.195 -12.075 ;
        RECT -18.525 -15.125 -18.195 -14.795 ;
        RECT -18.525 -16.25 -18.195 -15.92 ;
        RECT -18.52 -17.16 -18.2 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.525 -108.965 -18.195 -108.635 ;
        RECT -18.525 -110.325 -18.195 -109.995 ;
        RECT -18.525 -111.685 -18.195 -111.355 ;
        RECT -18.525 -113.045 -18.195 -112.715 ;
        RECT -18.525 -115.765 -18.195 -115.435 ;
        RECT -18.525 -117.125 -18.195 -116.795 ;
        RECT -18.525 -118.485 -18.195 -118.155 ;
        RECT -18.525 -119.845 -18.195 -119.515 ;
        RECT -18.525 -121.205 -18.195 -120.875 ;
        RECT -18.525 -122.565 -18.195 -122.235 ;
        RECT -18.525 -124.39 -18.195 -124.06 ;
        RECT -18.525 -125.285 -18.195 -124.955 ;
        RECT -18.525 -126.645 -18.195 -126.315 ;
        RECT -18.525 -128.005 -18.195 -127.675 ;
        RECT -18.525 -129.365 -18.195 -129.035 ;
        RECT -18.525 -133.445 -18.195 -133.115 ;
        RECT -18.525 -134.805 -18.195 -134.475 ;
        RECT -18.525 -136.165 -18.195 -135.835 ;
        RECT -18.525 -137.525 -18.195 -137.195 ;
        RECT -18.525 -148.405 -18.195 -148.075 ;
        RECT -18.525 -149.765 -18.195 -149.435 ;
        RECT -18.525 -151.125 -18.195 -150.795 ;
        RECT -18.525 -152.485 -18.195 -152.155 ;
        RECT -18.525 -155.205 -18.195 -154.875 ;
        RECT -18.525 -156.565 -18.195 -156.235 ;
        RECT -18.525 -157.925 -18.195 -157.595 ;
        RECT -18.525 -159.285 -18.195 -158.955 ;
        RECT -18.525 -160.645 -18.195 -160.315 ;
        RECT -18.525 -162.005 -18.195 -161.675 ;
        RECT -18.525 -163.365 -18.195 -163.035 ;
        RECT -18.525 -172.885 -18.195 -172.555 ;
        RECT -18.525 -175.605 -18.195 -175.275 ;
        RECT -18.525 -176.965 -18.195 -176.635 ;
        RECT -18.525 -182.405 -18.195 -182.075 ;
        RECT -18.525 -189.205 -18.195 -188.875 ;
        RECT -18.525 -190.565 -18.195 -190.235 ;
        RECT -18.525 -194.645 -18.195 -194.315 ;
        RECT -18.525 -196.005 -18.195 -195.675 ;
        RECT -18.525 -197.365 -18.195 -197.035 ;
        RECT -18.525 -198.725 -18.195 -198.395 ;
        RECT -18.525 -200.085 -18.195 -199.755 ;
        RECT -18.525 -201.445 -18.195 -201.115 ;
        RECT -18.525 -202.805 -18.195 -202.475 ;
        RECT -18.525 -204.165 -18.195 -203.835 ;
        RECT -18.525 -205.525 -18.195 -205.195 ;
        RECT -18.525 -208.245 -18.195 -207.915 ;
        RECT -18.525 -210.965 -18.195 -210.635 ;
        RECT -18.525 -212.325 -18.195 -211.995 ;
        RECT -18.525 -213.625 -18.195 -213.295 ;
        RECT -18.525 -215.045 -18.195 -214.715 ;
        RECT -18.525 -216.405 -18.195 -216.075 ;
        RECT -18.525 -217.765 -18.195 -217.435 ;
        RECT -18.525 -219.125 -18.195 -218.795 ;
        RECT -18.525 -221.37 -18.195 -220.24 ;
        RECT -18.52 -221.485 -18.2 -108.635 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.165 129.8 -16.835 130.93 ;
        RECT -17.165 127.675 -16.835 128.005 ;
        RECT -17.165 126.315 -16.835 126.645 ;
        RECT -17.165 124.955 -16.835 125.285 ;
        RECT -17.165 123.595 -16.835 123.925 ;
        RECT -17.165 122.235 -16.835 122.565 ;
        RECT -17.165 120.875 -16.835 121.205 ;
        RECT -17.165 119.515 -16.835 119.845 ;
        RECT -17.165 118.155 -16.835 118.485 ;
        RECT -17.165 116.795 -16.835 117.125 ;
        RECT -17.165 115.435 -16.835 115.765 ;
        RECT -17.165 114.075 -16.835 114.405 ;
        RECT -17.165 112.715 -16.835 113.045 ;
        RECT -17.165 111.355 -16.835 111.685 ;
        RECT -17.165 109.995 -16.835 110.325 ;
        RECT -17.165 108.635 -16.835 108.965 ;
        RECT -17.165 107.275 -16.835 107.605 ;
        RECT -17.165 105.915 -16.835 106.245 ;
        RECT -17.165 104.555 -16.835 104.885 ;
        RECT -17.165 103.195 -16.835 103.525 ;
        RECT -17.165 101.835 -16.835 102.165 ;
        RECT -17.165 100.475 -16.835 100.805 ;
        RECT -17.165 99.115 -16.835 99.445 ;
        RECT -17.165 97.755 -16.835 98.085 ;
        RECT -17.165 96.395 -16.835 96.725 ;
        RECT -17.165 95.035 -16.835 95.365 ;
        RECT -17.165 93.675 -16.835 94.005 ;
        RECT -17.165 92.315 -16.835 92.645 ;
        RECT -17.165 90.955 -16.835 91.285 ;
        RECT -17.165 89.595 -16.835 89.925 ;
        RECT -17.165 88.235 -16.835 88.565 ;
        RECT -17.165 86.875 -16.835 87.205 ;
        RECT -17.165 85.515 -16.835 85.845 ;
        RECT -17.165 84.155 -16.835 84.485 ;
        RECT -17.165 82.795 -16.835 83.125 ;
        RECT -17.165 81.435 -16.835 81.765 ;
        RECT -17.165 80.075 -16.835 80.405 ;
        RECT -17.165 78.715 -16.835 79.045 ;
        RECT -17.165 77.355 -16.835 77.685 ;
        RECT -17.165 75.995 -16.835 76.325 ;
        RECT -17.165 74.635 -16.835 74.965 ;
        RECT -17.165 73.275 -16.835 73.605 ;
        RECT -17.165 71.915 -16.835 72.245 ;
        RECT -17.165 70.555 -16.835 70.885 ;
        RECT -17.165 69.195 -16.835 69.525 ;
        RECT -17.165 67.835 -16.835 68.165 ;
        RECT -17.165 66.475 -16.835 66.805 ;
        RECT -17.165 65.115 -16.835 65.445 ;
        RECT -17.165 63.755 -16.835 64.085 ;
        RECT -17.165 62.395 -16.835 62.725 ;
        RECT -17.165 61.035 -16.835 61.365 ;
        RECT -17.165 59.675 -16.835 60.005 ;
        RECT -17.165 58.315 -16.835 58.645 ;
        RECT -17.165 56.955 -16.835 57.285 ;
        RECT -17.165 55.595 -16.835 55.925 ;
        RECT -17.165 54.235 -16.835 54.565 ;
        RECT -17.165 52.875 -16.835 53.205 ;
        RECT -17.165 51.515 -16.835 51.845 ;
        RECT -17.165 50.155 -16.835 50.485 ;
        RECT -17.165 48.795 -16.835 49.125 ;
        RECT -17.165 47.435 -16.835 47.765 ;
        RECT -17.165 46.075 -16.835 46.405 ;
        RECT -17.165 44.715 -16.835 45.045 ;
        RECT -17.165 43.355 -16.835 43.685 ;
        RECT -17.165 41.995 -16.835 42.325 ;
        RECT -17.165 40.635 -16.835 40.965 ;
        RECT -17.165 39.275 -16.835 39.605 ;
        RECT -17.165 37.915 -16.835 38.245 ;
        RECT -17.165 36.555 -16.835 36.885 ;
        RECT -17.165 35.195 -16.835 35.525 ;
        RECT -17.165 33.835 -16.835 34.165 ;
        RECT -17.165 32.475 -16.835 32.805 ;
        RECT -17.165 31.115 -16.835 31.445 ;
        RECT -17.165 29.755 -16.835 30.085 ;
        RECT -17.165 28.395 -16.835 28.725 ;
        RECT -17.165 27.035 -16.835 27.365 ;
        RECT -17.165 25.675 -16.835 26.005 ;
        RECT -17.165 24.315 -16.835 24.645 ;
        RECT -17.165 22.955 -16.835 23.285 ;
        RECT -17.165 21.595 -16.835 21.925 ;
        RECT -17.165 20.235 -16.835 20.565 ;
        RECT -17.165 18.875 -16.835 19.205 ;
        RECT -17.165 17.515 -16.835 17.845 ;
        RECT -17.165 16.155 -16.835 16.485 ;
        RECT -17.165 14.795 -16.835 15.125 ;
        RECT -17.165 13.435 -16.835 13.765 ;
        RECT -17.165 12.075 -16.835 12.405 ;
        RECT -17.165 10.715 -16.835 11.045 ;
        RECT -17.165 9.355 -16.835 9.685 ;
        RECT -17.165 7.995 -16.835 8.325 ;
        RECT -17.165 6.635 -16.835 6.965 ;
        RECT -17.165 5.275 -16.835 5.605 ;
        RECT -17.165 3.915 -16.835 4.245 ;
        RECT -17.165 2.555 -16.835 2.885 ;
        RECT -17.165 1.195 -16.835 1.525 ;
        RECT -17.165 -0.165 -16.835 0.165 ;
        RECT -17.165 -1.525 -16.835 -1.195 ;
        RECT -17.165 -2.885 -16.835 -2.555 ;
        RECT -17.165 -8.325 -16.835 -7.995 ;
        RECT -17.165 -9.685 -16.835 -9.355 ;
        RECT -17.165 -11.16 -16.835 -10.83 ;
        RECT -17.165 -12.405 -16.835 -12.075 ;
        RECT -17.165 -15.125 -16.835 -14.795 ;
        RECT -17.165 -16.25 -16.835 -15.92 ;
        RECT -17.165 -21.925 -16.835 -21.595 ;
        RECT -17.165 -23.285 -16.835 -22.955 ;
        RECT -17.165 -27.365 -16.835 -27.035 ;
        RECT -17.165 -30.085 -16.835 -29.755 ;
        RECT -17.165 -31.445 -16.835 -31.115 ;
        RECT -17.165 -32.34 -16.835 -32.01 ;
        RECT -17.165 -34.165 -16.835 -33.835 ;
        RECT -17.165 -37.43 -16.835 -37.1 ;
        RECT -17.165 -38.245 -16.835 -37.915 ;
        RECT -17.165 -43.685 -16.835 -43.355 ;
        RECT -17.165 -45.045 -16.835 -44.715 ;
        RECT -17.165 -46.405 -16.835 -46.075 ;
        RECT -17.165 -47.765 -16.835 -47.435 ;
        RECT -17.165 -49.125 -16.835 -48.795 ;
        RECT -17.165 -50.485 -16.835 -50.155 ;
        RECT -17.165 -53.205 -16.835 -52.875 ;
        RECT -17.165 -54.565 -16.835 -54.235 ;
        RECT -17.165 -55.925 -16.835 -55.595 ;
        RECT -17.165 -57.285 -16.835 -56.955 ;
        RECT -17.165 -58.645 -16.835 -58.315 ;
        RECT -17.165 -60.005 -16.835 -59.675 ;
        RECT -17.165 -61.67 -16.835 -61.34 ;
        RECT -17.165 -65.445 -16.835 -65.115 ;
        RECT -17.165 -66.805 -16.835 -66.475 ;
        RECT -17.165 -68.165 -16.835 -67.835 ;
        RECT -17.165 -69.525 -16.835 -69.195 ;
        RECT -17.165 -72.245 -16.835 -71.915 ;
        RECT -17.165 -73.605 -16.835 -73.275 ;
        RECT -17.165 -74.965 -16.835 -74.635 ;
        RECT -17.165 -76.325 -16.835 -75.995 ;
        RECT -17.165 -77.685 -16.835 -77.355 ;
        RECT -17.165 -79.045 -16.835 -78.715 ;
        RECT -17.165 -80.21 -16.835 -79.88 ;
        RECT -17.165 -81.765 -16.835 -81.435 ;
        RECT -17.165 -83.125 -16.835 -82.795 ;
        RECT -17.165 -84.485 -16.835 -84.155 ;
        RECT -17.165 -87.205 -16.835 -86.875 ;
        RECT -17.165 -88.565 -16.835 -88.235 ;
        RECT -17.165 -89.925 -16.835 -89.595 ;
        RECT -17.165 -91.285 -16.835 -90.955 ;
        RECT -17.165 -92.645 -16.835 -92.315 ;
        RECT -17.165 -94.005 -16.835 -93.675 ;
        RECT -17.165 -95.365 -16.835 -95.035 ;
        RECT -17.165 -98.085 -16.835 -97.755 ;
        RECT -17.165 -99.445 -16.835 -99.115 ;
        RECT -17.165 -100.805 -16.835 -100.475 ;
        RECT -17.165 -102.165 -16.835 -101.835 ;
        RECT -17.165 -103.525 -16.835 -103.195 ;
        RECT -17.165 -104.885 -16.835 -104.555 ;
        RECT -17.165 -105.85 -16.835 -105.52 ;
        RECT -17.165 -107.605 -16.835 -107.275 ;
        RECT -17.165 -108.965 -16.835 -108.635 ;
        RECT -17.165 -110.325 -16.835 -109.995 ;
        RECT -17.165 -111.685 -16.835 -111.355 ;
        RECT -17.165 -113.045 -16.835 -112.715 ;
        RECT -17.165 -115.765 -16.835 -115.435 ;
        RECT -17.165 -117.125 -16.835 -116.795 ;
        RECT -17.165 -118.485 -16.835 -118.155 ;
        RECT -17.165 -119.845 -16.835 -119.515 ;
        RECT -17.165 -121.205 -16.835 -120.875 ;
        RECT -17.165 -122.565 -16.835 -122.235 ;
        RECT -17.165 -124.39 -16.835 -124.06 ;
        RECT -17.165 -125.285 -16.835 -124.955 ;
        RECT -17.165 -126.645 -16.835 -126.315 ;
        RECT -17.165 -128.005 -16.835 -127.675 ;
        RECT -17.165 -129.365 -16.835 -129.035 ;
        RECT -17.165 -133.445 -16.835 -133.115 ;
        RECT -17.165 -134.805 -16.835 -134.475 ;
        RECT -17.165 -136.165 -16.835 -135.835 ;
        RECT -17.165 -137.525 -16.835 -137.195 ;
        RECT -17.165 -148.405 -16.835 -148.075 ;
        RECT -17.165 -149.765 -16.835 -149.435 ;
        RECT -17.165 -151.125 -16.835 -150.795 ;
        RECT -17.165 -152.485 -16.835 -152.155 ;
        RECT -17.165 -155.205 -16.835 -154.875 ;
        RECT -17.165 -156.565 -16.835 -156.235 ;
        RECT -17.165 -157.925 -16.835 -157.595 ;
        RECT -17.165 -159.285 -16.835 -158.955 ;
        RECT -17.165 -160.645 -16.835 -160.315 ;
        RECT -17.165 -162.005 -16.835 -161.675 ;
        RECT -17.165 -163.365 -16.835 -163.035 ;
        RECT -17.165 -175.605 -16.835 -175.275 ;
        RECT -17.165 -176.965 -16.835 -176.635 ;
        RECT -17.165 -182.405 -16.835 -182.075 ;
        RECT -17.165 -183.765 -16.835 -183.435 ;
        RECT -17.165 -189.205 -16.835 -188.875 ;
        RECT -17.165 -190.565 -16.835 -190.235 ;
        RECT -17.165 -194.645 -16.835 -194.315 ;
        RECT -17.165 -196.005 -16.835 -195.675 ;
        RECT -17.165 -197.365 -16.835 -197.035 ;
        RECT -17.165 -198.725 -16.835 -198.395 ;
        RECT -17.165 -200.085 -16.835 -199.755 ;
        RECT -17.165 -201.445 -16.835 -201.115 ;
        RECT -17.165 -202.805 -16.835 -202.475 ;
        RECT -17.165 -204.165 -16.835 -203.835 ;
        RECT -17.165 -205.525 -16.835 -205.195 ;
        RECT -17.16 -206.88 -16.84 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.165 -212.325 -16.835 -211.995 ;
        RECT -17.165 -213.625 -16.835 -213.295 ;
        RECT -17.165 -215.045 -16.835 -214.715 ;
        RECT -17.165 -216.405 -16.835 -216.075 ;
        RECT -17.165 -217.765 -16.835 -217.435 ;
        RECT -17.165 -219.125 -16.835 -218.795 ;
        RECT -17.165 -221.37 -16.835 -220.24 ;
        RECT -17.16 -221.485 -16.84 -211.995 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.805 129.8 -15.475 130.93 ;
        RECT -15.805 127.675 -15.475 128.005 ;
        RECT -15.805 126.315 -15.475 126.645 ;
        RECT -15.805 124.955 -15.475 125.285 ;
        RECT -15.805 123.595 -15.475 123.925 ;
        RECT -15.805 122.235 -15.475 122.565 ;
        RECT -15.805 120.875 -15.475 121.205 ;
        RECT -15.805 119.515 -15.475 119.845 ;
        RECT -15.805 118.155 -15.475 118.485 ;
        RECT -15.805 116.795 -15.475 117.125 ;
        RECT -15.805 115.435 -15.475 115.765 ;
        RECT -15.805 114.075 -15.475 114.405 ;
        RECT -15.805 112.715 -15.475 113.045 ;
        RECT -15.805 111.355 -15.475 111.685 ;
        RECT -15.805 109.995 -15.475 110.325 ;
        RECT -15.805 108.635 -15.475 108.965 ;
        RECT -15.805 107.275 -15.475 107.605 ;
        RECT -15.805 105.915 -15.475 106.245 ;
        RECT -15.805 104.555 -15.475 104.885 ;
        RECT -15.805 103.195 -15.475 103.525 ;
        RECT -15.805 101.835 -15.475 102.165 ;
        RECT -15.805 100.475 -15.475 100.805 ;
        RECT -15.805 99.115 -15.475 99.445 ;
        RECT -15.805 97.755 -15.475 98.085 ;
        RECT -15.805 96.395 -15.475 96.725 ;
        RECT -15.805 95.035 -15.475 95.365 ;
        RECT -15.805 93.675 -15.475 94.005 ;
        RECT -15.805 92.315 -15.475 92.645 ;
        RECT -15.805 90.955 -15.475 91.285 ;
        RECT -15.805 89.595 -15.475 89.925 ;
        RECT -15.805 88.235 -15.475 88.565 ;
        RECT -15.805 86.875 -15.475 87.205 ;
        RECT -15.805 85.515 -15.475 85.845 ;
        RECT -15.805 84.155 -15.475 84.485 ;
        RECT -15.805 82.795 -15.475 83.125 ;
        RECT -15.805 81.435 -15.475 81.765 ;
        RECT -15.805 80.075 -15.475 80.405 ;
        RECT -15.805 78.715 -15.475 79.045 ;
        RECT -15.805 77.355 -15.475 77.685 ;
        RECT -15.805 75.995 -15.475 76.325 ;
        RECT -15.805 74.635 -15.475 74.965 ;
        RECT -15.805 73.275 -15.475 73.605 ;
        RECT -15.805 71.915 -15.475 72.245 ;
        RECT -15.805 70.555 -15.475 70.885 ;
        RECT -15.805 69.195 -15.475 69.525 ;
        RECT -15.805 67.835 -15.475 68.165 ;
        RECT -15.805 66.475 -15.475 66.805 ;
        RECT -15.805 65.115 -15.475 65.445 ;
        RECT -15.805 63.755 -15.475 64.085 ;
        RECT -15.805 62.395 -15.475 62.725 ;
        RECT -15.805 61.035 -15.475 61.365 ;
        RECT -15.805 59.675 -15.475 60.005 ;
        RECT -15.805 58.315 -15.475 58.645 ;
        RECT -15.805 56.955 -15.475 57.285 ;
        RECT -15.805 55.595 -15.475 55.925 ;
        RECT -15.805 54.235 -15.475 54.565 ;
        RECT -15.805 52.875 -15.475 53.205 ;
        RECT -15.805 51.515 -15.475 51.845 ;
        RECT -15.805 50.155 -15.475 50.485 ;
        RECT -15.805 48.795 -15.475 49.125 ;
        RECT -15.805 47.435 -15.475 47.765 ;
        RECT -15.805 46.075 -15.475 46.405 ;
        RECT -15.805 44.715 -15.475 45.045 ;
        RECT -15.805 43.355 -15.475 43.685 ;
        RECT -15.805 41.995 -15.475 42.325 ;
        RECT -15.805 40.635 -15.475 40.965 ;
        RECT -15.805 39.275 -15.475 39.605 ;
        RECT -15.805 37.915 -15.475 38.245 ;
        RECT -15.805 36.555 -15.475 36.885 ;
        RECT -15.805 35.195 -15.475 35.525 ;
        RECT -15.805 33.835 -15.475 34.165 ;
        RECT -15.805 32.475 -15.475 32.805 ;
        RECT -15.805 31.115 -15.475 31.445 ;
        RECT -15.805 29.755 -15.475 30.085 ;
        RECT -15.805 28.395 -15.475 28.725 ;
        RECT -15.805 27.035 -15.475 27.365 ;
        RECT -15.805 25.675 -15.475 26.005 ;
        RECT -15.805 24.315 -15.475 24.645 ;
        RECT -15.805 22.955 -15.475 23.285 ;
        RECT -15.805 21.595 -15.475 21.925 ;
        RECT -15.805 20.235 -15.475 20.565 ;
        RECT -15.805 18.875 -15.475 19.205 ;
        RECT -15.805 17.515 -15.475 17.845 ;
        RECT -15.805 16.155 -15.475 16.485 ;
        RECT -15.805 14.795 -15.475 15.125 ;
        RECT -15.805 13.435 -15.475 13.765 ;
        RECT -15.805 12.075 -15.475 12.405 ;
        RECT -15.805 10.715 -15.475 11.045 ;
        RECT -15.805 9.355 -15.475 9.685 ;
        RECT -15.805 7.995 -15.475 8.325 ;
        RECT -15.805 6.635 -15.475 6.965 ;
        RECT -15.805 5.275 -15.475 5.605 ;
        RECT -15.805 3.915 -15.475 4.245 ;
        RECT -15.805 2.555 -15.475 2.885 ;
        RECT -15.805 1.195 -15.475 1.525 ;
        RECT -15.805 -0.165 -15.475 0.165 ;
        RECT -15.805 -1.525 -15.475 -1.195 ;
        RECT -15.805 -2.885 -15.475 -2.555 ;
        RECT -15.805 -4.245 -15.475 -3.915 ;
        RECT -15.805 -8.325 -15.475 -7.995 ;
        RECT -15.805 -9.685 -15.475 -9.355 ;
        RECT -15.805 -11.16 -15.475 -10.83 ;
        RECT -15.805 -12.405 -15.475 -12.075 ;
        RECT -15.805 -15.125 -15.475 -14.795 ;
        RECT -15.805 -16.25 -15.475 -15.92 ;
        RECT -15.805 -21.925 -15.475 -21.595 ;
        RECT -15.805 -23.285 -15.475 -22.955 ;
        RECT -15.805 -24.645 -15.475 -24.315 ;
        RECT -15.805 -27.365 -15.475 -27.035 ;
        RECT -15.805 -30.085 -15.475 -29.755 ;
        RECT -15.805 -31.445 -15.475 -31.115 ;
        RECT -15.805 -32.34 -15.475 -32.01 ;
        RECT -15.805 -34.165 -15.475 -33.835 ;
        RECT -15.805 -37.43 -15.475 -37.1 ;
        RECT -15.805 -38.245 -15.475 -37.915 ;
        RECT -15.805 -43.685 -15.475 -43.355 ;
        RECT -15.805 -45.045 -15.475 -44.715 ;
        RECT -15.805 -46.405 -15.475 -46.075 ;
        RECT -15.805 -47.765 -15.475 -47.435 ;
        RECT -15.805 -49.125 -15.475 -48.795 ;
        RECT -15.805 -50.485 -15.475 -50.155 ;
        RECT -15.805 -53.205 -15.475 -52.875 ;
        RECT -15.805 -54.565 -15.475 -54.235 ;
        RECT -15.805 -55.925 -15.475 -55.595 ;
        RECT -15.805 -57.285 -15.475 -56.955 ;
        RECT -15.805 -58.645 -15.475 -58.315 ;
        RECT -15.805 -60.005 -15.475 -59.675 ;
        RECT -15.805 -61.67 -15.475 -61.34 ;
        RECT -15.805 -65.445 -15.475 -65.115 ;
        RECT -15.805 -66.805 -15.475 -66.475 ;
        RECT -15.805 -68.165 -15.475 -67.835 ;
        RECT -15.805 -69.525 -15.475 -69.195 ;
        RECT -15.805 -72.245 -15.475 -71.915 ;
        RECT -15.805 -73.605 -15.475 -73.275 ;
        RECT -15.805 -74.965 -15.475 -74.635 ;
        RECT -15.805 -76.325 -15.475 -75.995 ;
        RECT -15.805 -77.685 -15.475 -77.355 ;
        RECT -15.805 -79.045 -15.475 -78.715 ;
        RECT -15.805 -80.21 -15.475 -79.88 ;
        RECT -15.805 -81.765 -15.475 -81.435 ;
        RECT -15.805 -83.125 -15.475 -82.795 ;
        RECT -15.805 -84.485 -15.475 -84.155 ;
        RECT -15.805 -87.205 -15.475 -86.875 ;
        RECT -15.805 -88.565 -15.475 -88.235 ;
        RECT -15.805 -89.925 -15.475 -89.595 ;
        RECT -15.805 -91.285 -15.475 -90.955 ;
        RECT -15.805 -92.645 -15.475 -92.315 ;
        RECT -15.805 -94.005 -15.475 -93.675 ;
        RECT -15.805 -95.365 -15.475 -95.035 ;
        RECT -15.805 -98.085 -15.475 -97.755 ;
        RECT -15.805 -99.445 -15.475 -99.115 ;
        RECT -15.805 -100.805 -15.475 -100.475 ;
        RECT -15.805 -102.165 -15.475 -101.835 ;
        RECT -15.805 -103.525 -15.475 -103.195 ;
        RECT -15.805 -104.885 -15.475 -104.555 ;
        RECT -15.805 -105.85 -15.475 -105.52 ;
        RECT -15.805 -107.605 -15.475 -107.275 ;
        RECT -15.805 -108.965 -15.475 -108.635 ;
        RECT -15.805 -110.325 -15.475 -109.995 ;
        RECT -15.805 -111.685 -15.475 -111.355 ;
        RECT -15.805 -113.045 -15.475 -112.715 ;
        RECT -15.805 -115.765 -15.475 -115.435 ;
        RECT -15.805 -117.125 -15.475 -116.795 ;
        RECT -15.805 -118.485 -15.475 -118.155 ;
        RECT -15.805 -119.845 -15.475 -119.515 ;
        RECT -15.805 -121.205 -15.475 -120.875 ;
        RECT -15.805 -122.565 -15.475 -122.235 ;
        RECT -15.805 -124.39 -15.475 -124.06 ;
        RECT -15.805 -125.285 -15.475 -124.955 ;
        RECT -15.805 -126.645 -15.475 -126.315 ;
        RECT -15.805 -128.005 -15.475 -127.675 ;
        RECT -15.805 -129.365 -15.475 -129.035 ;
        RECT -15.8 -130.04 -15.48 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.805 -212.325 -15.475 -211.995 ;
        RECT -15.805 -213.625 -15.475 -213.295 ;
        RECT -15.805 -215.045 -15.475 -214.715 ;
        RECT -15.805 -216.405 -15.475 -216.075 ;
        RECT -15.805 -217.765 -15.475 -217.435 ;
        RECT -15.805 -219.125 -15.475 -218.795 ;
        RECT -15.805 -221.37 -15.475 -220.24 ;
        RECT -15.8 -221.485 -15.48 -208.6 ;
    END
    PORT
      LAYER met3 ;
        RECT -14.445 9.355 -14.115 9.685 ;
        RECT -14.445 7.995 -14.115 8.325 ;
        RECT -14.445 6.635 -14.115 6.965 ;
        RECT -14.445 5.275 -14.115 5.605 ;
        RECT -14.445 3.915 -14.115 4.245 ;
        RECT -14.445 2.555 -14.115 2.885 ;
        RECT -14.445 1.195 -14.115 1.525 ;
        RECT -14.445 -0.165 -14.115 0.165 ;
        RECT -14.445 -1.525 -14.115 -1.195 ;
        RECT -14.445 -2.885 -14.115 -2.555 ;
        RECT -14.445 -4.245 -14.115 -3.915 ;
        RECT -14.445 -8.325 -14.115 -7.995 ;
        RECT -14.445 -9.685 -14.115 -9.355 ;
        RECT -14.445 -11.16 -14.115 -10.83 ;
        RECT -14.445 -12.405 -14.115 -12.075 ;
        RECT -14.445 -15.125 -14.115 -14.795 ;
        RECT -14.445 -16.25 -14.115 -15.92 ;
        RECT -14.445 -21.925 -14.115 -21.595 ;
        RECT -14.445 -23.285 -14.115 -22.955 ;
        RECT -14.445 -24.645 -14.115 -24.315 ;
        RECT -14.445 -27.365 -14.115 -27.035 ;
        RECT -14.445 -30.085 -14.115 -29.755 ;
        RECT -14.445 -31.445 -14.115 -31.115 ;
        RECT -14.445 -32.34 -14.115 -32.01 ;
        RECT -14.445 -34.165 -14.115 -33.835 ;
        RECT -14.445 -37.43 -14.115 -37.1 ;
        RECT -14.445 -38.245 -14.115 -37.915 ;
        RECT -14.445 -43.685 -14.115 -43.355 ;
        RECT -14.445 -45.045 -14.115 -44.715 ;
        RECT -14.445 -46.405 -14.115 -46.075 ;
        RECT -14.445 -47.765 -14.115 -47.435 ;
        RECT -14.445 -49.125 -14.115 -48.795 ;
        RECT -14.445 -50.485 -14.115 -50.155 ;
        RECT -14.445 -53.205 -14.115 -52.875 ;
        RECT -14.445 -54.565 -14.115 -54.235 ;
        RECT -14.445 -55.925 -14.115 -55.595 ;
        RECT -14.445 -57.285 -14.115 -56.955 ;
        RECT -14.445 -58.645 -14.115 -58.315 ;
        RECT -14.445 -60.005 -14.115 -59.675 ;
        RECT -14.445 -61.67 -14.115 -61.34 ;
        RECT -14.445 -65.445 -14.115 -65.115 ;
        RECT -14.445 -66.805 -14.115 -66.475 ;
        RECT -14.445 -68.165 -14.115 -67.835 ;
        RECT -14.445 -69.525 -14.115 -69.195 ;
        RECT -14.445 -72.245 -14.115 -71.915 ;
        RECT -14.445 -73.605 -14.115 -73.275 ;
        RECT -14.445 -74.965 -14.115 -74.635 ;
        RECT -14.445 -76.325 -14.115 -75.995 ;
        RECT -14.445 -77.685 -14.115 -77.355 ;
        RECT -14.445 -79.045 -14.115 -78.715 ;
        RECT -14.445 -80.21 -14.115 -79.88 ;
        RECT -14.445 -81.765 -14.115 -81.435 ;
        RECT -14.445 -83.125 -14.115 -82.795 ;
        RECT -14.445 -84.485 -14.115 -84.155 ;
        RECT -14.445 -87.205 -14.115 -86.875 ;
        RECT -14.445 -88.565 -14.115 -88.235 ;
        RECT -14.445 -89.925 -14.115 -89.595 ;
        RECT -14.445 -91.285 -14.115 -90.955 ;
        RECT -14.445 -92.645 -14.115 -92.315 ;
        RECT -14.445 -94.005 -14.115 -93.675 ;
        RECT -14.445 -95.365 -14.115 -95.035 ;
        RECT -14.445 -98.085 -14.115 -97.755 ;
        RECT -14.445 -99.445 -14.115 -99.115 ;
        RECT -14.445 -100.805 -14.115 -100.475 ;
        RECT -14.445 -102.165 -14.115 -101.835 ;
        RECT -14.445 -103.525 -14.115 -103.195 ;
        RECT -14.445 -104.885 -14.115 -104.555 ;
        RECT -14.445 -105.85 -14.115 -105.52 ;
        RECT -14.445 -107.605 -14.115 -107.275 ;
        RECT -14.445 -108.965 -14.115 -108.635 ;
        RECT -14.445 -110.325 -14.115 -109.995 ;
        RECT -14.445 -111.685 -14.115 -111.355 ;
        RECT -14.445 -113.045 -14.115 -112.715 ;
        RECT -14.445 -115.765 -14.115 -115.435 ;
        RECT -14.445 -117.125 -14.115 -116.795 ;
        RECT -14.445 -118.485 -14.115 -118.155 ;
        RECT -14.445 -119.845 -14.115 -119.515 ;
        RECT -14.445 -121.205 -14.115 -120.875 ;
        RECT -14.445 -122.565 -14.115 -122.235 ;
        RECT -14.445 -124.39 -14.115 -124.06 ;
        RECT -14.445 -125.285 -14.115 -124.955 ;
        RECT -14.445 -126.645 -14.115 -126.315 ;
        RECT -14.445 -128.005 -14.115 -127.675 ;
        RECT -14.445 -129.365 -14.115 -129.035 ;
        RECT -14.44 -129.365 -14.12 131.045 ;
        RECT -14.445 129.8 -14.115 130.93 ;
        RECT -14.445 127.675 -14.115 128.005 ;
        RECT -14.445 126.315 -14.115 126.645 ;
        RECT -14.445 124.955 -14.115 125.285 ;
        RECT -14.445 123.595 -14.115 123.925 ;
        RECT -14.445 122.235 -14.115 122.565 ;
        RECT -14.445 120.875 -14.115 121.205 ;
        RECT -14.445 119.515 -14.115 119.845 ;
        RECT -14.445 118.155 -14.115 118.485 ;
        RECT -14.445 116.795 -14.115 117.125 ;
        RECT -14.445 115.435 -14.115 115.765 ;
        RECT -14.445 114.075 -14.115 114.405 ;
        RECT -14.445 112.715 -14.115 113.045 ;
        RECT -14.445 111.355 -14.115 111.685 ;
        RECT -14.445 109.995 -14.115 110.325 ;
        RECT -14.445 108.635 -14.115 108.965 ;
        RECT -14.445 107.275 -14.115 107.605 ;
        RECT -14.445 105.915 -14.115 106.245 ;
        RECT -14.445 104.555 -14.115 104.885 ;
        RECT -14.445 103.195 -14.115 103.525 ;
        RECT -14.445 101.835 -14.115 102.165 ;
        RECT -14.445 100.475 -14.115 100.805 ;
        RECT -14.445 99.115 -14.115 99.445 ;
        RECT -14.445 97.755 -14.115 98.085 ;
        RECT -14.445 96.395 -14.115 96.725 ;
        RECT -14.445 95.035 -14.115 95.365 ;
        RECT -14.445 93.675 -14.115 94.005 ;
        RECT -14.445 92.315 -14.115 92.645 ;
        RECT -14.445 90.955 -14.115 91.285 ;
        RECT -14.445 89.595 -14.115 89.925 ;
        RECT -14.445 88.235 -14.115 88.565 ;
        RECT -14.445 86.875 -14.115 87.205 ;
        RECT -14.445 85.515 -14.115 85.845 ;
        RECT -14.445 84.155 -14.115 84.485 ;
        RECT -14.445 82.795 -14.115 83.125 ;
        RECT -14.445 81.435 -14.115 81.765 ;
        RECT -14.445 80.075 -14.115 80.405 ;
        RECT -14.445 78.715 -14.115 79.045 ;
        RECT -14.445 77.355 -14.115 77.685 ;
        RECT -14.445 75.995 -14.115 76.325 ;
        RECT -14.445 74.635 -14.115 74.965 ;
        RECT -14.445 73.275 -14.115 73.605 ;
        RECT -14.445 71.915 -14.115 72.245 ;
        RECT -14.445 70.555 -14.115 70.885 ;
        RECT -14.445 69.195 -14.115 69.525 ;
        RECT -14.445 67.835 -14.115 68.165 ;
        RECT -14.445 66.475 -14.115 66.805 ;
        RECT -14.445 65.115 -14.115 65.445 ;
        RECT -14.445 63.755 -14.115 64.085 ;
        RECT -14.445 62.395 -14.115 62.725 ;
        RECT -14.445 61.035 -14.115 61.365 ;
        RECT -14.445 59.675 -14.115 60.005 ;
        RECT -14.445 58.315 -14.115 58.645 ;
        RECT -14.445 56.955 -14.115 57.285 ;
        RECT -14.445 55.595 -14.115 55.925 ;
        RECT -14.445 54.235 -14.115 54.565 ;
        RECT -14.445 52.875 -14.115 53.205 ;
        RECT -14.445 51.515 -14.115 51.845 ;
        RECT -14.445 50.155 -14.115 50.485 ;
        RECT -14.445 48.795 -14.115 49.125 ;
        RECT -14.445 47.435 -14.115 47.765 ;
        RECT -14.445 46.075 -14.115 46.405 ;
        RECT -14.445 44.715 -14.115 45.045 ;
        RECT -14.445 43.355 -14.115 43.685 ;
        RECT -14.445 41.995 -14.115 42.325 ;
        RECT -14.445 40.635 -14.115 40.965 ;
        RECT -14.445 39.275 -14.115 39.605 ;
        RECT -14.445 37.915 -14.115 38.245 ;
        RECT -14.445 36.555 -14.115 36.885 ;
        RECT -14.445 35.195 -14.115 35.525 ;
        RECT -14.445 33.835 -14.115 34.165 ;
        RECT -14.445 32.475 -14.115 32.805 ;
        RECT -14.445 31.115 -14.115 31.445 ;
        RECT -14.445 29.755 -14.115 30.085 ;
        RECT -14.445 28.395 -14.115 28.725 ;
        RECT -14.445 27.035 -14.115 27.365 ;
        RECT -14.445 25.675 -14.115 26.005 ;
        RECT -14.445 24.315 -14.115 24.645 ;
        RECT -14.445 22.955 -14.115 23.285 ;
        RECT -14.445 21.595 -14.115 21.925 ;
        RECT -14.445 20.235 -14.115 20.565 ;
        RECT -14.445 18.875 -14.115 19.205 ;
        RECT -14.445 17.515 -14.115 17.845 ;
        RECT -14.445 16.155 -14.115 16.485 ;
        RECT -14.445 14.795 -14.115 15.125 ;
        RECT -14.445 13.435 -14.115 13.765 ;
        RECT -14.445 12.075 -14.115 12.405 ;
        RECT -14.445 10.715 -14.115 11.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.685 129.8 -26.355 130.93 ;
        RECT -26.685 127.675 -26.355 128.005 ;
        RECT -26.685 126.315 -26.355 126.645 ;
        RECT -26.685 124.955 -26.355 125.285 ;
        RECT -26.685 123.595 -26.355 123.925 ;
        RECT -26.685 122.235 -26.355 122.565 ;
        RECT -26.685 120.875 -26.355 121.205 ;
        RECT -26.685 119.515 -26.355 119.845 ;
        RECT -26.685 118.155 -26.355 118.485 ;
        RECT -26.685 116.795 -26.355 117.125 ;
        RECT -26.685 115.435 -26.355 115.765 ;
        RECT -26.685 114.075 -26.355 114.405 ;
        RECT -26.685 112.715 -26.355 113.045 ;
        RECT -26.685 111.355 -26.355 111.685 ;
        RECT -26.685 109.995 -26.355 110.325 ;
        RECT -26.685 108.635 -26.355 108.965 ;
        RECT -26.685 107.275 -26.355 107.605 ;
        RECT -26.685 105.915 -26.355 106.245 ;
        RECT -26.685 104.555 -26.355 104.885 ;
        RECT -26.685 103.195 -26.355 103.525 ;
        RECT -26.685 101.835 -26.355 102.165 ;
        RECT -26.685 100.475 -26.355 100.805 ;
        RECT -26.685 99.115 -26.355 99.445 ;
        RECT -26.685 97.755 -26.355 98.085 ;
        RECT -26.685 96.395 -26.355 96.725 ;
        RECT -26.685 95.035 -26.355 95.365 ;
        RECT -26.685 93.675 -26.355 94.005 ;
        RECT -26.685 92.315 -26.355 92.645 ;
        RECT -26.685 90.955 -26.355 91.285 ;
        RECT -26.685 89.595 -26.355 89.925 ;
        RECT -26.685 88.235 -26.355 88.565 ;
        RECT -26.685 86.875 -26.355 87.205 ;
        RECT -26.685 85.515 -26.355 85.845 ;
        RECT -26.685 84.155 -26.355 84.485 ;
        RECT -26.685 82.795 -26.355 83.125 ;
        RECT -26.685 81.435 -26.355 81.765 ;
        RECT -26.685 80.075 -26.355 80.405 ;
        RECT -26.685 78.715 -26.355 79.045 ;
        RECT -26.685 77.355 -26.355 77.685 ;
        RECT -26.685 75.995 -26.355 76.325 ;
        RECT -26.685 74.635 -26.355 74.965 ;
        RECT -26.685 73.275 -26.355 73.605 ;
        RECT -26.685 71.915 -26.355 72.245 ;
        RECT -26.685 70.555 -26.355 70.885 ;
        RECT -26.685 69.195 -26.355 69.525 ;
        RECT -26.685 67.835 -26.355 68.165 ;
        RECT -26.685 66.475 -26.355 66.805 ;
        RECT -26.685 65.115 -26.355 65.445 ;
        RECT -26.685 63.755 -26.355 64.085 ;
        RECT -26.685 62.395 -26.355 62.725 ;
        RECT -26.685 61.035 -26.355 61.365 ;
        RECT -26.685 59.675 -26.355 60.005 ;
        RECT -26.685 58.315 -26.355 58.645 ;
        RECT -26.685 56.955 -26.355 57.285 ;
        RECT -26.685 55.595 -26.355 55.925 ;
        RECT -26.685 54.235 -26.355 54.565 ;
        RECT -26.685 52.875 -26.355 53.205 ;
        RECT -26.685 51.515 -26.355 51.845 ;
        RECT -26.685 50.155 -26.355 50.485 ;
        RECT -26.685 48.795 -26.355 49.125 ;
        RECT -26.685 47.435 -26.355 47.765 ;
        RECT -26.685 46.075 -26.355 46.405 ;
        RECT -26.685 44.715 -26.355 45.045 ;
        RECT -26.685 43.355 -26.355 43.685 ;
        RECT -26.685 41.995 -26.355 42.325 ;
        RECT -26.685 40.635 -26.355 40.965 ;
        RECT -26.685 39.275 -26.355 39.605 ;
        RECT -26.685 37.915 -26.355 38.245 ;
        RECT -26.685 36.555 -26.355 36.885 ;
        RECT -26.685 35.195 -26.355 35.525 ;
        RECT -26.685 33.835 -26.355 34.165 ;
        RECT -26.685 32.475 -26.355 32.805 ;
        RECT -26.685 31.115 -26.355 31.445 ;
        RECT -26.685 29.755 -26.355 30.085 ;
        RECT -26.685 28.395 -26.355 28.725 ;
        RECT -26.685 27.035 -26.355 27.365 ;
        RECT -26.685 25.675 -26.355 26.005 ;
        RECT -26.685 24.315 -26.355 24.645 ;
        RECT -26.685 22.955 -26.355 23.285 ;
        RECT -26.685 21.595 -26.355 21.925 ;
        RECT -26.685 20.235 -26.355 20.565 ;
        RECT -26.685 18.875 -26.355 19.205 ;
        RECT -26.685 17.515 -26.355 17.845 ;
        RECT -26.685 16.155 -26.355 16.485 ;
        RECT -26.685 14.795 -26.355 15.125 ;
        RECT -26.685 13.435 -26.355 13.765 ;
        RECT -26.685 12.075 -26.355 12.405 ;
        RECT -26.685 10.715 -26.355 11.045 ;
        RECT -26.685 9.355 -26.355 9.685 ;
        RECT -26.685 7.995 -26.355 8.325 ;
        RECT -26.685 6.635 -26.355 6.965 ;
        RECT -26.685 5.275 -26.355 5.605 ;
        RECT -26.685 3.915 -26.355 4.245 ;
        RECT -26.685 2.555 -26.355 2.885 ;
        RECT -26.685 1.195 -26.355 1.525 ;
        RECT -26.685 -0.165 -26.355 0.165 ;
        RECT -26.685 -8.325 -26.355 -7.995 ;
        RECT -26.685 -9.685 -26.355 -9.355 ;
        RECT -26.685 -11.16 -26.355 -10.83 ;
        RECT -26.685 -12.405 -26.355 -12.075 ;
        RECT -26.685 -15.125 -26.355 -14.795 ;
        RECT -26.685 -16.25 -26.355 -15.92 ;
        RECT -26.685 -27.365 -26.355 -27.035 ;
        RECT -26.685 -30.085 -26.355 -29.755 ;
        RECT -26.685 -32.34 -26.355 -32.01 ;
        RECT -26.685 -37.43 -26.355 -37.1 ;
        RECT -26.685 -43.685 -26.355 -43.355 ;
        RECT -26.685 -45.045 -26.355 -44.715 ;
        RECT -26.685 -46.405 -26.355 -46.075 ;
        RECT -26.685 -47.765 -26.355 -47.435 ;
        RECT -26.685 -49.125 -26.355 -48.795 ;
        RECT -26.685 -50.485 -26.355 -50.155 ;
        RECT -26.685 -51.845 -26.355 -51.515 ;
        RECT -26.685 -53.205 -26.355 -52.875 ;
        RECT -26.685 -54.565 -26.355 -54.235 ;
        RECT -26.685 -55.925 -26.355 -55.595 ;
        RECT -26.685 -57.285 -26.355 -56.955 ;
        RECT -26.685 -58.645 -26.355 -58.315 ;
        RECT -26.685 -60.005 -26.355 -59.675 ;
        RECT -26.685 -61.365 -26.355 -61.035 ;
        RECT -26.685 -62.725 -26.355 -62.395 ;
        RECT -26.685 -64.085 -26.355 -63.755 ;
        RECT -26.685 -65.445 -26.355 -65.115 ;
        RECT -26.685 -66.805 -26.355 -66.475 ;
        RECT -26.685 -68.165 -26.355 -67.835 ;
        RECT -26.685 -69.525 -26.355 -69.195 ;
        RECT -26.685 -70.885 -26.355 -70.555 ;
        RECT -26.685 -72.245 -26.355 -71.915 ;
        RECT -26.685 -73.605 -26.355 -73.275 ;
        RECT -26.685 -74.965 -26.355 -74.635 ;
        RECT -26.685 -76.325 -26.355 -75.995 ;
        RECT -26.685 -77.685 -26.355 -77.355 ;
        RECT -26.685 -79.045 -26.355 -78.715 ;
        RECT -26.685 -80.405 -26.355 -80.075 ;
        RECT -26.685 -81.765 -26.355 -81.435 ;
        RECT -26.685 -83.125 -26.355 -82.795 ;
        RECT -26.685 -84.485 -26.355 -84.155 ;
        RECT -26.685 -85.845 -26.355 -85.515 ;
        RECT -26.685 -87.205 -26.355 -86.875 ;
        RECT -26.685 -88.565 -26.355 -88.235 ;
        RECT -26.685 -89.925 -26.355 -89.595 ;
        RECT -26.685 -91.285 -26.355 -90.955 ;
        RECT -26.685 -92.645 -26.355 -92.315 ;
        RECT -26.685 -94.005 -26.355 -93.675 ;
        RECT -26.685 -95.365 -26.355 -95.035 ;
        RECT -26.685 -96.725 -26.355 -96.395 ;
        RECT -26.685 -98.085 -26.355 -97.755 ;
        RECT -26.685 -99.445 -26.355 -99.115 ;
        RECT -26.685 -100.805 -26.355 -100.475 ;
        RECT -26.685 -102.165 -26.355 -101.835 ;
        RECT -26.685 -103.525 -26.355 -103.195 ;
        RECT -26.685 -108.965 -26.355 -108.635 ;
        RECT -26.685 -110.325 -26.355 -109.995 ;
        RECT -26.685 -113.045 -26.355 -112.715 ;
        RECT -26.685 -114.405 -26.355 -114.075 ;
        RECT -26.685 -115.765 -26.355 -115.435 ;
        RECT -26.685 -117.125 -26.355 -116.795 ;
        RECT -26.685 -118.485 -26.355 -118.155 ;
        RECT -26.685 -121.205 -26.355 -120.875 ;
        RECT -26.685 -122.565 -26.355 -122.235 ;
        RECT -26.685 -123.925 -26.355 -123.595 ;
        RECT -26.685 -126.645 -26.355 -126.315 ;
        RECT -26.685 -129.365 -26.355 -129.035 ;
        RECT -26.685 -130.725 -26.355 -130.395 ;
        RECT -26.685 -133.445 -26.355 -133.115 ;
        RECT -26.685 -134.805 -26.355 -134.475 ;
        RECT -26.685 -136.165 -26.355 -135.835 ;
        RECT -26.685 -137.525 -26.355 -137.195 ;
        RECT -26.685 -140.245 -26.355 -139.915 ;
        RECT -26.685 -142.965 -26.355 -142.635 ;
        RECT -26.685 -144.325 -26.355 -143.995 ;
        RECT -26.685 -145.685 -26.355 -145.355 ;
        RECT -26.685 -147.045 -26.355 -146.715 ;
        RECT -26.685 -148.405 -26.355 -148.075 ;
        RECT -26.685 -149.765 -26.355 -149.435 ;
        RECT -26.685 -151.125 -26.355 -150.795 ;
        RECT -26.685 -152.485 -26.355 -152.155 ;
        RECT -26.685 -153.845 -26.355 -153.515 ;
        RECT -26.685 -155.205 -26.355 -154.875 ;
        RECT -26.685 -156.565 -26.355 -156.235 ;
        RECT -26.685 -157.925 -26.355 -157.595 ;
        RECT -26.685 -159.285 -26.355 -158.955 ;
        RECT -26.685 -160.645 -26.355 -160.315 ;
        RECT -26.685 -162.005 -26.355 -161.675 ;
        RECT -26.685 -163.365 -26.355 -163.035 ;
        RECT -26.685 -166.085 -26.355 -165.755 ;
        RECT -26.685 -167.445 -26.355 -167.115 ;
        RECT -26.685 -171.525 -26.355 -171.195 ;
        RECT -26.685 -172.885 -26.355 -172.555 ;
        RECT -26.685 -174.245 -26.355 -173.915 ;
        RECT -26.685 -175.605 -26.355 -175.275 ;
        RECT -26.685 -176.965 -26.355 -176.635 ;
        RECT -26.685 -179.685 -26.355 -179.355 ;
        RECT -26.685 -181.045 -26.355 -180.715 ;
        RECT -26.685 -182.405 -26.355 -182.075 ;
        RECT -26.685 -183.765 -26.355 -183.435 ;
        RECT -26.685 -185.125 -26.355 -184.795 ;
        RECT -26.685 -186.485 -26.355 -186.155 ;
        RECT -26.685 -189.205 -26.355 -188.875 ;
        RECT -26.685 -190.565 -26.355 -190.235 ;
        RECT -26.685 -196.005 -26.355 -195.675 ;
        RECT -26.685 -197.365 -26.355 -197.035 ;
        RECT -26.685 -198.725 -26.355 -198.395 ;
        RECT -26.685 -200.085 -26.355 -199.755 ;
        RECT -26.685 -201.445 -26.355 -201.115 ;
        RECT -26.685 -202.805 -26.355 -202.475 ;
        RECT -26.685 -204.165 -26.355 -203.835 ;
        RECT -26.685 -205.525 -26.355 -205.195 ;
        RECT -26.685 -208.245 -26.355 -207.915 ;
        RECT -26.685 -210.965 -26.355 -210.635 ;
        RECT -26.685 -212.325 -26.355 -211.995 ;
        RECT -26.685 -213.625 -26.355 -213.295 ;
        RECT -26.685 -215.045 -26.355 -214.715 ;
        RECT -26.685 -216.405 -26.355 -216.075 ;
        RECT -26.685 -217.765 -26.355 -217.435 ;
        RECT -26.685 -219.125 -26.355 -218.795 ;
        RECT -26.685 -221.37 -26.355 -220.24 ;
        RECT -26.68 -221.485 -26.36 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -25.325 129.8 -24.995 130.93 ;
        RECT -25.325 127.675 -24.995 128.005 ;
        RECT -25.325 126.315 -24.995 126.645 ;
        RECT -25.325 124.955 -24.995 125.285 ;
        RECT -25.325 123.595 -24.995 123.925 ;
        RECT -25.325 122.235 -24.995 122.565 ;
        RECT -25.325 120.875 -24.995 121.205 ;
        RECT -25.325 119.515 -24.995 119.845 ;
        RECT -25.325 118.155 -24.995 118.485 ;
        RECT -25.325 116.795 -24.995 117.125 ;
        RECT -25.325 115.435 -24.995 115.765 ;
        RECT -25.325 114.075 -24.995 114.405 ;
        RECT -25.325 112.715 -24.995 113.045 ;
        RECT -25.325 111.355 -24.995 111.685 ;
        RECT -25.325 109.995 -24.995 110.325 ;
        RECT -25.325 108.635 -24.995 108.965 ;
        RECT -25.325 107.275 -24.995 107.605 ;
        RECT -25.325 105.915 -24.995 106.245 ;
        RECT -25.325 104.555 -24.995 104.885 ;
        RECT -25.325 103.195 -24.995 103.525 ;
        RECT -25.325 101.835 -24.995 102.165 ;
        RECT -25.325 100.475 -24.995 100.805 ;
        RECT -25.325 99.115 -24.995 99.445 ;
        RECT -25.325 97.755 -24.995 98.085 ;
        RECT -25.325 96.395 -24.995 96.725 ;
        RECT -25.325 95.035 -24.995 95.365 ;
        RECT -25.325 93.675 -24.995 94.005 ;
        RECT -25.325 92.315 -24.995 92.645 ;
        RECT -25.325 90.955 -24.995 91.285 ;
        RECT -25.325 89.595 -24.995 89.925 ;
        RECT -25.325 88.235 -24.995 88.565 ;
        RECT -25.325 86.875 -24.995 87.205 ;
        RECT -25.325 85.515 -24.995 85.845 ;
        RECT -25.325 84.155 -24.995 84.485 ;
        RECT -25.325 82.795 -24.995 83.125 ;
        RECT -25.325 81.435 -24.995 81.765 ;
        RECT -25.325 80.075 -24.995 80.405 ;
        RECT -25.325 78.715 -24.995 79.045 ;
        RECT -25.325 77.355 -24.995 77.685 ;
        RECT -25.325 75.995 -24.995 76.325 ;
        RECT -25.325 74.635 -24.995 74.965 ;
        RECT -25.325 73.275 -24.995 73.605 ;
        RECT -25.325 71.915 -24.995 72.245 ;
        RECT -25.325 70.555 -24.995 70.885 ;
        RECT -25.325 69.195 -24.995 69.525 ;
        RECT -25.325 67.835 -24.995 68.165 ;
        RECT -25.325 66.475 -24.995 66.805 ;
        RECT -25.325 65.115 -24.995 65.445 ;
        RECT -25.325 63.755 -24.995 64.085 ;
        RECT -25.325 62.395 -24.995 62.725 ;
        RECT -25.325 61.035 -24.995 61.365 ;
        RECT -25.325 59.675 -24.995 60.005 ;
        RECT -25.325 58.315 -24.995 58.645 ;
        RECT -25.325 56.955 -24.995 57.285 ;
        RECT -25.325 55.595 -24.995 55.925 ;
        RECT -25.325 54.235 -24.995 54.565 ;
        RECT -25.325 52.875 -24.995 53.205 ;
        RECT -25.325 51.515 -24.995 51.845 ;
        RECT -25.325 50.155 -24.995 50.485 ;
        RECT -25.325 48.795 -24.995 49.125 ;
        RECT -25.325 47.435 -24.995 47.765 ;
        RECT -25.325 46.075 -24.995 46.405 ;
        RECT -25.325 44.715 -24.995 45.045 ;
        RECT -25.325 43.355 -24.995 43.685 ;
        RECT -25.325 41.995 -24.995 42.325 ;
        RECT -25.325 40.635 -24.995 40.965 ;
        RECT -25.325 39.275 -24.995 39.605 ;
        RECT -25.325 37.915 -24.995 38.245 ;
        RECT -25.325 36.555 -24.995 36.885 ;
        RECT -25.325 35.195 -24.995 35.525 ;
        RECT -25.325 33.835 -24.995 34.165 ;
        RECT -25.325 32.475 -24.995 32.805 ;
        RECT -25.325 31.115 -24.995 31.445 ;
        RECT -25.325 29.755 -24.995 30.085 ;
        RECT -25.325 28.395 -24.995 28.725 ;
        RECT -25.325 27.035 -24.995 27.365 ;
        RECT -25.325 25.675 -24.995 26.005 ;
        RECT -25.325 24.315 -24.995 24.645 ;
        RECT -25.325 22.955 -24.995 23.285 ;
        RECT -25.325 21.595 -24.995 21.925 ;
        RECT -25.325 20.235 -24.995 20.565 ;
        RECT -25.325 18.875 -24.995 19.205 ;
        RECT -25.325 17.515 -24.995 17.845 ;
        RECT -25.325 16.155 -24.995 16.485 ;
        RECT -25.325 14.795 -24.995 15.125 ;
        RECT -25.325 13.435 -24.995 13.765 ;
        RECT -25.325 12.075 -24.995 12.405 ;
        RECT -25.325 10.715 -24.995 11.045 ;
        RECT -25.325 9.355 -24.995 9.685 ;
        RECT -25.325 7.995 -24.995 8.325 ;
        RECT -25.325 6.635 -24.995 6.965 ;
        RECT -25.325 5.275 -24.995 5.605 ;
        RECT -25.325 3.915 -24.995 4.245 ;
        RECT -25.325 2.555 -24.995 2.885 ;
        RECT -25.325 1.195 -24.995 1.525 ;
        RECT -25.325 -0.165 -24.995 0.165 ;
        RECT -25.325 -1.525 -24.995 -1.195 ;
        RECT -25.325 -8.325 -24.995 -7.995 ;
        RECT -25.325 -9.685 -24.995 -9.355 ;
        RECT -25.325 -11.16 -24.995 -10.83 ;
        RECT -25.325 -12.405 -24.995 -12.075 ;
        RECT -25.325 -15.125 -24.995 -14.795 ;
        RECT -25.325 -16.25 -24.995 -15.92 ;
        RECT -25.325 -21.925 -24.995 -21.595 ;
        RECT -25.325 -27.365 -24.995 -27.035 ;
        RECT -25.325 -30.085 -24.995 -29.755 ;
        RECT -25.325 -32.34 -24.995 -32.01 ;
        RECT -25.325 -37.43 -24.995 -37.1 ;
        RECT -25.325 -43.685 -24.995 -43.355 ;
        RECT -25.325 -45.045 -24.995 -44.715 ;
        RECT -25.325 -46.405 -24.995 -46.075 ;
        RECT -25.325 -47.765 -24.995 -47.435 ;
        RECT -25.325 -49.125 -24.995 -48.795 ;
        RECT -25.325 -50.485 -24.995 -50.155 ;
        RECT -25.325 -51.845 -24.995 -51.515 ;
        RECT -25.325 -53.205 -24.995 -52.875 ;
        RECT -25.325 -54.565 -24.995 -54.235 ;
        RECT -25.325 -55.925 -24.995 -55.595 ;
        RECT -25.325 -57.285 -24.995 -56.955 ;
        RECT -25.325 -58.645 -24.995 -58.315 ;
        RECT -25.325 -60.005 -24.995 -59.675 ;
        RECT -25.325 -61.365 -24.995 -61.035 ;
        RECT -25.325 -62.725 -24.995 -62.395 ;
        RECT -25.325 -64.085 -24.995 -63.755 ;
        RECT -25.325 -65.445 -24.995 -65.115 ;
        RECT -25.325 -66.805 -24.995 -66.475 ;
        RECT -25.325 -68.165 -24.995 -67.835 ;
        RECT -25.325 -69.525 -24.995 -69.195 ;
        RECT -25.325 -70.885 -24.995 -70.555 ;
        RECT -25.325 -72.245 -24.995 -71.915 ;
        RECT -25.325 -73.605 -24.995 -73.275 ;
        RECT -25.325 -74.965 -24.995 -74.635 ;
        RECT -25.325 -76.325 -24.995 -75.995 ;
        RECT -25.325 -77.685 -24.995 -77.355 ;
        RECT -25.325 -79.045 -24.995 -78.715 ;
        RECT -25.325 -80.405 -24.995 -80.075 ;
        RECT -25.325 -81.765 -24.995 -81.435 ;
        RECT -25.325 -83.125 -24.995 -82.795 ;
        RECT -25.325 -84.485 -24.995 -84.155 ;
        RECT -25.325 -85.845 -24.995 -85.515 ;
        RECT -25.325 -87.205 -24.995 -86.875 ;
        RECT -25.325 -88.565 -24.995 -88.235 ;
        RECT -25.325 -89.925 -24.995 -89.595 ;
        RECT -25.325 -91.285 -24.995 -90.955 ;
        RECT -25.325 -92.645 -24.995 -92.315 ;
        RECT -25.325 -94.005 -24.995 -93.675 ;
        RECT -25.325 -95.365 -24.995 -95.035 ;
        RECT -25.325 -96.725 -24.995 -96.395 ;
        RECT -25.325 -98.085 -24.995 -97.755 ;
        RECT -25.325 -99.445 -24.995 -99.115 ;
        RECT -25.325 -100.805 -24.995 -100.475 ;
        RECT -25.325 -102.165 -24.995 -101.835 ;
        RECT -25.325 -103.525 -24.995 -103.195 ;
        RECT -25.325 -108.965 -24.995 -108.635 ;
        RECT -25.325 -110.325 -24.995 -109.995 ;
        RECT -25.325 -111.685 -24.995 -111.355 ;
        RECT -25.325 -113.045 -24.995 -112.715 ;
        RECT -25.325 -114.405 -24.995 -114.075 ;
        RECT -25.325 -115.765 -24.995 -115.435 ;
        RECT -25.325 -117.125 -24.995 -116.795 ;
        RECT -25.325 -118.485 -24.995 -118.155 ;
        RECT -25.325 -119.845 -24.995 -119.515 ;
        RECT -25.325 -121.205 -24.995 -120.875 ;
        RECT -25.325 -122.565 -24.995 -122.235 ;
        RECT -25.325 -123.925 -24.995 -123.595 ;
        RECT -25.325 -125.285 -24.995 -124.955 ;
        RECT -25.325 -126.645 -24.995 -126.315 ;
        RECT -25.325 -128.005 -24.995 -127.675 ;
        RECT -25.325 -129.365 -24.995 -129.035 ;
        RECT -25.325 -130.725 -24.995 -130.395 ;
        RECT -25.325 -132.085 -24.995 -131.755 ;
        RECT -25.325 -133.445 -24.995 -133.115 ;
        RECT -25.325 -134.805 -24.995 -134.475 ;
        RECT -25.325 -136.165 -24.995 -135.835 ;
        RECT -25.325 -137.525 -24.995 -137.195 ;
        RECT -25.325 -140.245 -24.995 -139.915 ;
        RECT -25.325 -142.965 -24.995 -142.635 ;
        RECT -25.325 -144.325 -24.995 -143.995 ;
        RECT -25.325 -145.685 -24.995 -145.355 ;
        RECT -25.325 -147.045 -24.995 -146.715 ;
        RECT -25.325 -148.405 -24.995 -148.075 ;
        RECT -25.325 -149.765 -24.995 -149.435 ;
        RECT -25.325 -151.125 -24.995 -150.795 ;
        RECT -25.325 -152.485 -24.995 -152.155 ;
        RECT -25.325 -153.845 -24.995 -153.515 ;
        RECT -25.325 -155.205 -24.995 -154.875 ;
        RECT -25.325 -156.565 -24.995 -156.235 ;
        RECT -25.325 -157.925 -24.995 -157.595 ;
        RECT -25.325 -159.285 -24.995 -158.955 ;
        RECT -25.325 -160.645 -24.995 -160.315 ;
        RECT -25.325 -162.005 -24.995 -161.675 ;
        RECT -25.325 -163.365 -24.995 -163.035 ;
        RECT -25.325 -166.085 -24.995 -165.755 ;
        RECT -25.325 -167.445 -24.995 -167.115 ;
        RECT -25.325 -172.885 -24.995 -172.555 ;
        RECT -25.325 -174.245 -24.995 -173.915 ;
        RECT -25.325 -175.605 -24.995 -175.275 ;
        RECT -25.325 -176.965 -24.995 -176.635 ;
        RECT -25.325 -179.685 -24.995 -179.355 ;
        RECT -25.325 -181.045 -24.995 -180.715 ;
        RECT -25.325 -182.405 -24.995 -182.075 ;
        RECT -25.325 -185.125 -24.995 -184.795 ;
        RECT -25.325 -186.485 -24.995 -186.155 ;
        RECT -25.325 -189.205 -24.995 -188.875 ;
        RECT -25.325 -190.565 -24.995 -190.235 ;
        RECT -25.325 -196.005 -24.995 -195.675 ;
        RECT -25.325 -197.365 -24.995 -197.035 ;
        RECT -25.325 -198.725 -24.995 -198.395 ;
        RECT -25.325 -200.085 -24.995 -199.755 ;
        RECT -25.325 -201.445 -24.995 -201.115 ;
        RECT -25.325 -202.805 -24.995 -202.475 ;
        RECT -25.325 -204.165 -24.995 -203.835 ;
        RECT -25.325 -205.525 -24.995 -205.195 ;
        RECT -25.325 -208.245 -24.995 -207.915 ;
        RECT -25.325 -210.965 -24.995 -210.635 ;
        RECT -25.325 -212.325 -24.995 -211.995 ;
        RECT -25.325 -213.625 -24.995 -213.295 ;
        RECT -25.325 -215.045 -24.995 -214.715 ;
        RECT -25.325 -216.405 -24.995 -216.075 ;
        RECT -25.325 -217.765 -24.995 -217.435 ;
        RECT -25.325 -219.125 -24.995 -218.795 ;
        RECT -25.325 -221.37 -24.995 -220.24 ;
        RECT -25.32 -221.485 -25 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.965 129.8 -23.635 130.93 ;
        RECT -23.965 127.675 -23.635 128.005 ;
        RECT -23.965 126.315 -23.635 126.645 ;
        RECT -23.965 124.955 -23.635 125.285 ;
        RECT -23.965 123.595 -23.635 123.925 ;
        RECT -23.965 122.235 -23.635 122.565 ;
        RECT -23.965 120.875 -23.635 121.205 ;
        RECT -23.965 119.515 -23.635 119.845 ;
        RECT -23.965 118.155 -23.635 118.485 ;
        RECT -23.965 116.795 -23.635 117.125 ;
        RECT -23.965 115.435 -23.635 115.765 ;
        RECT -23.965 114.075 -23.635 114.405 ;
        RECT -23.965 112.715 -23.635 113.045 ;
        RECT -23.965 111.355 -23.635 111.685 ;
        RECT -23.965 109.995 -23.635 110.325 ;
        RECT -23.965 108.635 -23.635 108.965 ;
        RECT -23.965 107.275 -23.635 107.605 ;
        RECT -23.965 105.915 -23.635 106.245 ;
        RECT -23.965 104.555 -23.635 104.885 ;
        RECT -23.965 103.195 -23.635 103.525 ;
        RECT -23.965 101.835 -23.635 102.165 ;
        RECT -23.965 100.475 -23.635 100.805 ;
        RECT -23.965 99.115 -23.635 99.445 ;
        RECT -23.965 97.755 -23.635 98.085 ;
        RECT -23.965 96.395 -23.635 96.725 ;
        RECT -23.965 95.035 -23.635 95.365 ;
        RECT -23.965 93.675 -23.635 94.005 ;
        RECT -23.965 92.315 -23.635 92.645 ;
        RECT -23.965 90.955 -23.635 91.285 ;
        RECT -23.965 89.595 -23.635 89.925 ;
        RECT -23.965 88.235 -23.635 88.565 ;
        RECT -23.965 86.875 -23.635 87.205 ;
        RECT -23.965 85.515 -23.635 85.845 ;
        RECT -23.965 84.155 -23.635 84.485 ;
        RECT -23.965 82.795 -23.635 83.125 ;
        RECT -23.965 81.435 -23.635 81.765 ;
        RECT -23.965 80.075 -23.635 80.405 ;
        RECT -23.965 78.715 -23.635 79.045 ;
        RECT -23.965 77.355 -23.635 77.685 ;
        RECT -23.965 75.995 -23.635 76.325 ;
        RECT -23.965 74.635 -23.635 74.965 ;
        RECT -23.965 73.275 -23.635 73.605 ;
        RECT -23.965 71.915 -23.635 72.245 ;
        RECT -23.965 70.555 -23.635 70.885 ;
        RECT -23.965 69.195 -23.635 69.525 ;
        RECT -23.965 67.835 -23.635 68.165 ;
        RECT -23.965 66.475 -23.635 66.805 ;
        RECT -23.965 65.115 -23.635 65.445 ;
        RECT -23.965 63.755 -23.635 64.085 ;
        RECT -23.965 62.395 -23.635 62.725 ;
        RECT -23.965 61.035 -23.635 61.365 ;
        RECT -23.965 59.675 -23.635 60.005 ;
        RECT -23.965 58.315 -23.635 58.645 ;
        RECT -23.965 56.955 -23.635 57.285 ;
        RECT -23.965 55.595 -23.635 55.925 ;
        RECT -23.965 54.235 -23.635 54.565 ;
        RECT -23.965 52.875 -23.635 53.205 ;
        RECT -23.965 51.515 -23.635 51.845 ;
        RECT -23.965 50.155 -23.635 50.485 ;
        RECT -23.965 48.795 -23.635 49.125 ;
        RECT -23.965 47.435 -23.635 47.765 ;
        RECT -23.965 46.075 -23.635 46.405 ;
        RECT -23.965 44.715 -23.635 45.045 ;
        RECT -23.965 43.355 -23.635 43.685 ;
        RECT -23.965 41.995 -23.635 42.325 ;
        RECT -23.965 40.635 -23.635 40.965 ;
        RECT -23.965 39.275 -23.635 39.605 ;
        RECT -23.965 37.915 -23.635 38.245 ;
        RECT -23.965 36.555 -23.635 36.885 ;
        RECT -23.965 35.195 -23.635 35.525 ;
        RECT -23.965 33.835 -23.635 34.165 ;
        RECT -23.965 32.475 -23.635 32.805 ;
        RECT -23.965 31.115 -23.635 31.445 ;
        RECT -23.965 29.755 -23.635 30.085 ;
        RECT -23.965 28.395 -23.635 28.725 ;
        RECT -23.965 27.035 -23.635 27.365 ;
        RECT -23.965 25.675 -23.635 26.005 ;
        RECT -23.965 24.315 -23.635 24.645 ;
        RECT -23.965 22.955 -23.635 23.285 ;
        RECT -23.965 21.595 -23.635 21.925 ;
        RECT -23.965 20.235 -23.635 20.565 ;
        RECT -23.965 18.875 -23.635 19.205 ;
        RECT -23.965 17.515 -23.635 17.845 ;
        RECT -23.965 16.155 -23.635 16.485 ;
        RECT -23.965 14.795 -23.635 15.125 ;
        RECT -23.965 13.435 -23.635 13.765 ;
        RECT -23.965 12.075 -23.635 12.405 ;
        RECT -23.965 10.715 -23.635 11.045 ;
        RECT -23.965 9.355 -23.635 9.685 ;
        RECT -23.965 7.995 -23.635 8.325 ;
        RECT -23.965 6.635 -23.635 6.965 ;
        RECT -23.965 5.275 -23.635 5.605 ;
        RECT -23.965 3.915 -23.635 4.245 ;
        RECT -23.965 2.555 -23.635 2.885 ;
        RECT -23.965 1.195 -23.635 1.525 ;
        RECT -23.965 -0.165 -23.635 0.165 ;
        RECT -23.965 -1.525 -23.635 -1.195 ;
        RECT -23.965 -8.325 -23.635 -7.995 ;
        RECT -23.965 -9.685 -23.635 -9.355 ;
        RECT -23.965 -11.16 -23.635 -10.83 ;
        RECT -23.965 -12.405 -23.635 -12.075 ;
        RECT -23.965 -15.125 -23.635 -14.795 ;
        RECT -23.965 -16.25 -23.635 -15.92 ;
        RECT -23.965 -21.925 -23.635 -21.595 ;
        RECT -23.965 -27.365 -23.635 -27.035 ;
        RECT -23.965 -30.085 -23.635 -29.755 ;
        RECT -23.965 -32.34 -23.635 -32.01 ;
        RECT -23.965 -37.43 -23.635 -37.1 ;
        RECT -23.965 -43.685 -23.635 -43.355 ;
        RECT -23.965 -45.045 -23.635 -44.715 ;
        RECT -23.965 -46.405 -23.635 -46.075 ;
        RECT -23.965 -47.765 -23.635 -47.435 ;
        RECT -23.965 -49.125 -23.635 -48.795 ;
        RECT -23.965 -50.485 -23.635 -50.155 ;
        RECT -23.965 -51.845 -23.635 -51.515 ;
        RECT -23.965 -53.205 -23.635 -52.875 ;
        RECT -23.965 -54.565 -23.635 -54.235 ;
        RECT -23.965 -55.925 -23.635 -55.595 ;
        RECT -23.965 -57.285 -23.635 -56.955 ;
        RECT -23.965 -58.645 -23.635 -58.315 ;
        RECT -23.965 -60.005 -23.635 -59.675 ;
        RECT -23.965 -61.365 -23.635 -61.035 ;
        RECT -23.965 -62.725 -23.635 -62.395 ;
        RECT -23.965 -64.085 -23.635 -63.755 ;
        RECT -23.965 -65.445 -23.635 -65.115 ;
        RECT -23.965 -66.805 -23.635 -66.475 ;
        RECT -23.965 -68.165 -23.635 -67.835 ;
        RECT -23.965 -69.525 -23.635 -69.195 ;
        RECT -23.965 -70.885 -23.635 -70.555 ;
        RECT -23.965 -72.245 -23.635 -71.915 ;
        RECT -23.965 -73.605 -23.635 -73.275 ;
        RECT -23.965 -74.965 -23.635 -74.635 ;
        RECT -23.965 -76.325 -23.635 -75.995 ;
        RECT -23.965 -77.685 -23.635 -77.355 ;
        RECT -23.965 -79.045 -23.635 -78.715 ;
        RECT -23.965 -80.405 -23.635 -80.075 ;
        RECT -23.965 -81.765 -23.635 -81.435 ;
        RECT -23.965 -83.125 -23.635 -82.795 ;
        RECT -23.965 -84.485 -23.635 -84.155 ;
        RECT -23.965 -85.845 -23.635 -85.515 ;
        RECT -23.965 -87.205 -23.635 -86.875 ;
        RECT -23.965 -88.565 -23.635 -88.235 ;
        RECT -23.965 -89.925 -23.635 -89.595 ;
        RECT -23.965 -91.285 -23.635 -90.955 ;
        RECT -23.965 -92.645 -23.635 -92.315 ;
        RECT -23.965 -94.005 -23.635 -93.675 ;
        RECT -23.965 -95.365 -23.635 -95.035 ;
        RECT -23.965 -96.725 -23.635 -96.395 ;
        RECT -23.965 -98.085 -23.635 -97.755 ;
        RECT -23.965 -99.445 -23.635 -99.115 ;
        RECT -23.965 -100.805 -23.635 -100.475 ;
        RECT -23.965 -102.165 -23.635 -101.835 ;
        RECT -23.965 -103.525 -23.635 -103.195 ;
        RECT -23.965 -108.965 -23.635 -108.635 ;
        RECT -23.965 -110.325 -23.635 -109.995 ;
        RECT -23.965 -111.685 -23.635 -111.355 ;
        RECT -23.965 -113.045 -23.635 -112.715 ;
        RECT -23.965 -114.405 -23.635 -114.075 ;
        RECT -23.965 -115.765 -23.635 -115.435 ;
        RECT -23.965 -117.125 -23.635 -116.795 ;
        RECT -23.965 -118.485 -23.635 -118.155 ;
        RECT -23.965 -119.845 -23.635 -119.515 ;
        RECT -23.965 -121.205 -23.635 -120.875 ;
        RECT -23.965 -122.565 -23.635 -122.235 ;
        RECT -23.965 -123.925 -23.635 -123.595 ;
        RECT -23.965 -125.285 -23.635 -124.955 ;
        RECT -23.965 -126.645 -23.635 -126.315 ;
        RECT -23.965 -128.005 -23.635 -127.675 ;
        RECT -23.965 -129.365 -23.635 -129.035 ;
        RECT -23.965 -130.725 -23.635 -130.395 ;
        RECT -23.965 -132.085 -23.635 -131.755 ;
        RECT -23.965 -133.445 -23.635 -133.115 ;
        RECT -23.965 -134.805 -23.635 -134.475 ;
        RECT -23.965 -136.165 -23.635 -135.835 ;
        RECT -23.965 -137.525 -23.635 -137.195 ;
        RECT -23.965 -140.245 -23.635 -139.915 ;
        RECT -23.965 -142.965 -23.635 -142.635 ;
        RECT -23.965 -144.325 -23.635 -143.995 ;
        RECT -23.965 -145.685 -23.635 -145.355 ;
        RECT -23.965 -147.045 -23.635 -146.715 ;
        RECT -23.965 -148.405 -23.635 -148.075 ;
        RECT -23.965 -149.765 -23.635 -149.435 ;
        RECT -23.965 -151.125 -23.635 -150.795 ;
        RECT -23.965 -152.485 -23.635 -152.155 ;
        RECT -23.965 -153.845 -23.635 -153.515 ;
        RECT -23.965 -155.205 -23.635 -154.875 ;
        RECT -23.965 -156.565 -23.635 -156.235 ;
        RECT -23.965 -157.925 -23.635 -157.595 ;
        RECT -23.965 -159.285 -23.635 -158.955 ;
        RECT -23.965 -160.645 -23.635 -160.315 ;
        RECT -23.965 -162.005 -23.635 -161.675 ;
        RECT -23.965 -163.365 -23.635 -163.035 ;
        RECT -23.965 -166.085 -23.635 -165.755 ;
        RECT -23.965 -172.885 -23.635 -172.555 ;
        RECT -23.965 -174.245 -23.635 -173.915 ;
        RECT -23.965 -175.605 -23.635 -175.275 ;
        RECT -23.965 -176.965 -23.635 -176.635 ;
        RECT -23.965 -179.685 -23.635 -179.355 ;
        RECT -23.965 -181.045 -23.635 -180.715 ;
        RECT -23.965 -185.125 -23.635 -184.795 ;
        RECT -23.965 -186.485 -23.635 -186.155 ;
        RECT -23.965 -189.205 -23.635 -188.875 ;
        RECT -23.965 -190.565 -23.635 -190.235 ;
        RECT -23.965 -196.005 -23.635 -195.675 ;
        RECT -23.965 -197.365 -23.635 -197.035 ;
        RECT -23.965 -198.725 -23.635 -198.395 ;
        RECT -23.965 -200.085 -23.635 -199.755 ;
        RECT -23.965 -201.445 -23.635 -201.115 ;
        RECT -23.965 -202.805 -23.635 -202.475 ;
        RECT -23.965 -204.165 -23.635 -203.835 ;
        RECT -23.965 -205.525 -23.635 -205.195 ;
        RECT -23.965 -208.245 -23.635 -207.915 ;
        RECT -23.965 -212.325 -23.635 -211.995 ;
        RECT -23.965 -213.625 -23.635 -213.295 ;
        RECT -23.965 -215.045 -23.635 -214.715 ;
        RECT -23.965 -216.405 -23.635 -216.075 ;
        RECT -23.965 -217.765 -23.635 -217.435 ;
        RECT -23.965 -219.125 -23.635 -218.795 ;
        RECT -23.965 -221.37 -23.635 -220.24 ;
        RECT -23.96 -221.485 -23.64 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -22.605 81.435 -22.275 81.765 ;
        RECT -22.605 80.075 -22.275 80.405 ;
        RECT -22.605 78.715 -22.275 79.045 ;
        RECT -22.605 77.355 -22.275 77.685 ;
        RECT -22.605 75.995 -22.275 76.325 ;
        RECT -22.605 74.635 -22.275 74.965 ;
        RECT -22.605 73.275 -22.275 73.605 ;
        RECT -22.605 71.915 -22.275 72.245 ;
        RECT -22.605 70.555 -22.275 70.885 ;
        RECT -22.605 69.195 -22.275 69.525 ;
        RECT -22.605 67.835 -22.275 68.165 ;
        RECT -22.605 66.475 -22.275 66.805 ;
        RECT -22.605 65.115 -22.275 65.445 ;
        RECT -22.605 63.755 -22.275 64.085 ;
        RECT -22.605 62.395 -22.275 62.725 ;
        RECT -22.605 61.035 -22.275 61.365 ;
        RECT -22.605 59.675 -22.275 60.005 ;
        RECT -22.605 58.315 -22.275 58.645 ;
        RECT -22.605 56.955 -22.275 57.285 ;
        RECT -22.605 55.595 -22.275 55.925 ;
        RECT -22.605 54.235 -22.275 54.565 ;
        RECT -22.605 52.875 -22.275 53.205 ;
        RECT -22.605 51.515 -22.275 51.845 ;
        RECT -22.605 50.155 -22.275 50.485 ;
        RECT -22.605 48.795 -22.275 49.125 ;
        RECT -22.605 47.435 -22.275 47.765 ;
        RECT -22.605 46.075 -22.275 46.405 ;
        RECT -22.605 44.715 -22.275 45.045 ;
        RECT -22.605 43.355 -22.275 43.685 ;
        RECT -22.605 41.995 -22.275 42.325 ;
        RECT -22.605 40.635 -22.275 40.965 ;
        RECT -22.605 39.275 -22.275 39.605 ;
        RECT -22.605 37.915 -22.275 38.245 ;
        RECT -22.605 36.555 -22.275 36.885 ;
        RECT -22.605 35.195 -22.275 35.525 ;
        RECT -22.605 33.835 -22.275 34.165 ;
        RECT -22.605 32.475 -22.275 32.805 ;
        RECT -22.605 31.115 -22.275 31.445 ;
        RECT -22.605 29.755 -22.275 30.085 ;
        RECT -22.605 28.395 -22.275 28.725 ;
        RECT -22.605 27.035 -22.275 27.365 ;
        RECT -22.605 25.675 -22.275 26.005 ;
        RECT -22.605 24.315 -22.275 24.645 ;
        RECT -22.605 22.955 -22.275 23.285 ;
        RECT -22.605 21.595 -22.275 21.925 ;
        RECT -22.605 20.235 -22.275 20.565 ;
        RECT -22.605 18.875 -22.275 19.205 ;
        RECT -22.605 17.515 -22.275 17.845 ;
        RECT -22.605 16.155 -22.275 16.485 ;
        RECT -22.605 14.795 -22.275 15.125 ;
        RECT -22.605 13.435 -22.275 13.765 ;
        RECT -22.605 12.075 -22.275 12.405 ;
        RECT -22.605 10.715 -22.275 11.045 ;
        RECT -22.605 9.355 -22.275 9.685 ;
        RECT -22.605 7.995 -22.275 8.325 ;
        RECT -22.605 6.635 -22.275 6.965 ;
        RECT -22.605 5.275 -22.275 5.605 ;
        RECT -22.605 3.915 -22.275 4.245 ;
        RECT -22.605 2.555 -22.275 2.885 ;
        RECT -22.605 1.195 -22.275 1.525 ;
        RECT -22.605 -0.165 -22.275 0.165 ;
        RECT -22.605 -1.525 -22.275 -1.195 ;
        RECT -22.605 -8.325 -22.275 -7.995 ;
        RECT -22.605 -9.685 -22.275 -9.355 ;
        RECT -22.605 -11.16 -22.275 -10.83 ;
        RECT -22.605 -12.405 -22.275 -12.075 ;
        RECT -22.605 -15.125 -22.275 -14.795 ;
        RECT -22.605 -16.25 -22.275 -15.92 ;
        RECT -22.605 -21.925 -22.275 -21.595 ;
        RECT -22.605 -27.365 -22.275 -27.035 ;
        RECT -22.605 -30.085 -22.275 -29.755 ;
        RECT -22.605 -32.34 -22.275 -32.01 ;
        RECT -22.605 -37.43 -22.275 -37.1 ;
        RECT -22.605 -43.685 -22.275 -43.355 ;
        RECT -22.605 -45.045 -22.275 -44.715 ;
        RECT -22.605 -46.405 -22.275 -46.075 ;
        RECT -22.605 -47.765 -22.275 -47.435 ;
        RECT -22.605 -49.125 -22.275 -48.795 ;
        RECT -22.605 -50.485 -22.275 -50.155 ;
        RECT -22.605 -51.845 -22.275 -51.515 ;
        RECT -22.605 -53.205 -22.275 -52.875 ;
        RECT -22.605 -54.565 -22.275 -54.235 ;
        RECT -22.605 -55.925 -22.275 -55.595 ;
        RECT -22.605 -57.285 -22.275 -56.955 ;
        RECT -22.605 -58.645 -22.275 -58.315 ;
        RECT -22.605 -60.005 -22.275 -59.675 ;
        RECT -22.605 -61.365 -22.275 -61.035 ;
        RECT -22.605 -62.725 -22.275 -62.395 ;
        RECT -22.605 -64.085 -22.275 -63.755 ;
        RECT -22.605 -65.445 -22.275 -65.115 ;
        RECT -22.605 -66.805 -22.275 -66.475 ;
        RECT -22.605 -68.165 -22.275 -67.835 ;
        RECT -22.605 -69.525 -22.275 -69.195 ;
        RECT -22.605 -70.885 -22.275 -70.555 ;
        RECT -22.605 -72.245 -22.275 -71.915 ;
        RECT -22.605 -73.605 -22.275 -73.275 ;
        RECT -22.605 -74.965 -22.275 -74.635 ;
        RECT -22.605 -76.325 -22.275 -75.995 ;
        RECT -22.605 -77.685 -22.275 -77.355 ;
        RECT -22.605 -79.045 -22.275 -78.715 ;
        RECT -22.605 -80.405 -22.275 -80.075 ;
        RECT -22.605 -81.765 -22.275 -81.435 ;
        RECT -22.605 -83.125 -22.275 -82.795 ;
        RECT -22.605 -84.485 -22.275 -84.155 ;
        RECT -22.605 -85.845 -22.275 -85.515 ;
        RECT -22.605 -87.205 -22.275 -86.875 ;
        RECT -22.605 -88.565 -22.275 -88.235 ;
        RECT -22.605 -89.925 -22.275 -89.595 ;
        RECT -22.605 -91.285 -22.275 -90.955 ;
        RECT -22.605 -92.645 -22.275 -92.315 ;
        RECT -22.605 -94.005 -22.275 -93.675 ;
        RECT -22.605 -95.365 -22.275 -95.035 ;
        RECT -22.605 -96.725 -22.275 -96.395 ;
        RECT -22.605 -98.085 -22.275 -97.755 ;
        RECT -22.605 -99.445 -22.275 -99.115 ;
        RECT -22.605 -100.805 -22.275 -100.475 ;
        RECT -22.605 -102.165 -22.275 -101.835 ;
        RECT -22.605 -103.525 -22.275 -103.195 ;
        RECT -22.605 -108.965 -22.275 -108.635 ;
        RECT -22.605 -110.325 -22.275 -109.995 ;
        RECT -22.605 -111.685 -22.275 -111.355 ;
        RECT -22.605 -113.045 -22.275 -112.715 ;
        RECT -22.605 -114.405 -22.275 -114.075 ;
        RECT -22.605 -115.765 -22.275 -115.435 ;
        RECT -22.605 -117.125 -22.275 -116.795 ;
        RECT -22.605 -118.485 -22.275 -118.155 ;
        RECT -22.605 -119.845 -22.275 -119.515 ;
        RECT -22.605 -121.205 -22.275 -120.875 ;
        RECT -22.605 -122.565 -22.275 -122.235 ;
        RECT -22.605 -123.925 -22.275 -123.595 ;
        RECT -22.605 -125.285 -22.275 -124.955 ;
        RECT -22.605 -126.645 -22.275 -126.315 ;
        RECT -22.605 -128.005 -22.275 -127.675 ;
        RECT -22.605 -129.365 -22.275 -129.035 ;
        RECT -22.605 -130.725 -22.275 -130.395 ;
        RECT -22.605 -132.085 -22.275 -131.755 ;
        RECT -22.605 -133.445 -22.275 -133.115 ;
        RECT -22.605 -134.805 -22.275 -134.475 ;
        RECT -22.605 -136.165 -22.275 -135.835 ;
        RECT -22.605 -137.525 -22.275 -137.195 ;
        RECT -22.605 -140.245 -22.275 -139.915 ;
        RECT -22.605 -142.965 -22.275 -142.635 ;
        RECT -22.605 -144.325 -22.275 -143.995 ;
        RECT -22.605 -145.685 -22.275 -145.355 ;
        RECT -22.605 -147.045 -22.275 -146.715 ;
        RECT -22.605 -148.405 -22.275 -148.075 ;
        RECT -22.605 -149.765 -22.275 -149.435 ;
        RECT -22.605 -151.125 -22.275 -150.795 ;
        RECT -22.605 -152.485 -22.275 -152.155 ;
        RECT -22.605 -155.205 -22.275 -154.875 ;
        RECT -22.605 -156.565 -22.275 -156.235 ;
        RECT -22.605 -157.925 -22.275 -157.595 ;
        RECT -22.605 -159.285 -22.275 -158.955 ;
        RECT -22.605 -160.645 -22.275 -160.315 ;
        RECT -22.605 -162.005 -22.275 -161.675 ;
        RECT -22.605 -163.365 -22.275 -163.035 ;
        RECT -22.605 -172.885 -22.275 -172.555 ;
        RECT -22.605 -174.245 -22.275 -173.915 ;
        RECT -22.605 -175.605 -22.275 -175.275 ;
        RECT -22.605 -176.965 -22.275 -176.635 ;
        RECT -22.605 -179.685 -22.275 -179.355 ;
        RECT -22.605 -181.045 -22.275 -180.715 ;
        RECT -22.605 -183.765 -22.275 -183.435 ;
        RECT -22.605 -185.125 -22.275 -184.795 ;
        RECT -22.605 -186.485 -22.275 -186.155 ;
        RECT -22.605 -189.205 -22.275 -188.875 ;
        RECT -22.605 -190.565 -22.275 -190.235 ;
        RECT -22.605 -196.005 -22.275 -195.675 ;
        RECT -22.605 -197.365 -22.275 -197.035 ;
        RECT -22.605 -198.725 -22.275 -198.395 ;
        RECT -22.605 -200.085 -22.275 -199.755 ;
        RECT -22.605 -201.445 -22.275 -201.115 ;
        RECT -22.605 -202.805 -22.275 -202.475 ;
        RECT -22.605 -204.165 -22.275 -203.835 ;
        RECT -22.605 -205.525 -22.275 -205.195 ;
        RECT -22.605 -208.245 -22.275 -207.915 ;
        RECT -22.605 -212.325 -22.275 -211.995 ;
        RECT -22.605 -215.045 -22.275 -214.715 ;
        RECT -22.605 -216.405 -22.275 -216.075 ;
        RECT -22.605 -217.765 -22.275 -217.435 ;
        RECT -22.605 -219.125 -22.275 -218.795 ;
        RECT -22.605 -221.37 -22.275 -220.24 ;
        RECT -22.6 -221.485 -22.28 131.045 ;
        RECT -22.605 129.8 -22.275 130.93 ;
        RECT -22.605 127.675 -22.275 128.005 ;
        RECT -22.605 126.315 -22.275 126.645 ;
        RECT -22.605 124.955 -22.275 125.285 ;
        RECT -22.605 123.595 -22.275 123.925 ;
        RECT -22.605 122.235 -22.275 122.565 ;
        RECT -22.605 120.875 -22.275 121.205 ;
        RECT -22.605 119.515 -22.275 119.845 ;
        RECT -22.605 118.155 -22.275 118.485 ;
        RECT -22.605 116.795 -22.275 117.125 ;
        RECT -22.605 115.435 -22.275 115.765 ;
        RECT -22.605 114.075 -22.275 114.405 ;
        RECT -22.605 112.715 -22.275 113.045 ;
        RECT -22.605 111.355 -22.275 111.685 ;
        RECT -22.605 109.995 -22.275 110.325 ;
        RECT -22.605 108.635 -22.275 108.965 ;
        RECT -22.605 107.275 -22.275 107.605 ;
        RECT -22.605 105.915 -22.275 106.245 ;
        RECT -22.605 104.555 -22.275 104.885 ;
        RECT -22.605 103.195 -22.275 103.525 ;
        RECT -22.605 101.835 -22.275 102.165 ;
        RECT -22.605 100.475 -22.275 100.805 ;
        RECT -22.605 99.115 -22.275 99.445 ;
        RECT -22.605 97.755 -22.275 98.085 ;
        RECT -22.605 96.395 -22.275 96.725 ;
        RECT -22.605 95.035 -22.275 95.365 ;
        RECT -22.605 93.675 -22.275 94.005 ;
        RECT -22.605 92.315 -22.275 92.645 ;
        RECT -22.605 90.955 -22.275 91.285 ;
        RECT -22.605 89.595 -22.275 89.925 ;
        RECT -22.605 88.235 -22.275 88.565 ;
        RECT -22.605 86.875 -22.275 87.205 ;
        RECT -22.605 85.515 -22.275 85.845 ;
        RECT -22.605 84.155 -22.275 84.485 ;
        RECT -22.605 82.795 -22.275 83.125 ;
    END
    PORT
      LAYER met3 ;
        RECT -34.845 -212.325 -34.515 -211.995 ;
        RECT -34.845 -215.045 -34.515 -214.715 ;
        RECT -34.845 -216.405 -34.515 -216.075 ;
        RECT -34.845 -217.765 -34.515 -217.435 ;
        RECT -34.845 -219.125 -34.515 -218.795 ;
        RECT -34.845 -221.37 -34.515 -220.24 ;
        RECT -34.84 -221.485 -34.52 -211.995 ;
    END
    PORT
      LAYER met3 ;
        RECT -33.485 129.8 -33.155 130.93 ;
        RECT -33.485 127.675 -33.155 128.005 ;
        RECT -33.485 126.315 -33.155 126.645 ;
        RECT -33.485 124.955 -33.155 125.285 ;
        RECT -33.485 123.595 -33.155 123.925 ;
        RECT -33.485 122.235 -33.155 122.565 ;
        RECT -33.485 120.875 -33.155 121.205 ;
        RECT -33.485 119.515 -33.155 119.845 ;
        RECT -33.485 118.155 -33.155 118.485 ;
        RECT -33.485 116.795 -33.155 117.125 ;
        RECT -33.485 115.435 -33.155 115.765 ;
        RECT -33.485 114.075 -33.155 114.405 ;
        RECT -33.485 112.715 -33.155 113.045 ;
        RECT -33.485 111.355 -33.155 111.685 ;
        RECT -33.485 109.995 -33.155 110.325 ;
        RECT -33.485 108.635 -33.155 108.965 ;
        RECT -33.485 107.275 -33.155 107.605 ;
        RECT -33.485 105.915 -33.155 106.245 ;
        RECT -33.485 104.555 -33.155 104.885 ;
        RECT -33.485 103.195 -33.155 103.525 ;
        RECT -33.485 101.835 -33.155 102.165 ;
        RECT -33.485 100.475 -33.155 100.805 ;
        RECT -33.485 99.115 -33.155 99.445 ;
        RECT -33.485 97.755 -33.155 98.085 ;
        RECT -33.485 96.395 -33.155 96.725 ;
        RECT -33.485 95.035 -33.155 95.365 ;
        RECT -33.485 93.675 -33.155 94.005 ;
        RECT -33.485 92.315 -33.155 92.645 ;
        RECT -33.485 90.955 -33.155 91.285 ;
        RECT -33.485 89.595 -33.155 89.925 ;
        RECT -33.485 88.235 -33.155 88.565 ;
        RECT -33.485 86.875 -33.155 87.205 ;
        RECT -33.485 85.515 -33.155 85.845 ;
        RECT -33.485 84.155 -33.155 84.485 ;
        RECT -33.485 82.795 -33.155 83.125 ;
        RECT -33.485 81.435 -33.155 81.765 ;
        RECT -33.485 80.075 -33.155 80.405 ;
        RECT -33.485 78.715 -33.155 79.045 ;
        RECT -33.485 77.355 -33.155 77.685 ;
        RECT -33.485 75.995 -33.155 76.325 ;
        RECT -33.485 74.635 -33.155 74.965 ;
        RECT -33.485 73.275 -33.155 73.605 ;
        RECT -33.485 71.915 -33.155 72.245 ;
        RECT -33.485 70.555 -33.155 70.885 ;
        RECT -33.485 69.195 -33.155 69.525 ;
        RECT -33.485 67.835 -33.155 68.165 ;
        RECT -33.485 66.475 -33.155 66.805 ;
        RECT -33.485 65.115 -33.155 65.445 ;
        RECT -33.485 63.755 -33.155 64.085 ;
        RECT -33.485 62.395 -33.155 62.725 ;
        RECT -33.485 61.035 -33.155 61.365 ;
        RECT -33.485 59.675 -33.155 60.005 ;
        RECT -33.485 58.315 -33.155 58.645 ;
        RECT -33.485 56.955 -33.155 57.285 ;
        RECT -33.485 55.595 -33.155 55.925 ;
        RECT -33.485 54.235 -33.155 54.565 ;
        RECT -33.485 52.875 -33.155 53.205 ;
        RECT -33.485 51.515 -33.155 51.845 ;
        RECT -33.485 50.155 -33.155 50.485 ;
        RECT -33.485 48.795 -33.155 49.125 ;
        RECT -33.485 47.435 -33.155 47.765 ;
        RECT -33.485 46.075 -33.155 46.405 ;
        RECT -33.485 44.715 -33.155 45.045 ;
        RECT -33.485 43.355 -33.155 43.685 ;
        RECT -33.485 41.995 -33.155 42.325 ;
        RECT -33.485 40.635 -33.155 40.965 ;
        RECT -33.485 39.275 -33.155 39.605 ;
        RECT -33.485 37.915 -33.155 38.245 ;
        RECT -33.485 36.555 -33.155 36.885 ;
        RECT -33.485 35.195 -33.155 35.525 ;
        RECT -33.485 33.835 -33.155 34.165 ;
        RECT -33.485 32.475 -33.155 32.805 ;
        RECT -33.485 31.115 -33.155 31.445 ;
        RECT -33.485 29.755 -33.155 30.085 ;
        RECT -33.485 28.395 -33.155 28.725 ;
        RECT -33.485 27.035 -33.155 27.365 ;
        RECT -33.485 25.675 -33.155 26.005 ;
        RECT -33.485 24.315 -33.155 24.645 ;
        RECT -33.485 22.955 -33.155 23.285 ;
        RECT -33.485 21.595 -33.155 21.925 ;
        RECT -33.485 20.235 -33.155 20.565 ;
        RECT -33.485 18.875 -33.155 19.205 ;
        RECT -33.485 17.515 -33.155 17.845 ;
        RECT -33.485 16.155 -33.155 16.485 ;
        RECT -33.485 14.795 -33.155 15.125 ;
        RECT -33.485 13.435 -33.155 13.765 ;
        RECT -33.485 12.075 -33.155 12.405 ;
        RECT -33.485 10.715 -33.155 11.045 ;
        RECT -33.485 9.355 -33.155 9.685 ;
        RECT -33.485 7.995 -33.155 8.325 ;
        RECT -33.485 6.635 -33.155 6.965 ;
        RECT -33.485 5.275 -33.155 5.605 ;
        RECT -33.485 3.915 -33.155 4.245 ;
        RECT -33.485 2.555 -33.155 2.885 ;
        RECT -33.485 1.195 -33.155 1.525 ;
        RECT -33.485 -0.165 -33.155 0.165 ;
        RECT -33.485 -6.965 -33.155 -6.635 ;
        RECT -33.485 -8.325 -33.155 -7.995 ;
        RECT -33.485 -9.685 -33.155 -9.355 ;
        RECT -33.485 -11.045 -33.155 -10.715 ;
        RECT -33.485 -12.405 -33.155 -12.075 ;
        RECT -33.485 -13.765 -33.155 -13.435 ;
        RECT -33.485 -15.125 -33.155 -14.795 ;
        RECT -33.485 -16.485 -33.155 -16.155 ;
        RECT -33.485 -17.845 -33.155 -17.515 ;
        RECT -33.485 -19.205 -33.155 -18.875 ;
        RECT -33.485 -20.565 -33.155 -20.235 ;
        RECT -33.485 -27.365 -33.155 -27.035 ;
        RECT -33.485 -28.725 -33.155 -28.395 ;
        RECT -33.485 -30.085 -33.155 -29.755 ;
        RECT -33.485 -32.805 -33.155 -32.475 ;
        RECT -33.485 -35.525 -33.155 -35.195 ;
        RECT -33.485 -36.885 -33.155 -36.555 ;
        RECT -33.485 -39.605 -33.155 -39.275 ;
        RECT -33.485 -40.965 -33.155 -40.635 ;
        RECT -33.485 -42.325 -33.155 -41.995 ;
        RECT -33.485 -43.685 -33.155 -43.355 ;
        RECT -33.485 -45.045 -33.155 -44.715 ;
        RECT -33.485 -46.405 -33.155 -46.075 ;
        RECT -33.485 -47.765 -33.155 -47.435 ;
        RECT -33.485 -49.125 -33.155 -48.795 ;
        RECT -33.485 -50.485 -33.155 -50.155 ;
        RECT -33.485 -51.845 -33.155 -51.515 ;
        RECT -33.485 -53.205 -33.155 -52.875 ;
        RECT -33.485 -54.565 -33.155 -54.235 ;
        RECT -33.485 -55.925 -33.155 -55.595 ;
        RECT -33.485 -57.285 -33.155 -56.955 ;
        RECT -33.485 -58.645 -33.155 -58.315 ;
        RECT -33.485 -60.005 -33.155 -59.675 ;
        RECT -33.485 -61.365 -33.155 -61.035 ;
        RECT -33.485 -62.725 -33.155 -62.395 ;
        RECT -33.485 -64.085 -33.155 -63.755 ;
        RECT -33.485 -65.445 -33.155 -65.115 ;
        RECT -33.485 -66.805 -33.155 -66.475 ;
        RECT -33.485 -68.165 -33.155 -67.835 ;
        RECT -33.485 -69.525 -33.155 -69.195 ;
        RECT -33.485 -70.885 -33.155 -70.555 ;
        RECT -33.485 -72.245 -33.155 -71.915 ;
        RECT -33.485 -73.605 -33.155 -73.275 ;
        RECT -33.485 -74.965 -33.155 -74.635 ;
        RECT -33.485 -76.325 -33.155 -75.995 ;
        RECT -33.485 -77.685 -33.155 -77.355 ;
        RECT -33.485 -79.045 -33.155 -78.715 ;
        RECT -33.485 -80.405 -33.155 -80.075 ;
        RECT -33.485 -81.765 -33.155 -81.435 ;
        RECT -33.485 -83.125 -33.155 -82.795 ;
        RECT -33.485 -84.485 -33.155 -84.155 ;
        RECT -33.485 -85.845 -33.155 -85.515 ;
        RECT -33.485 -87.205 -33.155 -86.875 ;
        RECT -33.485 -88.565 -33.155 -88.235 ;
        RECT -33.485 -89.925 -33.155 -89.595 ;
        RECT -33.485 -91.285 -33.155 -90.955 ;
        RECT -33.485 -92.645 -33.155 -92.315 ;
        RECT -33.485 -94.005 -33.155 -93.675 ;
        RECT -33.485 -95.365 -33.155 -95.035 ;
        RECT -33.485 -96.725 -33.155 -96.395 ;
        RECT -33.485 -98.085 -33.155 -97.755 ;
        RECT -33.485 -99.445 -33.155 -99.115 ;
        RECT -33.485 -100.805 -33.155 -100.475 ;
        RECT -33.485 -102.165 -33.155 -101.835 ;
        RECT -33.485 -103.525 -33.155 -103.195 ;
        RECT -33.485 -106.245 -33.155 -105.915 ;
        RECT -33.485 -108.965 -33.155 -108.635 ;
        RECT -33.485 -110.325 -33.155 -109.995 ;
        RECT -33.485 -113.045 -33.155 -112.715 ;
        RECT -33.485 -114.405 -33.155 -114.075 ;
        RECT -33.485 -115.765 -33.155 -115.435 ;
        RECT -33.485 -117.125 -33.155 -116.795 ;
        RECT -33.485 -118.485 -33.155 -118.155 ;
        RECT -33.485 -119.79 -33.155 -119.46 ;
        RECT -33.485 -121.205 -33.155 -120.875 ;
        RECT -33.485 -122.565 -33.155 -122.235 ;
        RECT -33.485 -123.925 -33.155 -123.595 ;
        RECT -33.485 -126.645 -33.155 -126.315 ;
        RECT -33.485 -128.43 -33.155 -128.1 ;
        RECT -33.485 -129.365 -33.155 -129.035 ;
        RECT -33.485 -130.725 -33.155 -130.395 ;
        RECT -33.485 -133.445 -33.155 -133.115 ;
        RECT -33.485 -134.805 -33.155 -134.475 ;
        RECT -33.485 -136.165 -33.155 -135.835 ;
        RECT -33.485 -137.525 -33.155 -137.195 ;
        RECT -33.485 -140.245 -33.155 -139.915 ;
        RECT -33.485 -142.965 -33.155 -142.635 ;
        RECT -33.485 -144.325 -33.155 -143.995 ;
        RECT -33.485 -145.685 -33.155 -145.355 ;
        RECT -33.485 -147.045 -33.155 -146.715 ;
        RECT -33.485 -148.405 -33.155 -148.075 ;
        RECT -33.485 -149.765 -33.155 -149.435 ;
        RECT -33.485 -151.125 -33.155 -150.795 ;
        RECT -33.485 -152.485 -33.155 -152.155 ;
        RECT -33.485 -153.845 -33.155 -153.515 ;
        RECT -33.485 -155.205 -33.155 -154.875 ;
        RECT -33.485 -156.565 -33.155 -156.235 ;
        RECT -33.485 -157.925 -33.155 -157.595 ;
        RECT -33.485 -159.285 -33.155 -158.955 ;
        RECT -33.485 -160.645 -33.155 -160.315 ;
        RECT -33.485 -162.005 -33.155 -161.675 ;
        RECT -33.485 -163.365 -33.155 -163.035 ;
        RECT -33.485 -164.725 -33.155 -164.395 ;
        RECT -33.485 -166.085 -33.155 -165.755 ;
        RECT -33.485 -167.445 -33.155 -167.115 ;
        RECT -33.485 -168.805 -33.155 -168.475 ;
        RECT -33.485 -171.525 -33.155 -171.195 ;
        RECT -33.485 -172.885 -33.155 -172.555 ;
        RECT -33.485 -174.245 -33.155 -173.915 ;
        RECT -33.485 -175.605 -33.155 -175.275 ;
        RECT -33.485 -176.965 -33.155 -176.635 ;
        RECT -33.485 -178.325 -33.155 -177.995 ;
        RECT -33.485 -179.685 -33.155 -179.355 ;
        RECT -33.485 -181.045 -33.155 -180.715 ;
        RECT -33.485 -182.405 -33.155 -182.075 ;
        RECT -33.485 -183.765 -33.155 -183.435 ;
        RECT -33.485 -185.125 -33.155 -184.795 ;
        RECT -33.485 -186.485 -33.155 -186.155 ;
        RECT -33.485 -189.205 -33.155 -188.875 ;
        RECT -33.485 -190.565 -33.155 -190.235 ;
        RECT -33.485 -193.285 -33.155 -192.955 ;
        RECT -33.485 -196.005 -33.155 -195.675 ;
        RECT -33.485 -197.365 -33.155 -197.035 ;
        RECT -33.485 -198.725 -33.155 -198.395 ;
        RECT -33.485 -200.085 -33.155 -199.755 ;
        RECT -33.485 -201.445 -33.155 -201.115 ;
        RECT -33.485 -202.805 -33.155 -202.475 ;
        RECT -33.485 -204.165 -33.155 -203.835 ;
        RECT -33.485 -205.525 -33.155 -205.195 ;
        RECT -33.485 -208.245 -33.155 -207.915 ;
        RECT -33.485 -212.325 -33.155 -211.995 ;
        RECT -33.485 -213.625 -33.155 -213.295 ;
        RECT -33.485 -215.045 -33.155 -214.715 ;
        RECT -33.485 -216.405 -33.155 -216.075 ;
        RECT -33.485 -217.765 -33.155 -217.435 ;
        RECT -33.485 -219.125 -33.155 -218.795 ;
        RECT -33.485 -221.37 -33.155 -220.24 ;
        RECT -33.48 -221.485 -33.16 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -32.125 129.8 -31.795 130.93 ;
        RECT -32.125 127.675 -31.795 128.005 ;
        RECT -32.125 126.315 -31.795 126.645 ;
        RECT -32.125 124.955 -31.795 125.285 ;
        RECT -32.125 123.595 -31.795 123.925 ;
        RECT -32.125 122.235 -31.795 122.565 ;
        RECT -32.125 120.875 -31.795 121.205 ;
        RECT -32.125 119.515 -31.795 119.845 ;
        RECT -32.125 118.155 -31.795 118.485 ;
        RECT -32.125 116.795 -31.795 117.125 ;
        RECT -32.125 115.435 -31.795 115.765 ;
        RECT -32.125 114.075 -31.795 114.405 ;
        RECT -32.125 112.715 -31.795 113.045 ;
        RECT -32.125 111.355 -31.795 111.685 ;
        RECT -32.125 109.995 -31.795 110.325 ;
        RECT -32.125 108.635 -31.795 108.965 ;
        RECT -32.125 107.275 -31.795 107.605 ;
        RECT -32.125 105.915 -31.795 106.245 ;
        RECT -32.125 104.555 -31.795 104.885 ;
        RECT -32.125 103.195 -31.795 103.525 ;
        RECT -32.125 101.835 -31.795 102.165 ;
        RECT -32.125 100.475 -31.795 100.805 ;
        RECT -32.125 99.115 -31.795 99.445 ;
        RECT -32.125 97.755 -31.795 98.085 ;
        RECT -32.125 96.395 -31.795 96.725 ;
        RECT -32.125 95.035 -31.795 95.365 ;
        RECT -32.125 93.675 -31.795 94.005 ;
        RECT -32.125 92.315 -31.795 92.645 ;
        RECT -32.125 90.955 -31.795 91.285 ;
        RECT -32.125 89.595 -31.795 89.925 ;
        RECT -32.125 88.235 -31.795 88.565 ;
        RECT -32.125 86.875 -31.795 87.205 ;
        RECT -32.125 85.515 -31.795 85.845 ;
        RECT -32.125 84.155 -31.795 84.485 ;
        RECT -32.125 82.795 -31.795 83.125 ;
        RECT -32.125 81.435 -31.795 81.765 ;
        RECT -32.125 80.075 -31.795 80.405 ;
        RECT -32.125 78.715 -31.795 79.045 ;
        RECT -32.125 77.355 -31.795 77.685 ;
        RECT -32.125 75.995 -31.795 76.325 ;
        RECT -32.125 74.635 -31.795 74.965 ;
        RECT -32.125 73.275 -31.795 73.605 ;
        RECT -32.125 71.915 -31.795 72.245 ;
        RECT -32.125 70.555 -31.795 70.885 ;
        RECT -32.125 69.195 -31.795 69.525 ;
        RECT -32.125 67.835 -31.795 68.165 ;
        RECT -32.125 66.475 -31.795 66.805 ;
        RECT -32.125 65.115 -31.795 65.445 ;
        RECT -32.125 63.755 -31.795 64.085 ;
        RECT -32.125 62.395 -31.795 62.725 ;
        RECT -32.125 61.035 -31.795 61.365 ;
        RECT -32.125 59.675 -31.795 60.005 ;
        RECT -32.125 58.315 -31.795 58.645 ;
        RECT -32.125 56.955 -31.795 57.285 ;
        RECT -32.125 55.595 -31.795 55.925 ;
        RECT -32.125 54.235 -31.795 54.565 ;
        RECT -32.125 52.875 -31.795 53.205 ;
        RECT -32.125 51.515 -31.795 51.845 ;
        RECT -32.125 50.155 -31.795 50.485 ;
        RECT -32.125 48.795 -31.795 49.125 ;
        RECT -32.125 47.435 -31.795 47.765 ;
        RECT -32.125 46.075 -31.795 46.405 ;
        RECT -32.125 44.715 -31.795 45.045 ;
        RECT -32.125 43.355 -31.795 43.685 ;
        RECT -32.125 41.995 -31.795 42.325 ;
        RECT -32.125 40.635 -31.795 40.965 ;
        RECT -32.125 39.275 -31.795 39.605 ;
        RECT -32.125 37.915 -31.795 38.245 ;
        RECT -32.125 36.555 -31.795 36.885 ;
        RECT -32.125 35.195 -31.795 35.525 ;
        RECT -32.125 33.835 -31.795 34.165 ;
        RECT -32.125 32.475 -31.795 32.805 ;
        RECT -32.125 31.115 -31.795 31.445 ;
        RECT -32.125 29.755 -31.795 30.085 ;
        RECT -32.125 28.395 -31.795 28.725 ;
        RECT -32.125 27.035 -31.795 27.365 ;
        RECT -32.125 25.675 -31.795 26.005 ;
        RECT -32.125 24.315 -31.795 24.645 ;
        RECT -32.125 22.955 -31.795 23.285 ;
        RECT -32.125 21.595 -31.795 21.925 ;
        RECT -32.125 20.235 -31.795 20.565 ;
        RECT -32.125 18.875 -31.795 19.205 ;
        RECT -32.125 17.515 -31.795 17.845 ;
        RECT -32.125 16.155 -31.795 16.485 ;
        RECT -32.125 14.795 -31.795 15.125 ;
        RECT -32.125 13.435 -31.795 13.765 ;
        RECT -32.125 12.075 -31.795 12.405 ;
        RECT -32.125 10.715 -31.795 11.045 ;
        RECT -32.125 9.355 -31.795 9.685 ;
        RECT -32.125 7.995 -31.795 8.325 ;
        RECT -32.125 6.635 -31.795 6.965 ;
        RECT -32.125 5.275 -31.795 5.605 ;
        RECT -32.125 3.915 -31.795 4.245 ;
        RECT -32.125 2.555 -31.795 2.885 ;
        RECT -32.125 1.195 -31.795 1.525 ;
        RECT -32.125 -0.165 -31.795 0.165 ;
        RECT -32.125 -6.965 -31.795 -6.635 ;
        RECT -32.125 -8.325 -31.795 -7.995 ;
        RECT -32.125 -9.685 -31.795 -9.355 ;
        RECT -32.125 -11.045 -31.795 -10.715 ;
        RECT -32.125 -12.405 -31.795 -12.075 ;
        RECT -32.125 -13.765 -31.795 -13.435 ;
        RECT -32.125 -15.125 -31.795 -14.795 ;
        RECT -32.125 -16.485 -31.795 -16.155 ;
        RECT -32.125 -17.845 -31.795 -17.515 ;
        RECT -32.125 -19.205 -31.795 -18.875 ;
        RECT -32.125 -20.565 -31.795 -20.235 ;
        RECT -32.125 -27.365 -31.795 -27.035 ;
        RECT -32.125 -28.725 -31.795 -28.395 ;
        RECT -32.125 -30.085 -31.795 -29.755 ;
        RECT -32.125 -32.805 -31.795 -32.475 ;
        RECT -32.125 -35.525 -31.795 -35.195 ;
        RECT -32.125 -36.885 -31.795 -36.555 ;
        RECT -32.125 -39.605 -31.795 -39.275 ;
        RECT -32.125 -40.965 -31.795 -40.635 ;
        RECT -32.125 -42.325 -31.795 -41.995 ;
        RECT -32.125 -43.685 -31.795 -43.355 ;
        RECT -32.125 -45.045 -31.795 -44.715 ;
        RECT -32.125 -46.405 -31.795 -46.075 ;
        RECT -32.125 -47.765 -31.795 -47.435 ;
        RECT -32.125 -49.125 -31.795 -48.795 ;
        RECT -32.125 -50.485 -31.795 -50.155 ;
        RECT -32.125 -51.845 -31.795 -51.515 ;
        RECT -32.125 -53.205 -31.795 -52.875 ;
        RECT -32.125 -54.565 -31.795 -54.235 ;
        RECT -32.125 -55.925 -31.795 -55.595 ;
        RECT -32.125 -57.285 -31.795 -56.955 ;
        RECT -32.125 -58.645 -31.795 -58.315 ;
        RECT -32.125 -60.005 -31.795 -59.675 ;
        RECT -32.125 -61.365 -31.795 -61.035 ;
        RECT -32.125 -62.725 -31.795 -62.395 ;
        RECT -32.125 -64.085 -31.795 -63.755 ;
        RECT -32.125 -65.445 -31.795 -65.115 ;
        RECT -32.125 -66.805 -31.795 -66.475 ;
        RECT -32.125 -68.165 -31.795 -67.835 ;
        RECT -32.125 -69.525 -31.795 -69.195 ;
        RECT -32.125 -70.885 -31.795 -70.555 ;
        RECT -32.125 -72.245 -31.795 -71.915 ;
        RECT -32.125 -73.605 -31.795 -73.275 ;
        RECT -32.125 -74.965 -31.795 -74.635 ;
        RECT -32.125 -76.325 -31.795 -75.995 ;
        RECT -32.125 -77.685 -31.795 -77.355 ;
        RECT -32.125 -79.045 -31.795 -78.715 ;
        RECT -32.125 -80.405 -31.795 -80.075 ;
        RECT -32.125 -81.765 -31.795 -81.435 ;
        RECT -32.125 -83.125 -31.795 -82.795 ;
        RECT -32.125 -84.485 -31.795 -84.155 ;
        RECT -32.125 -85.845 -31.795 -85.515 ;
        RECT -32.125 -87.205 -31.795 -86.875 ;
        RECT -32.125 -88.565 -31.795 -88.235 ;
        RECT -32.125 -89.925 -31.795 -89.595 ;
        RECT -32.125 -91.285 -31.795 -90.955 ;
        RECT -32.125 -92.645 -31.795 -92.315 ;
        RECT -32.125 -94.005 -31.795 -93.675 ;
        RECT -32.125 -95.365 -31.795 -95.035 ;
        RECT -32.125 -96.725 -31.795 -96.395 ;
        RECT -32.125 -98.085 -31.795 -97.755 ;
        RECT -32.125 -99.445 -31.795 -99.115 ;
        RECT -32.125 -100.805 -31.795 -100.475 ;
        RECT -32.125 -102.165 -31.795 -101.835 ;
        RECT -32.125 -103.525 -31.795 -103.195 ;
        RECT -32.125 -106.245 -31.795 -105.915 ;
        RECT -32.125 -108.965 -31.795 -108.635 ;
        RECT -32.125 -110.325 -31.795 -109.995 ;
        RECT -32.125 -113.045 -31.795 -112.715 ;
        RECT -32.125 -114.405 -31.795 -114.075 ;
        RECT -32.125 -115.765 -31.795 -115.435 ;
        RECT -32.125 -117.125 -31.795 -116.795 ;
        RECT -32.125 -118.485 -31.795 -118.155 ;
        RECT -32.125 -119.79 -31.795 -119.46 ;
        RECT -32.125 -121.205 -31.795 -120.875 ;
        RECT -32.125 -122.565 -31.795 -122.235 ;
        RECT -32.125 -123.925 -31.795 -123.595 ;
        RECT -32.125 -126.645 -31.795 -126.315 ;
        RECT -32.125 -128.43 -31.795 -128.1 ;
        RECT -32.125 -129.365 -31.795 -129.035 ;
        RECT -32.125 -130.725 -31.795 -130.395 ;
        RECT -32.125 -133.445 -31.795 -133.115 ;
        RECT -32.125 -134.805 -31.795 -134.475 ;
        RECT -32.125 -136.165 -31.795 -135.835 ;
        RECT -32.125 -137.525 -31.795 -137.195 ;
        RECT -32.125 -140.245 -31.795 -139.915 ;
        RECT -32.125 -142.965 -31.795 -142.635 ;
        RECT -32.125 -144.325 -31.795 -143.995 ;
        RECT -32.125 -145.685 -31.795 -145.355 ;
        RECT -32.125 -147.045 -31.795 -146.715 ;
        RECT -32.125 -148.405 -31.795 -148.075 ;
        RECT -32.125 -149.765 -31.795 -149.435 ;
        RECT -32.125 -151.125 -31.795 -150.795 ;
        RECT -32.125 -152.485 -31.795 -152.155 ;
        RECT -32.125 -153.845 -31.795 -153.515 ;
        RECT -32.125 -155.205 -31.795 -154.875 ;
        RECT -32.125 -156.565 -31.795 -156.235 ;
        RECT -32.125 -157.925 -31.795 -157.595 ;
        RECT -32.125 -159.285 -31.795 -158.955 ;
        RECT -32.125 -160.645 -31.795 -160.315 ;
        RECT -32.125 -162.005 -31.795 -161.675 ;
        RECT -32.125 -163.365 -31.795 -163.035 ;
        RECT -32.125 -164.725 -31.795 -164.395 ;
        RECT -32.125 -166.085 -31.795 -165.755 ;
        RECT -32.125 -167.445 -31.795 -167.115 ;
        RECT -32.125 -171.525 -31.795 -171.195 ;
        RECT -32.125 -172.885 -31.795 -172.555 ;
        RECT -32.125 -174.245 -31.795 -173.915 ;
        RECT -32.125 -175.605 -31.795 -175.275 ;
        RECT -32.125 -176.965 -31.795 -176.635 ;
        RECT -32.125 -178.325 -31.795 -177.995 ;
        RECT -32.125 -179.685 -31.795 -179.355 ;
        RECT -32.125 -181.045 -31.795 -180.715 ;
        RECT -32.125 -182.405 -31.795 -182.075 ;
        RECT -32.125 -183.765 -31.795 -183.435 ;
        RECT -32.125 -185.125 -31.795 -184.795 ;
        RECT -32.125 -186.485 -31.795 -186.155 ;
        RECT -32.125 -189.205 -31.795 -188.875 ;
        RECT -32.125 -190.565 -31.795 -190.235 ;
        RECT -32.125 -194.645 -31.795 -194.315 ;
        RECT -32.125 -196.005 -31.795 -195.675 ;
        RECT -32.125 -197.365 -31.795 -197.035 ;
        RECT -32.125 -198.725 -31.795 -198.395 ;
        RECT -32.125 -200.085 -31.795 -199.755 ;
        RECT -32.125 -201.445 -31.795 -201.115 ;
        RECT -32.125 -202.805 -31.795 -202.475 ;
        RECT -32.125 -204.165 -31.795 -203.835 ;
        RECT -32.125 -205.525 -31.795 -205.195 ;
        RECT -32.125 -208.245 -31.795 -207.915 ;
        RECT -32.125 -210.965 -31.795 -210.635 ;
        RECT -32.125 -212.325 -31.795 -211.995 ;
        RECT -32.125 -213.625 -31.795 -213.295 ;
        RECT -32.125 -215.045 -31.795 -214.715 ;
        RECT -32.125 -216.405 -31.795 -216.075 ;
        RECT -32.125 -217.765 -31.795 -217.435 ;
        RECT -32.125 -219.125 -31.795 -218.795 ;
        RECT -32.125 -221.37 -31.795 -220.24 ;
        RECT -32.12 -221.485 -31.8 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.765 129.8 -30.435 130.93 ;
        RECT -30.765 127.675 -30.435 128.005 ;
        RECT -30.765 126.315 -30.435 126.645 ;
        RECT -30.765 124.955 -30.435 125.285 ;
        RECT -30.765 123.595 -30.435 123.925 ;
        RECT -30.765 122.235 -30.435 122.565 ;
        RECT -30.765 120.875 -30.435 121.205 ;
        RECT -30.765 119.515 -30.435 119.845 ;
        RECT -30.765 118.155 -30.435 118.485 ;
        RECT -30.765 116.795 -30.435 117.125 ;
        RECT -30.765 115.435 -30.435 115.765 ;
        RECT -30.765 114.075 -30.435 114.405 ;
        RECT -30.765 112.715 -30.435 113.045 ;
        RECT -30.765 111.355 -30.435 111.685 ;
        RECT -30.765 109.995 -30.435 110.325 ;
        RECT -30.765 108.635 -30.435 108.965 ;
        RECT -30.765 107.275 -30.435 107.605 ;
        RECT -30.765 105.915 -30.435 106.245 ;
        RECT -30.765 104.555 -30.435 104.885 ;
        RECT -30.765 103.195 -30.435 103.525 ;
        RECT -30.765 101.835 -30.435 102.165 ;
        RECT -30.765 100.475 -30.435 100.805 ;
        RECT -30.765 99.115 -30.435 99.445 ;
        RECT -30.765 97.755 -30.435 98.085 ;
        RECT -30.765 96.395 -30.435 96.725 ;
        RECT -30.765 95.035 -30.435 95.365 ;
        RECT -30.765 93.675 -30.435 94.005 ;
        RECT -30.765 92.315 -30.435 92.645 ;
        RECT -30.765 90.955 -30.435 91.285 ;
        RECT -30.765 89.595 -30.435 89.925 ;
        RECT -30.765 88.235 -30.435 88.565 ;
        RECT -30.765 86.875 -30.435 87.205 ;
        RECT -30.765 85.515 -30.435 85.845 ;
        RECT -30.765 84.155 -30.435 84.485 ;
        RECT -30.765 82.795 -30.435 83.125 ;
        RECT -30.765 81.435 -30.435 81.765 ;
        RECT -30.765 80.075 -30.435 80.405 ;
        RECT -30.765 78.715 -30.435 79.045 ;
        RECT -30.765 77.355 -30.435 77.685 ;
        RECT -30.765 75.995 -30.435 76.325 ;
        RECT -30.765 74.635 -30.435 74.965 ;
        RECT -30.765 73.275 -30.435 73.605 ;
        RECT -30.765 71.915 -30.435 72.245 ;
        RECT -30.765 70.555 -30.435 70.885 ;
        RECT -30.765 69.195 -30.435 69.525 ;
        RECT -30.765 67.835 -30.435 68.165 ;
        RECT -30.765 66.475 -30.435 66.805 ;
        RECT -30.765 65.115 -30.435 65.445 ;
        RECT -30.765 63.755 -30.435 64.085 ;
        RECT -30.765 62.395 -30.435 62.725 ;
        RECT -30.765 61.035 -30.435 61.365 ;
        RECT -30.765 59.675 -30.435 60.005 ;
        RECT -30.765 58.315 -30.435 58.645 ;
        RECT -30.765 56.955 -30.435 57.285 ;
        RECT -30.765 55.595 -30.435 55.925 ;
        RECT -30.765 54.235 -30.435 54.565 ;
        RECT -30.765 52.875 -30.435 53.205 ;
        RECT -30.765 51.515 -30.435 51.845 ;
        RECT -30.765 50.155 -30.435 50.485 ;
        RECT -30.765 48.795 -30.435 49.125 ;
        RECT -30.765 47.435 -30.435 47.765 ;
        RECT -30.765 46.075 -30.435 46.405 ;
        RECT -30.765 44.715 -30.435 45.045 ;
        RECT -30.765 43.355 -30.435 43.685 ;
        RECT -30.765 41.995 -30.435 42.325 ;
        RECT -30.765 40.635 -30.435 40.965 ;
        RECT -30.765 39.275 -30.435 39.605 ;
        RECT -30.765 37.915 -30.435 38.245 ;
        RECT -30.765 36.555 -30.435 36.885 ;
        RECT -30.765 35.195 -30.435 35.525 ;
        RECT -30.765 33.835 -30.435 34.165 ;
        RECT -30.765 32.475 -30.435 32.805 ;
        RECT -30.765 31.115 -30.435 31.445 ;
        RECT -30.765 29.755 -30.435 30.085 ;
        RECT -30.765 28.395 -30.435 28.725 ;
        RECT -30.765 27.035 -30.435 27.365 ;
        RECT -30.765 25.675 -30.435 26.005 ;
        RECT -30.765 24.315 -30.435 24.645 ;
        RECT -30.765 22.955 -30.435 23.285 ;
        RECT -30.765 21.595 -30.435 21.925 ;
        RECT -30.765 20.235 -30.435 20.565 ;
        RECT -30.765 18.875 -30.435 19.205 ;
        RECT -30.765 17.515 -30.435 17.845 ;
        RECT -30.765 16.155 -30.435 16.485 ;
        RECT -30.765 14.795 -30.435 15.125 ;
        RECT -30.765 13.435 -30.435 13.765 ;
        RECT -30.765 12.075 -30.435 12.405 ;
        RECT -30.765 10.715 -30.435 11.045 ;
        RECT -30.765 9.355 -30.435 9.685 ;
        RECT -30.765 7.995 -30.435 8.325 ;
        RECT -30.765 6.635 -30.435 6.965 ;
        RECT -30.765 5.275 -30.435 5.605 ;
        RECT -30.765 3.915 -30.435 4.245 ;
        RECT -30.765 2.555 -30.435 2.885 ;
        RECT -30.765 1.195 -30.435 1.525 ;
        RECT -30.765 -0.165 -30.435 0.165 ;
        RECT -30.765 -6.965 -30.435 -6.635 ;
        RECT -30.765 -8.325 -30.435 -7.995 ;
        RECT -30.765 -9.685 -30.435 -9.355 ;
        RECT -30.765 -11.045 -30.435 -10.715 ;
        RECT -30.765 -12.405 -30.435 -12.075 ;
        RECT -30.765 -13.765 -30.435 -13.435 ;
        RECT -30.765 -15.125 -30.435 -14.795 ;
        RECT -30.765 -16.485 -30.435 -16.155 ;
        RECT -30.765 -17.845 -30.435 -17.515 ;
        RECT -30.765 -19.205 -30.435 -18.875 ;
        RECT -30.765 -20.565 -30.435 -20.235 ;
        RECT -30.765 -27.365 -30.435 -27.035 ;
        RECT -30.765 -28.725 -30.435 -28.395 ;
        RECT -30.765 -30.085 -30.435 -29.755 ;
        RECT -30.765 -32.805 -30.435 -32.475 ;
        RECT -30.765 -35.525 -30.435 -35.195 ;
        RECT -30.765 -36.885 -30.435 -36.555 ;
        RECT -30.765 -39.605 -30.435 -39.275 ;
        RECT -30.765 -40.965 -30.435 -40.635 ;
        RECT -30.765 -42.325 -30.435 -41.995 ;
        RECT -30.765 -43.685 -30.435 -43.355 ;
        RECT -30.765 -45.045 -30.435 -44.715 ;
        RECT -30.765 -46.405 -30.435 -46.075 ;
        RECT -30.765 -47.765 -30.435 -47.435 ;
        RECT -30.765 -49.125 -30.435 -48.795 ;
        RECT -30.765 -50.485 -30.435 -50.155 ;
        RECT -30.765 -51.845 -30.435 -51.515 ;
        RECT -30.765 -53.205 -30.435 -52.875 ;
        RECT -30.765 -54.565 -30.435 -54.235 ;
        RECT -30.765 -55.925 -30.435 -55.595 ;
        RECT -30.765 -57.285 -30.435 -56.955 ;
        RECT -30.765 -58.645 -30.435 -58.315 ;
        RECT -30.765 -60.005 -30.435 -59.675 ;
        RECT -30.765 -61.365 -30.435 -61.035 ;
        RECT -30.765 -62.725 -30.435 -62.395 ;
        RECT -30.765 -64.085 -30.435 -63.755 ;
        RECT -30.765 -65.445 -30.435 -65.115 ;
        RECT -30.765 -66.805 -30.435 -66.475 ;
        RECT -30.765 -68.165 -30.435 -67.835 ;
        RECT -30.765 -69.525 -30.435 -69.195 ;
        RECT -30.765 -70.885 -30.435 -70.555 ;
        RECT -30.765 -72.245 -30.435 -71.915 ;
        RECT -30.765 -73.605 -30.435 -73.275 ;
        RECT -30.765 -74.965 -30.435 -74.635 ;
        RECT -30.765 -76.325 -30.435 -75.995 ;
        RECT -30.765 -77.685 -30.435 -77.355 ;
        RECT -30.765 -79.045 -30.435 -78.715 ;
        RECT -30.765 -80.405 -30.435 -80.075 ;
        RECT -30.765 -81.765 -30.435 -81.435 ;
        RECT -30.765 -83.125 -30.435 -82.795 ;
        RECT -30.765 -84.485 -30.435 -84.155 ;
        RECT -30.765 -85.845 -30.435 -85.515 ;
        RECT -30.765 -87.205 -30.435 -86.875 ;
        RECT -30.765 -88.565 -30.435 -88.235 ;
        RECT -30.765 -89.925 -30.435 -89.595 ;
        RECT -30.765 -91.285 -30.435 -90.955 ;
        RECT -30.765 -92.645 -30.435 -92.315 ;
        RECT -30.765 -94.005 -30.435 -93.675 ;
        RECT -30.765 -95.365 -30.435 -95.035 ;
        RECT -30.765 -96.725 -30.435 -96.395 ;
        RECT -30.765 -98.085 -30.435 -97.755 ;
        RECT -30.765 -99.445 -30.435 -99.115 ;
        RECT -30.765 -100.805 -30.435 -100.475 ;
        RECT -30.765 -102.165 -30.435 -101.835 ;
        RECT -30.765 -103.525 -30.435 -103.195 ;
        RECT -30.765 -106.245 -30.435 -105.915 ;
        RECT -30.765 -108.965 -30.435 -108.635 ;
        RECT -30.765 -110.325 -30.435 -109.995 ;
        RECT -30.765 -113.045 -30.435 -112.715 ;
        RECT -30.765 -114.405 -30.435 -114.075 ;
        RECT -30.765 -115.765 -30.435 -115.435 ;
        RECT -30.765 -117.125 -30.435 -116.795 ;
        RECT -30.765 -118.485 -30.435 -118.155 ;
        RECT -30.765 -119.79 -30.435 -119.46 ;
        RECT -30.765 -121.205 -30.435 -120.875 ;
        RECT -30.765 -122.565 -30.435 -122.235 ;
        RECT -30.765 -123.925 -30.435 -123.595 ;
        RECT -30.765 -126.645 -30.435 -126.315 ;
        RECT -30.765 -128.43 -30.435 -128.1 ;
        RECT -30.765 -129.365 -30.435 -129.035 ;
        RECT -30.765 -130.725 -30.435 -130.395 ;
        RECT -30.765 -133.445 -30.435 -133.115 ;
        RECT -30.765 -134.805 -30.435 -134.475 ;
        RECT -30.765 -136.165 -30.435 -135.835 ;
        RECT -30.765 -137.525 -30.435 -137.195 ;
        RECT -30.765 -140.245 -30.435 -139.915 ;
        RECT -30.765 -142.965 -30.435 -142.635 ;
        RECT -30.765 -144.325 -30.435 -143.995 ;
        RECT -30.765 -145.685 -30.435 -145.355 ;
        RECT -30.765 -147.045 -30.435 -146.715 ;
        RECT -30.765 -148.405 -30.435 -148.075 ;
        RECT -30.765 -149.765 -30.435 -149.435 ;
        RECT -30.765 -151.125 -30.435 -150.795 ;
        RECT -30.765 -152.485 -30.435 -152.155 ;
        RECT -30.765 -153.845 -30.435 -153.515 ;
        RECT -30.765 -155.205 -30.435 -154.875 ;
        RECT -30.765 -156.565 -30.435 -156.235 ;
        RECT -30.765 -157.925 -30.435 -157.595 ;
        RECT -30.765 -159.285 -30.435 -158.955 ;
        RECT -30.765 -160.645 -30.435 -160.315 ;
        RECT -30.765 -162.005 -30.435 -161.675 ;
        RECT -30.765 -163.365 -30.435 -163.035 ;
        RECT -30.765 -164.725 -30.435 -164.395 ;
        RECT -30.765 -166.085 -30.435 -165.755 ;
        RECT -30.765 -167.445 -30.435 -167.115 ;
        RECT -30.765 -171.525 -30.435 -171.195 ;
        RECT -30.765 -172.885 -30.435 -172.555 ;
        RECT -30.765 -174.245 -30.435 -173.915 ;
        RECT -30.765 -175.605 -30.435 -175.275 ;
        RECT -30.765 -176.965 -30.435 -176.635 ;
        RECT -30.765 -178.325 -30.435 -177.995 ;
        RECT -30.765 -179.685 -30.435 -179.355 ;
        RECT -30.765 -181.045 -30.435 -180.715 ;
        RECT -30.765 -182.405 -30.435 -182.075 ;
        RECT -30.765 -183.765 -30.435 -183.435 ;
        RECT -30.765 -185.125 -30.435 -184.795 ;
        RECT -30.765 -186.485 -30.435 -186.155 ;
        RECT -30.765 -189.205 -30.435 -188.875 ;
        RECT -30.765 -190.565 -30.435 -190.235 ;
        RECT -30.765 -194.645 -30.435 -194.315 ;
        RECT -30.765 -196.005 -30.435 -195.675 ;
        RECT -30.765 -197.365 -30.435 -197.035 ;
        RECT -30.765 -198.725 -30.435 -198.395 ;
        RECT -30.765 -200.085 -30.435 -199.755 ;
        RECT -30.765 -201.445 -30.435 -201.115 ;
        RECT -30.765 -202.805 -30.435 -202.475 ;
        RECT -30.765 -204.165 -30.435 -203.835 ;
        RECT -30.765 -205.525 -30.435 -205.195 ;
        RECT -30.765 -208.245 -30.435 -207.915 ;
        RECT -30.765 -210.965 -30.435 -210.635 ;
        RECT -30.765 -212.325 -30.435 -211.995 ;
        RECT -30.765 -213.625 -30.435 -213.295 ;
        RECT -30.765 -215.045 -30.435 -214.715 ;
        RECT -30.765 -216.405 -30.435 -216.075 ;
        RECT -30.765 -217.765 -30.435 -217.435 ;
        RECT -30.765 -219.125 -30.435 -218.795 ;
        RECT -30.765 -221.37 -30.435 -220.24 ;
        RECT -30.76 -221.485 -30.44 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.405 129.8 -29.075 130.93 ;
        RECT -29.405 127.675 -29.075 128.005 ;
        RECT -29.405 126.315 -29.075 126.645 ;
        RECT -29.405 124.955 -29.075 125.285 ;
        RECT -29.405 123.595 -29.075 123.925 ;
        RECT -29.405 122.235 -29.075 122.565 ;
        RECT -29.405 120.875 -29.075 121.205 ;
        RECT -29.405 119.515 -29.075 119.845 ;
        RECT -29.405 118.155 -29.075 118.485 ;
        RECT -29.405 116.795 -29.075 117.125 ;
        RECT -29.405 115.435 -29.075 115.765 ;
        RECT -29.405 114.075 -29.075 114.405 ;
        RECT -29.405 112.715 -29.075 113.045 ;
        RECT -29.405 111.355 -29.075 111.685 ;
        RECT -29.405 109.995 -29.075 110.325 ;
        RECT -29.405 108.635 -29.075 108.965 ;
        RECT -29.405 107.275 -29.075 107.605 ;
        RECT -29.405 105.915 -29.075 106.245 ;
        RECT -29.405 104.555 -29.075 104.885 ;
        RECT -29.405 103.195 -29.075 103.525 ;
        RECT -29.405 101.835 -29.075 102.165 ;
        RECT -29.405 100.475 -29.075 100.805 ;
        RECT -29.405 99.115 -29.075 99.445 ;
        RECT -29.405 97.755 -29.075 98.085 ;
        RECT -29.405 96.395 -29.075 96.725 ;
        RECT -29.405 95.035 -29.075 95.365 ;
        RECT -29.405 93.675 -29.075 94.005 ;
        RECT -29.405 92.315 -29.075 92.645 ;
        RECT -29.405 90.955 -29.075 91.285 ;
        RECT -29.405 89.595 -29.075 89.925 ;
        RECT -29.405 88.235 -29.075 88.565 ;
        RECT -29.405 86.875 -29.075 87.205 ;
        RECT -29.405 85.515 -29.075 85.845 ;
        RECT -29.405 84.155 -29.075 84.485 ;
        RECT -29.405 82.795 -29.075 83.125 ;
        RECT -29.405 81.435 -29.075 81.765 ;
        RECT -29.405 80.075 -29.075 80.405 ;
        RECT -29.405 78.715 -29.075 79.045 ;
        RECT -29.405 77.355 -29.075 77.685 ;
        RECT -29.405 75.995 -29.075 76.325 ;
        RECT -29.405 74.635 -29.075 74.965 ;
        RECT -29.405 73.275 -29.075 73.605 ;
        RECT -29.405 71.915 -29.075 72.245 ;
        RECT -29.405 70.555 -29.075 70.885 ;
        RECT -29.405 69.195 -29.075 69.525 ;
        RECT -29.405 67.835 -29.075 68.165 ;
        RECT -29.405 66.475 -29.075 66.805 ;
        RECT -29.405 65.115 -29.075 65.445 ;
        RECT -29.405 63.755 -29.075 64.085 ;
        RECT -29.405 62.395 -29.075 62.725 ;
        RECT -29.405 61.035 -29.075 61.365 ;
        RECT -29.405 59.675 -29.075 60.005 ;
        RECT -29.405 58.315 -29.075 58.645 ;
        RECT -29.405 56.955 -29.075 57.285 ;
        RECT -29.405 55.595 -29.075 55.925 ;
        RECT -29.405 54.235 -29.075 54.565 ;
        RECT -29.405 52.875 -29.075 53.205 ;
        RECT -29.405 51.515 -29.075 51.845 ;
        RECT -29.405 50.155 -29.075 50.485 ;
        RECT -29.405 48.795 -29.075 49.125 ;
        RECT -29.405 47.435 -29.075 47.765 ;
        RECT -29.405 46.075 -29.075 46.405 ;
        RECT -29.405 44.715 -29.075 45.045 ;
        RECT -29.405 43.355 -29.075 43.685 ;
        RECT -29.405 41.995 -29.075 42.325 ;
        RECT -29.405 40.635 -29.075 40.965 ;
        RECT -29.405 39.275 -29.075 39.605 ;
        RECT -29.405 37.915 -29.075 38.245 ;
        RECT -29.405 36.555 -29.075 36.885 ;
        RECT -29.405 35.195 -29.075 35.525 ;
        RECT -29.405 33.835 -29.075 34.165 ;
        RECT -29.405 32.475 -29.075 32.805 ;
        RECT -29.405 31.115 -29.075 31.445 ;
        RECT -29.405 29.755 -29.075 30.085 ;
        RECT -29.405 28.395 -29.075 28.725 ;
        RECT -29.405 27.035 -29.075 27.365 ;
        RECT -29.405 25.675 -29.075 26.005 ;
        RECT -29.405 24.315 -29.075 24.645 ;
        RECT -29.405 22.955 -29.075 23.285 ;
        RECT -29.405 21.595 -29.075 21.925 ;
        RECT -29.405 20.235 -29.075 20.565 ;
        RECT -29.405 18.875 -29.075 19.205 ;
        RECT -29.405 17.515 -29.075 17.845 ;
        RECT -29.405 16.155 -29.075 16.485 ;
        RECT -29.405 14.795 -29.075 15.125 ;
        RECT -29.405 13.435 -29.075 13.765 ;
        RECT -29.405 12.075 -29.075 12.405 ;
        RECT -29.405 10.715 -29.075 11.045 ;
        RECT -29.405 9.355 -29.075 9.685 ;
        RECT -29.405 7.995 -29.075 8.325 ;
        RECT -29.405 6.635 -29.075 6.965 ;
        RECT -29.405 5.275 -29.075 5.605 ;
        RECT -29.405 3.915 -29.075 4.245 ;
        RECT -29.405 2.555 -29.075 2.885 ;
        RECT -29.405 1.195 -29.075 1.525 ;
        RECT -29.405 -0.165 -29.075 0.165 ;
        RECT -29.405 -8.325 -29.075 -7.995 ;
        RECT -29.405 -9.685 -29.075 -9.355 ;
        RECT -29.405 -11.16 -29.075 -10.83 ;
        RECT -29.405 -12.405 -29.075 -12.075 ;
        RECT -29.405 -15.125 -29.075 -14.795 ;
        RECT -29.405 -16.25 -29.075 -15.92 ;
        RECT -29.405 -27.365 -29.075 -27.035 ;
        RECT -29.405 -30.085 -29.075 -29.755 ;
        RECT -29.405 -32.34 -29.075 -32.01 ;
        RECT -29.405 -37.43 -29.075 -37.1 ;
        RECT -29.405 -43.685 -29.075 -43.355 ;
        RECT -29.405 -45.045 -29.075 -44.715 ;
        RECT -29.405 -46.405 -29.075 -46.075 ;
        RECT -29.405 -47.765 -29.075 -47.435 ;
        RECT -29.405 -49.125 -29.075 -48.795 ;
        RECT -29.405 -50.485 -29.075 -50.155 ;
        RECT -29.405 -51.845 -29.075 -51.515 ;
        RECT -29.405 -53.205 -29.075 -52.875 ;
        RECT -29.405 -54.565 -29.075 -54.235 ;
        RECT -29.405 -55.925 -29.075 -55.595 ;
        RECT -29.405 -57.285 -29.075 -56.955 ;
        RECT -29.405 -58.645 -29.075 -58.315 ;
        RECT -29.405 -60.005 -29.075 -59.675 ;
        RECT -29.405 -61.365 -29.075 -61.035 ;
        RECT -29.405 -62.725 -29.075 -62.395 ;
        RECT -29.405 -64.085 -29.075 -63.755 ;
        RECT -29.405 -65.445 -29.075 -65.115 ;
        RECT -29.405 -66.805 -29.075 -66.475 ;
        RECT -29.405 -68.165 -29.075 -67.835 ;
        RECT -29.405 -69.525 -29.075 -69.195 ;
        RECT -29.405 -70.885 -29.075 -70.555 ;
        RECT -29.405 -72.245 -29.075 -71.915 ;
        RECT -29.405 -73.605 -29.075 -73.275 ;
        RECT -29.405 -74.965 -29.075 -74.635 ;
        RECT -29.405 -76.325 -29.075 -75.995 ;
        RECT -29.405 -77.685 -29.075 -77.355 ;
        RECT -29.405 -79.045 -29.075 -78.715 ;
        RECT -29.405 -80.405 -29.075 -80.075 ;
        RECT -29.405 -81.765 -29.075 -81.435 ;
        RECT -29.405 -83.125 -29.075 -82.795 ;
        RECT -29.405 -84.485 -29.075 -84.155 ;
        RECT -29.405 -85.845 -29.075 -85.515 ;
        RECT -29.405 -87.205 -29.075 -86.875 ;
        RECT -29.405 -88.565 -29.075 -88.235 ;
        RECT -29.405 -89.925 -29.075 -89.595 ;
        RECT -29.405 -91.285 -29.075 -90.955 ;
        RECT -29.405 -92.645 -29.075 -92.315 ;
        RECT -29.405 -94.005 -29.075 -93.675 ;
        RECT -29.405 -95.365 -29.075 -95.035 ;
        RECT -29.405 -96.725 -29.075 -96.395 ;
        RECT -29.405 -98.085 -29.075 -97.755 ;
        RECT -29.405 -99.445 -29.075 -99.115 ;
        RECT -29.405 -100.805 -29.075 -100.475 ;
        RECT -29.405 -102.165 -29.075 -101.835 ;
        RECT -29.405 -103.525 -29.075 -103.195 ;
        RECT -29.405 -108.965 -29.075 -108.635 ;
        RECT -29.405 -110.325 -29.075 -109.995 ;
        RECT -29.405 -113.045 -29.075 -112.715 ;
        RECT -29.405 -114.405 -29.075 -114.075 ;
        RECT -29.405 -115.765 -29.075 -115.435 ;
        RECT -29.405 -117.125 -29.075 -116.795 ;
        RECT -29.405 -118.485 -29.075 -118.155 ;
        RECT -29.405 -119.79 -29.075 -119.46 ;
        RECT -29.405 -121.205 -29.075 -120.875 ;
        RECT -29.405 -122.565 -29.075 -122.235 ;
        RECT -29.405 -123.925 -29.075 -123.595 ;
        RECT -29.405 -126.645 -29.075 -126.315 ;
        RECT -29.405 -128.43 -29.075 -128.1 ;
        RECT -29.405 -129.365 -29.075 -129.035 ;
        RECT -29.405 -130.725 -29.075 -130.395 ;
        RECT -29.4 -132.08 -29.08 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.405 -212.325 -29.075 -211.995 ;
        RECT -29.405 -213.625 -29.075 -213.295 ;
        RECT -29.405 -215.045 -29.075 -214.715 ;
        RECT -29.405 -216.405 -29.075 -216.075 ;
        RECT -29.405 -217.765 -29.075 -217.435 ;
        RECT -29.405 -219.125 -29.075 -218.795 ;
        RECT -29.405 -221.37 -29.075 -220.24 ;
        RECT -29.4 -221.485 -29.08 -211.995 ;
    END
    PORT
      LAYER met3 ;
        RECT -28.045 -117.125 -27.715 -116.795 ;
        RECT -28.045 -118.485 -27.715 -118.155 ;
        RECT -28.045 -119.79 -27.715 -119.46 ;
        RECT -28.045 -121.205 -27.715 -120.875 ;
        RECT -28.045 -122.565 -27.715 -122.235 ;
        RECT -28.045 -123.925 -27.715 -123.595 ;
        RECT -28.045 -126.645 -27.715 -126.315 ;
        RECT -28.045 -128.43 -27.715 -128.1 ;
        RECT -28.045 -129.365 -27.715 -129.035 ;
        RECT -28.045 -130.725 -27.715 -130.395 ;
        RECT -28.045 -133.445 -27.715 -133.115 ;
        RECT -28.045 -134.805 -27.715 -134.475 ;
        RECT -28.045 -136.165 -27.715 -135.835 ;
        RECT -28.045 -137.525 -27.715 -137.195 ;
        RECT -28.045 -140.245 -27.715 -139.915 ;
        RECT -28.045 -142.965 -27.715 -142.635 ;
        RECT -28.045 -144.325 -27.715 -143.995 ;
        RECT -28.045 -145.685 -27.715 -145.355 ;
        RECT -28.045 -147.045 -27.715 -146.715 ;
        RECT -28.045 -148.405 -27.715 -148.075 ;
        RECT -28.045 -149.765 -27.715 -149.435 ;
        RECT -28.045 -151.125 -27.715 -150.795 ;
        RECT -28.045 -152.485 -27.715 -152.155 ;
        RECT -28.045 -153.845 -27.715 -153.515 ;
        RECT -28.045 -155.205 -27.715 -154.875 ;
        RECT -28.045 -156.565 -27.715 -156.235 ;
        RECT -28.045 -157.925 -27.715 -157.595 ;
        RECT -28.045 -159.285 -27.715 -158.955 ;
        RECT -28.045 -160.645 -27.715 -160.315 ;
        RECT -28.045 -162.005 -27.715 -161.675 ;
        RECT -28.045 -163.365 -27.715 -163.035 ;
        RECT -28.045 -164.725 -27.715 -164.395 ;
        RECT -28.045 -166.085 -27.715 -165.755 ;
        RECT -28.045 -167.445 -27.715 -167.115 ;
        RECT -28.045 -171.525 -27.715 -171.195 ;
        RECT -28.045 -172.885 -27.715 -172.555 ;
        RECT -28.045 -174.245 -27.715 -173.915 ;
        RECT -28.045 -175.605 -27.715 -175.275 ;
        RECT -28.045 -176.965 -27.715 -176.635 ;
        RECT -28.045 -179.685 -27.715 -179.355 ;
        RECT -28.045 -181.045 -27.715 -180.715 ;
        RECT -28.045 -182.405 -27.715 -182.075 ;
        RECT -28.045 -183.765 -27.715 -183.435 ;
        RECT -28.045 -185.125 -27.715 -184.795 ;
        RECT -28.045 -186.485 -27.715 -186.155 ;
        RECT -28.045 -189.205 -27.715 -188.875 ;
        RECT -28.045 -190.565 -27.715 -190.235 ;
        RECT -28.045 -196.005 -27.715 -195.675 ;
        RECT -28.045 -197.365 -27.715 -197.035 ;
        RECT -28.045 -198.725 -27.715 -198.395 ;
        RECT -28.045 -200.085 -27.715 -199.755 ;
        RECT -28.045 -201.445 -27.715 -201.115 ;
        RECT -28.045 -202.805 -27.715 -202.475 ;
        RECT -28.045 -204.165 -27.715 -203.835 ;
        RECT -28.045 -205.525 -27.715 -205.195 ;
        RECT -28.045 -208.245 -27.715 -207.915 ;
        RECT -28.04 -209.6 -27.72 131.045 ;
        RECT -28.045 129.8 -27.715 130.93 ;
        RECT -28.045 127.675 -27.715 128.005 ;
        RECT -28.045 126.315 -27.715 126.645 ;
        RECT -28.045 124.955 -27.715 125.285 ;
        RECT -28.045 123.595 -27.715 123.925 ;
        RECT -28.045 122.235 -27.715 122.565 ;
        RECT -28.045 120.875 -27.715 121.205 ;
        RECT -28.045 119.515 -27.715 119.845 ;
        RECT -28.045 118.155 -27.715 118.485 ;
        RECT -28.045 116.795 -27.715 117.125 ;
        RECT -28.045 115.435 -27.715 115.765 ;
        RECT -28.045 114.075 -27.715 114.405 ;
        RECT -28.045 112.715 -27.715 113.045 ;
        RECT -28.045 111.355 -27.715 111.685 ;
        RECT -28.045 109.995 -27.715 110.325 ;
        RECT -28.045 108.635 -27.715 108.965 ;
        RECT -28.045 107.275 -27.715 107.605 ;
        RECT -28.045 105.915 -27.715 106.245 ;
        RECT -28.045 104.555 -27.715 104.885 ;
        RECT -28.045 103.195 -27.715 103.525 ;
        RECT -28.045 101.835 -27.715 102.165 ;
        RECT -28.045 100.475 -27.715 100.805 ;
        RECT -28.045 99.115 -27.715 99.445 ;
        RECT -28.045 97.755 -27.715 98.085 ;
        RECT -28.045 96.395 -27.715 96.725 ;
        RECT -28.045 95.035 -27.715 95.365 ;
        RECT -28.045 93.675 -27.715 94.005 ;
        RECT -28.045 92.315 -27.715 92.645 ;
        RECT -28.045 90.955 -27.715 91.285 ;
        RECT -28.045 89.595 -27.715 89.925 ;
        RECT -28.045 88.235 -27.715 88.565 ;
        RECT -28.045 86.875 -27.715 87.205 ;
        RECT -28.045 85.515 -27.715 85.845 ;
        RECT -28.045 84.155 -27.715 84.485 ;
        RECT -28.045 82.795 -27.715 83.125 ;
        RECT -28.045 81.435 -27.715 81.765 ;
        RECT -28.045 80.075 -27.715 80.405 ;
        RECT -28.045 78.715 -27.715 79.045 ;
        RECT -28.045 77.355 -27.715 77.685 ;
        RECT -28.045 75.995 -27.715 76.325 ;
        RECT -28.045 74.635 -27.715 74.965 ;
        RECT -28.045 73.275 -27.715 73.605 ;
        RECT -28.045 71.915 -27.715 72.245 ;
        RECT -28.045 70.555 -27.715 70.885 ;
        RECT -28.045 69.195 -27.715 69.525 ;
        RECT -28.045 67.835 -27.715 68.165 ;
        RECT -28.045 66.475 -27.715 66.805 ;
        RECT -28.045 65.115 -27.715 65.445 ;
        RECT -28.045 63.755 -27.715 64.085 ;
        RECT -28.045 62.395 -27.715 62.725 ;
        RECT -28.045 61.035 -27.715 61.365 ;
        RECT -28.045 59.675 -27.715 60.005 ;
        RECT -28.045 58.315 -27.715 58.645 ;
        RECT -28.045 56.955 -27.715 57.285 ;
        RECT -28.045 55.595 -27.715 55.925 ;
        RECT -28.045 54.235 -27.715 54.565 ;
        RECT -28.045 52.875 -27.715 53.205 ;
        RECT -28.045 51.515 -27.715 51.845 ;
        RECT -28.045 50.155 -27.715 50.485 ;
        RECT -28.045 48.795 -27.715 49.125 ;
        RECT -28.045 47.435 -27.715 47.765 ;
        RECT -28.045 46.075 -27.715 46.405 ;
        RECT -28.045 44.715 -27.715 45.045 ;
        RECT -28.045 43.355 -27.715 43.685 ;
        RECT -28.045 41.995 -27.715 42.325 ;
        RECT -28.045 40.635 -27.715 40.965 ;
        RECT -28.045 39.275 -27.715 39.605 ;
        RECT -28.045 37.915 -27.715 38.245 ;
        RECT -28.045 36.555 -27.715 36.885 ;
        RECT -28.045 35.195 -27.715 35.525 ;
        RECT -28.045 33.835 -27.715 34.165 ;
        RECT -28.045 32.475 -27.715 32.805 ;
        RECT -28.045 31.115 -27.715 31.445 ;
        RECT -28.045 29.755 -27.715 30.085 ;
        RECT -28.045 28.395 -27.715 28.725 ;
        RECT -28.045 27.035 -27.715 27.365 ;
        RECT -28.045 25.675 -27.715 26.005 ;
        RECT -28.045 24.315 -27.715 24.645 ;
        RECT -28.045 22.955 -27.715 23.285 ;
        RECT -28.045 21.595 -27.715 21.925 ;
        RECT -28.045 20.235 -27.715 20.565 ;
        RECT -28.045 18.875 -27.715 19.205 ;
        RECT -28.045 17.515 -27.715 17.845 ;
        RECT -28.045 16.155 -27.715 16.485 ;
        RECT -28.045 14.795 -27.715 15.125 ;
        RECT -28.045 13.435 -27.715 13.765 ;
        RECT -28.045 12.075 -27.715 12.405 ;
        RECT -28.045 10.715 -27.715 11.045 ;
        RECT -28.045 9.355 -27.715 9.685 ;
        RECT -28.045 7.995 -27.715 8.325 ;
        RECT -28.045 6.635 -27.715 6.965 ;
        RECT -28.045 5.275 -27.715 5.605 ;
        RECT -28.045 3.915 -27.715 4.245 ;
        RECT -28.045 2.555 -27.715 2.885 ;
        RECT -28.045 1.195 -27.715 1.525 ;
        RECT -28.045 -0.165 -27.715 0.165 ;
        RECT -28.045 -8.325 -27.715 -7.995 ;
        RECT -28.045 -9.685 -27.715 -9.355 ;
        RECT -28.045 -11.16 -27.715 -10.83 ;
        RECT -28.045 -12.405 -27.715 -12.075 ;
        RECT -28.045 -15.125 -27.715 -14.795 ;
        RECT -28.045 -16.25 -27.715 -15.92 ;
        RECT -28.045 -27.365 -27.715 -27.035 ;
        RECT -28.045 -30.085 -27.715 -29.755 ;
        RECT -28.045 -32.34 -27.715 -32.01 ;
        RECT -28.045 -37.43 -27.715 -37.1 ;
        RECT -28.045 -43.685 -27.715 -43.355 ;
        RECT -28.045 -45.045 -27.715 -44.715 ;
        RECT -28.045 -46.405 -27.715 -46.075 ;
        RECT -28.045 -47.765 -27.715 -47.435 ;
        RECT -28.045 -49.125 -27.715 -48.795 ;
        RECT -28.045 -50.485 -27.715 -50.155 ;
        RECT -28.045 -51.845 -27.715 -51.515 ;
        RECT -28.045 -53.205 -27.715 -52.875 ;
        RECT -28.045 -54.565 -27.715 -54.235 ;
        RECT -28.045 -55.925 -27.715 -55.595 ;
        RECT -28.045 -57.285 -27.715 -56.955 ;
        RECT -28.045 -58.645 -27.715 -58.315 ;
        RECT -28.045 -60.005 -27.715 -59.675 ;
        RECT -28.045 -61.365 -27.715 -61.035 ;
        RECT -28.045 -62.725 -27.715 -62.395 ;
        RECT -28.045 -64.085 -27.715 -63.755 ;
        RECT -28.045 -65.445 -27.715 -65.115 ;
        RECT -28.045 -66.805 -27.715 -66.475 ;
        RECT -28.045 -68.165 -27.715 -67.835 ;
        RECT -28.045 -69.525 -27.715 -69.195 ;
        RECT -28.045 -70.885 -27.715 -70.555 ;
        RECT -28.045 -72.245 -27.715 -71.915 ;
        RECT -28.045 -73.605 -27.715 -73.275 ;
        RECT -28.045 -74.965 -27.715 -74.635 ;
        RECT -28.045 -76.325 -27.715 -75.995 ;
        RECT -28.045 -77.685 -27.715 -77.355 ;
        RECT -28.045 -79.045 -27.715 -78.715 ;
        RECT -28.045 -80.405 -27.715 -80.075 ;
        RECT -28.045 -81.765 -27.715 -81.435 ;
        RECT -28.045 -83.125 -27.715 -82.795 ;
        RECT -28.045 -84.485 -27.715 -84.155 ;
        RECT -28.045 -85.845 -27.715 -85.515 ;
        RECT -28.045 -87.205 -27.715 -86.875 ;
        RECT -28.045 -88.565 -27.715 -88.235 ;
        RECT -28.045 -89.925 -27.715 -89.595 ;
        RECT -28.045 -91.285 -27.715 -90.955 ;
        RECT -28.045 -92.645 -27.715 -92.315 ;
        RECT -28.045 -94.005 -27.715 -93.675 ;
        RECT -28.045 -95.365 -27.715 -95.035 ;
        RECT -28.045 -96.725 -27.715 -96.395 ;
        RECT -28.045 -98.085 -27.715 -97.755 ;
        RECT -28.045 -99.445 -27.715 -99.115 ;
        RECT -28.045 -100.805 -27.715 -100.475 ;
        RECT -28.045 -102.165 -27.715 -101.835 ;
        RECT -28.045 -103.525 -27.715 -103.195 ;
        RECT -28.045 -108.965 -27.715 -108.635 ;
        RECT -28.045 -110.325 -27.715 -109.995 ;
        RECT -28.045 -113.045 -27.715 -112.715 ;
        RECT -28.045 -114.405 -27.715 -114.075 ;
        RECT -28.045 -115.765 -27.715 -115.435 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.925 129.8 -38.595 130.93 ;
        RECT -38.925 127.675 -38.595 128.005 ;
        RECT -38.925 126.315 -38.595 126.645 ;
        RECT -38.925 124.955 -38.595 125.285 ;
        RECT -38.925 123.595 -38.595 123.925 ;
        RECT -38.925 122.235 -38.595 122.565 ;
        RECT -38.925 120.875 -38.595 121.205 ;
        RECT -38.925 119.515 -38.595 119.845 ;
        RECT -38.925 118.155 -38.595 118.485 ;
        RECT -38.925 116.795 -38.595 117.125 ;
        RECT -38.925 115.435 -38.595 115.765 ;
        RECT -38.925 114.075 -38.595 114.405 ;
        RECT -38.925 112.715 -38.595 113.045 ;
        RECT -38.925 111.355 -38.595 111.685 ;
        RECT -38.925 109.995 -38.595 110.325 ;
        RECT -38.925 108.635 -38.595 108.965 ;
        RECT -38.925 107.275 -38.595 107.605 ;
        RECT -38.925 105.915 -38.595 106.245 ;
        RECT -38.925 104.555 -38.595 104.885 ;
        RECT -38.925 103.195 -38.595 103.525 ;
        RECT -38.925 101.835 -38.595 102.165 ;
        RECT -38.925 100.475 -38.595 100.805 ;
        RECT -38.925 99.115 -38.595 99.445 ;
        RECT -38.925 97.755 -38.595 98.085 ;
        RECT -38.925 96.395 -38.595 96.725 ;
        RECT -38.925 95.035 -38.595 95.365 ;
        RECT -38.925 93.675 -38.595 94.005 ;
        RECT -38.925 92.315 -38.595 92.645 ;
        RECT -38.925 90.955 -38.595 91.285 ;
        RECT -38.925 89.595 -38.595 89.925 ;
        RECT -38.925 88.235 -38.595 88.565 ;
        RECT -38.925 86.875 -38.595 87.205 ;
        RECT -38.925 85.515 -38.595 85.845 ;
        RECT -38.925 84.155 -38.595 84.485 ;
        RECT -38.925 82.795 -38.595 83.125 ;
        RECT -38.925 81.435 -38.595 81.765 ;
        RECT -38.925 80.075 -38.595 80.405 ;
        RECT -38.925 78.715 -38.595 79.045 ;
        RECT -38.925 77.355 -38.595 77.685 ;
        RECT -38.925 75.995 -38.595 76.325 ;
        RECT -38.925 74.635 -38.595 74.965 ;
        RECT -38.925 73.275 -38.595 73.605 ;
        RECT -38.925 71.915 -38.595 72.245 ;
        RECT -38.925 70.555 -38.595 70.885 ;
        RECT -38.925 69.195 -38.595 69.525 ;
        RECT -38.925 67.835 -38.595 68.165 ;
        RECT -38.925 66.475 -38.595 66.805 ;
        RECT -38.925 65.115 -38.595 65.445 ;
        RECT -38.925 63.755 -38.595 64.085 ;
        RECT -38.925 62.395 -38.595 62.725 ;
        RECT -38.925 61.035 -38.595 61.365 ;
        RECT -38.925 59.675 -38.595 60.005 ;
        RECT -38.925 58.315 -38.595 58.645 ;
        RECT -38.925 56.955 -38.595 57.285 ;
        RECT -38.925 55.595 -38.595 55.925 ;
        RECT -38.925 54.235 -38.595 54.565 ;
        RECT -38.925 52.875 -38.595 53.205 ;
        RECT -38.925 51.515 -38.595 51.845 ;
        RECT -38.925 50.155 -38.595 50.485 ;
        RECT -38.925 48.795 -38.595 49.125 ;
        RECT -38.925 47.435 -38.595 47.765 ;
        RECT -38.925 46.075 -38.595 46.405 ;
        RECT -38.925 44.715 -38.595 45.045 ;
        RECT -38.925 43.355 -38.595 43.685 ;
        RECT -38.925 41.995 -38.595 42.325 ;
        RECT -38.925 40.635 -38.595 40.965 ;
        RECT -38.925 39.275 -38.595 39.605 ;
        RECT -38.925 37.915 -38.595 38.245 ;
        RECT -38.925 36.555 -38.595 36.885 ;
        RECT -38.925 35.195 -38.595 35.525 ;
        RECT -38.925 33.835 -38.595 34.165 ;
        RECT -38.925 32.475 -38.595 32.805 ;
        RECT -38.925 31.115 -38.595 31.445 ;
        RECT -38.925 29.755 -38.595 30.085 ;
        RECT -38.925 28.395 -38.595 28.725 ;
        RECT -38.925 27.035 -38.595 27.365 ;
        RECT -38.925 25.675 -38.595 26.005 ;
        RECT -38.925 24.315 -38.595 24.645 ;
        RECT -38.925 22.955 -38.595 23.285 ;
        RECT -38.925 21.595 -38.595 21.925 ;
        RECT -38.925 20.235 -38.595 20.565 ;
        RECT -38.925 18.875 -38.595 19.205 ;
        RECT -38.925 17.515 -38.595 17.845 ;
        RECT -38.925 16.155 -38.595 16.485 ;
        RECT -38.925 14.795 -38.595 15.125 ;
        RECT -38.925 13.435 -38.595 13.765 ;
        RECT -38.925 12.075 -38.595 12.405 ;
        RECT -38.925 10.715 -38.595 11.045 ;
        RECT -38.925 9.355 -38.595 9.685 ;
        RECT -38.925 7.995 -38.595 8.325 ;
        RECT -38.925 6.635 -38.595 6.965 ;
        RECT -38.925 5.275 -38.595 5.605 ;
        RECT -38.925 3.915 -38.595 4.245 ;
        RECT -38.925 2.555 -38.595 2.885 ;
        RECT -38.925 1.195 -38.595 1.525 ;
        RECT -38.925 -0.165 -38.595 0.165 ;
        RECT -38.925 -1.525 -38.595 -1.195 ;
        RECT -38.925 -2.885 -38.595 -2.555 ;
        RECT -38.925 -4.245 -38.595 -3.915 ;
        RECT -38.925 -5.605 -38.595 -5.275 ;
        RECT -38.925 -6.965 -38.595 -6.635 ;
        RECT -38.925 -8.325 -38.595 -7.995 ;
        RECT -38.925 -9.685 -38.595 -9.355 ;
        RECT -38.925 -11.045 -38.595 -10.715 ;
        RECT -38.925 -12.405 -38.595 -12.075 ;
        RECT -38.925 -13.765 -38.595 -13.435 ;
        RECT -38.925 -15.125 -38.595 -14.795 ;
        RECT -38.925 -16.485 -38.595 -16.155 ;
        RECT -38.925 -17.845 -38.595 -17.515 ;
        RECT -38.925 -19.205 -38.595 -18.875 ;
        RECT -38.925 -20.565 -38.595 -20.235 ;
        RECT -38.925 -27.365 -38.595 -27.035 ;
        RECT -38.925 -28.725 -38.595 -28.395 ;
        RECT -38.925 -30.085 -38.595 -29.755 ;
        RECT -38.925 -32.805 -38.595 -32.475 ;
        RECT -38.925 -35.525 -38.595 -35.195 ;
        RECT -38.925 -36.885 -38.595 -36.555 ;
        RECT -38.925 -39.605 -38.595 -39.275 ;
        RECT -38.925 -40.965 -38.595 -40.635 ;
        RECT -38.925 -42.325 -38.595 -41.995 ;
        RECT -38.925 -43.685 -38.595 -43.355 ;
        RECT -38.925 -45.045 -38.595 -44.715 ;
        RECT -38.925 -46.405 -38.595 -46.075 ;
        RECT -38.925 -47.765 -38.595 -47.435 ;
        RECT -38.925 -49.125 -38.595 -48.795 ;
        RECT -38.925 -50.485 -38.595 -50.155 ;
        RECT -38.925 -51.845 -38.595 -51.515 ;
        RECT -38.925 -53.205 -38.595 -52.875 ;
        RECT -38.925 -54.565 -38.595 -54.235 ;
        RECT -38.925 -55.925 -38.595 -55.595 ;
        RECT -38.925 -57.285 -38.595 -56.955 ;
        RECT -38.925 -58.645 -38.595 -58.315 ;
        RECT -38.925 -60.005 -38.595 -59.675 ;
        RECT -38.925 -61.365 -38.595 -61.035 ;
        RECT -38.925 -62.725 -38.595 -62.395 ;
        RECT -38.925 -64.085 -38.595 -63.755 ;
        RECT -38.925 -65.445 -38.595 -65.115 ;
        RECT -38.925 -66.805 -38.595 -66.475 ;
        RECT -38.925 -68.165 -38.595 -67.835 ;
        RECT -38.925 -69.525 -38.595 -69.195 ;
        RECT -38.925 -70.885 -38.595 -70.555 ;
        RECT -38.925 -72.245 -38.595 -71.915 ;
        RECT -38.925 -73.605 -38.595 -73.275 ;
        RECT -38.925 -74.965 -38.595 -74.635 ;
        RECT -38.925 -76.325 -38.595 -75.995 ;
        RECT -38.925 -77.685 -38.595 -77.355 ;
        RECT -38.925 -79.045 -38.595 -78.715 ;
        RECT -38.925 -80.405 -38.595 -80.075 ;
        RECT -38.925 -81.765 -38.595 -81.435 ;
        RECT -38.925 -83.125 -38.595 -82.795 ;
        RECT -38.925 -84.485 -38.595 -84.155 ;
        RECT -38.925 -85.845 -38.595 -85.515 ;
        RECT -38.925 -87.205 -38.595 -86.875 ;
        RECT -38.925 -88.565 -38.595 -88.235 ;
        RECT -38.925 -89.925 -38.595 -89.595 ;
        RECT -38.925 -91.285 -38.595 -90.955 ;
        RECT -38.925 -92.645 -38.595 -92.315 ;
        RECT -38.925 -94.005 -38.595 -93.675 ;
        RECT -38.925 -95.365 -38.595 -95.035 ;
        RECT -38.925 -96.725 -38.595 -96.395 ;
        RECT -38.925 -98.085 -38.595 -97.755 ;
        RECT -38.925 -99.445 -38.595 -99.115 ;
        RECT -38.925 -100.805 -38.595 -100.475 ;
        RECT -38.925 -102.165 -38.595 -101.835 ;
        RECT -38.925 -103.525 -38.595 -103.195 ;
        RECT -38.925 -104.885 -38.595 -104.555 ;
        RECT -38.925 -106.245 -38.595 -105.915 ;
        RECT -38.925 -108.965 -38.595 -108.635 ;
        RECT -38.925 -110.325 -38.595 -109.995 ;
        RECT -38.925 -113.045 -38.595 -112.715 ;
        RECT -38.925 -114.405 -38.595 -114.075 ;
        RECT -38.925 -115.765 -38.595 -115.435 ;
        RECT -38.925 -117.125 -38.595 -116.795 ;
        RECT -38.925 -118.485 -38.595 -118.155 ;
        RECT -38.925 -119.79 -38.595 -119.46 ;
        RECT -38.925 -121.205 -38.595 -120.875 ;
        RECT -38.925 -122.565 -38.595 -122.235 ;
        RECT -38.925 -123.925 -38.595 -123.595 ;
        RECT -38.925 -126.645 -38.595 -126.315 ;
        RECT -38.925 -128.43 -38.595 -128.1 ;
        RECT -38.925 -129.365 -38.595 -129.035 ;
        RECT -38.925 -130.725 -38.595 -130.395 ;
        RECT -38.92 -132.08 -38.6 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.925 -212.325 -38.595 -211.995 ;
        RECT -38.925 -213.625 -38.595 -213.295 ;
        RECT -38.925 -215.045 -38.595 -214.715 ;
        RECT -38.925 -216.405 -38.595 -216.075 ;
        RECT -38.925 -217.765 -38.595 -217.435 ;
        RECT -38.925 -219.125 -38.595 -218.795 ;
        RECT -38.925 -221.37 -38.595 -220.24 ;
        RECT -38.92 -221.485 -38.6 -211.995 ;
    END
    PORT
      LAYER met3 ;
        RECT -37.565 129.8 -37.235 130.93 ;
        RECT -37.565 127.675 -37.235 128.005 ;
        RECT -37.565 126.315 -37.235 126.645 ;
        RECT -37.565 124.955 -37.235 125.285 ;
        RECT -37.565 123.595 -37.235 123.925 ;
        RECT -37.565 122.235 -37.235 122.565 ;
        RECT -37.565 120.875 -37.235 121.205 ;
        RECT -37.565 119.515 -37.235 119.845 ;
        RECT -37.565 118.155 -37.235 118.485 ;
        RECT -37.565 116.795 -37.235 117.125 ;
        RECT -37.565 115.435 -37.235 115.765 ;
        RECT -37.565 114.075 -37.235 114.405 ;
        RECT -37.565 112.715 -37.235 113.045 ;
        RECT -37.565 111.355 -37.235 111.685 ;
        RECT -37.565 109.995 -37.235 110.325 ;
        RECT -37.565 108.635 -37.235 108.965 ;
        RECT -37.565 107.275 -37.235 107.605 ;
        RECT -37.565 105.915 -37.235 106.245 ;
        RECT -37.565 104.555 -37.235 104.885 ;
        RECT -37.565 103.195 -37.235 103.525 ;
        RECT -37.565 101.835 -37.235 102.165 ;
        RECT -37.565 100.475 -37.235 100.805 ;
        RECT -37.565 99.115 -37.235 99.445 ;
        RECT -37.565 97.755 -37.235 98.085 ;
        RECT -37.565 96.395 -37.235 96.725 ;
        RECT -37.565 95.035 -37.235 95.365 ;
        RECT -37.565 93.675 -37.235 94.005 ;
        RECT -37.565 92.315 -37.235 92.645 ;
        RECT -37.565 90.955 -37.235 91.285 ;
        RECT -37.565 89.595 -37.235 89.925 ;
        RECT -37.565 88.235 -37.235 88.565 ;
        RECT -37.565 86.875 -37.235 87.205 ;
        RECT -37.565 85.515 -37.235 85.845 ;
        RECT -37.565 84.155 -37.235 84.485 ;
        RECT -37.565 82.795 -37.235 83.125 ;
        RECT -37.565 81.435 -37.235 81.765 ;
        RECT -37.565 80.075 -37.235 80.405 ;
        RECT -37.565 78.715 -37.235 79.045 ;
        RECT -37.565 77.355 -37.235 77.685 ;
        RECT -37.565 75.995 -37.235 76.325 ;
        RECT -37.565 74.635 -37.235 74.965 ;
        RECT -37.565 73.275 -37.235 73.605 ;
        RECT -37.565 71.915 -37.235 72.245 ;
        RECT -37.565 70.555 -37.235 70.885 ;
        RECT -37.565 69.195 -37.235 69.525 ;
        RECT -37.565 67.835 -37.235 68.165 ;
        RECT -37.565 66.475 -37.235 66.805 ;
        RECT -37.565 65.115 -37.235 65.445 ;
        RECT -37.565 63.755 -37.235 64.085 ;
        RECT -37.565 62.395 -37.235 62.725 ;
        RECT -37.565 61.035 -37.235 61.365 ;
        RECT -37.565 59.675 -37.235 60.005 ;
        RECT -37.565 58.315 -37.235 58.645 ;
        RECT -37.565 56.955 -37.235 57.285 ;
        RECT -37.565 55.595 -37.235 55.925 ;
        RECT -37.565 54.235 -37.235 54.565 ;
        RECT -37.565 52.875 -37.235 53.205 ;
        RECT -37.565 51.515 -37.235 51.845 ;
        RECT -37.565 50.155 -37.235 50.485 ;
        RECT -37.565 48.795 -37.235 49.125 ;
        RECT -37.565 47.435 -37.235 47.765 ;
        RECT -37.565 46.075 -37.235 46.405 ;
        RECT -37.565 44.715 -37.235 45.045 ;
        RECT -37.565 43.355 -37.235 43.685 ;
        RECT -37.565 41.995 -37.235 42.325 ;
        RECT -37.565 40.635 -37.235 40.965 ;
        RECT -37.565 39.275 -37.235 39.605 ;
        RECT -37.565 37.915 -37.235 38.245 ;
        RECT -37.565 36.555 -37.235 36.885 ;
        RECT -37.565 35.195 -37.235 35.525 ;
        RECT -37.565 33.835 -37.235 34.165 ;
        RECT -37.565 32.475 -37.235 32.805 ;
        RECT -37.565 31.115 -37.235 31.445 ;
        RECT -37.565 29.755 -37.235 30.085 ;
        RECT -37.565 28.395 -37.235 28.725 ;
        RECT -37.565 27.035 -37.235 27.365 ;
        RECT -37.565 25.675 -37.235 26.005 ;
        RECT -37.565 24.315 -37.235 24.645 ;
        RECT -37.565 22.955 -37.235 23.285 ;
        RECT -37.565 21.595 -37.235 21.925 ;
        RECT -37.565 20.235 -37.235 20.565 ;
        RECT -37.565 18.875 -37.235 19.205 ;
        RECT -37.565 17.515 -37.235 17.845 ;
        RECT -37.565 16.155 -37.235 16.485 ;
        RECT -37.565 14.795 -37.235 15.125 ;
        RECT -37.565 13.435 -37.235 13.765 ;
        RECT -37.565 12.075 -37.235 12.405 ;
        RECT -37.565 10.715 -37.235 11.045 ;
        RECT -37.565 9.355 -37.235 9.685 ;
        RECT -37.565 7.995 -37.235 8.325 ;
        RECT -37.565 6.635 -37.235 6.965 ;
        RECT -37.565 5.275 -37.235 5.605 ;
        RECT -37.565 3.915 -37.235 4.245 ;
        RECT -37.565 2.555 -37.235 2.885 ;
        RECT -37.565 1.195 -37.235 1.525 ;
        RECT -37.565 -0.165 -37.235 0.165 ;
        RECT -37.565 -1.525 -37.235 -1.195 ;
        RECT -37.565 -2.885 -37.235 -2.555 ;
        RECT -37.565 -4.245 -37.235 -3.915 ;
        RECT -37.565 -6.965 -37.235 -6.635 ;
        RECT -37.565 -8.325 -37.235 -7.995 ;
        RECT -37.565 -9.685 -37.235 -9.355 ;
        RECT -37.565 -11.045 -37.235 -10.715 ;
        RECT -37.565 -12.405 -37.235 -12.075 ;
        RECT -37.565 -13.765 -37.235 -13.435 ;
        RECT -37.565 -15.125 -37.235 -14.795 ;
        RECT -37.565 -16.485 -37.235 -16.155 ;
        RECT -37.565 -17.845 -37.235 -17.515 ;
        RECT -37.565 -19.205 -37.235 -18.875 ;
        RECT -37.565 -20.565 -37.235 -20.235 ;
        RECT -37.565 -27.365 -37.235 -27.035 ;
        RECT -37.565 -28.725 -37.235 -28.395 ;
        RECT -37.565 -30.085 -37.235 -29.755 ;
        RECT -37.565 -32.805 -37.235 -32.475 ;
        RECT -37.565 -35.525 -37.235 -35.195 ;
        RECT -37.565 -36.885 -37.235 -36.555 ;
        RECT -37.565 -39.605 -37.235 -39.275 ;
        RECT -37.565 -40.965 -37.235 -40.635 ;
        RECT -37.565 -42.325 -37.235 -41.995 ;
        RECT -37.565 -43.685 -37.235 -43.355 ;
        RECT -37.565 -45.045 -37.235 -44.715 ;
        RECT -37.565 -46.405 -37.235 -46.075 ;
        RECT -37.565 -47.765 -37.235 -47.435 ;
        RECT -37.565 -49.125 -37.235 -48.795 ;
        RECT -37.565 -50.485 -37.235 -50.155 ;
        RECT -37.565 -51.845 -37.235 -51.515 ;
        RECT -37.565 -53.205 -37.235 -52.875 ;
        RECT -37.565 -54.565 -37.235 -54.235 ;
        RECT -37.565 -55.925 -37.235 -55.595 ;
        RECT -37.565 -57.285 -37.235 -56.955 ;
        RECT -37.565 -58.645 -37.235 -58.315 ;
        RECT -37.565 -60.005 -37.235 -59.675 ;
        RECT -37.565 -61.365 -37.235 -61.035 ;
        RECT -37.565 -62.725 -37.235 -62.395 ;
        RECT -37.565 -64.085 -37.235 -63.755 ;
        RECT -37.565 -65.445 -37.235 -65.115 ;
        RECT -37.565 -66.805 -37.235 -66.475 ;
        RECT -37.565 -68.165 -37.235 -67.835 ;
        RECT -37.565 -69.525 -37.235 -69.195 ;
        RECT -37.565 -70.885 -37.235 -70.555 ;
        RECT -37.565 -72.245 -37.235 -71.915 ;
        RECT -37.565 -73.605 -37.235 -73.275 ;
        RECT -37.565 -74.965 -37.235 -74.635 ;
        RECT -37.565 -76.325 -37.235 -75.995 ;
        RECT -37.565 -77.685 -37.235 -77.355 ;
        RECT -37.565 -79.045 -37.235 -78.715 ;
        RECT -37.565 -80.405 -37.235 -80.075 ;
        RECT -37.565 -81.765 -37.235 -81.435 ;
        RECT -37.565 -83.125 -37.235 -82.795 ;
        RECT -37.565 -84.485 -37.235 -84.155 ;
        RECT -37.565 -85.845 -37.235 -85.515 ;
        RECT -37.565 -87.205 -37.235 -86.875 ;
        RECT -37.565 -88.565 -37.235 -88.235 ;
        RECT -37.565 -89.925 -37.235 -89.595 ;
        RECT -37.565 -91.285 -37.235 -90.955 ;
        RECT -37.565 -92.645 -37.235 -92.315 ;
        RECT -37.565 -94.005 -37.235 -93.675 ;
        RECT -37.565 -95.365 -37.235 -95.035 ;
        RECT -37.565 -96.725 -37.235 -96.395 ;
        RECT -37.565 -98.085 -37.235 -97.755 ;
        RECT -37.565 -99.445 -37.235 -99.115 ;
        RECT -37.565 -100.805 -37.235 -100.475 ;
        RECT -37.565 -102.165 -37.235 -101.835 ;
        RECT -37.565 -103.525 -37.235 -103.195 ;
        RECT -37.565 -104.885 -37.235 -104.555 ;
        RECT -37.565 -106.245 -37.235 -105.915 ;
        RECT -37.565 -108.965 -37.235 -108.635 ;
        RECT -37.565 -110.325 -37.235 -109.995 ;
        RECT -37.565 -113.045 -37.235 -112.715 ;
        RECT -37.565 -114.405 -37.235 -114.075 ;
        RECT -37.565 -115.765 -37.235 -115.435 ;
        RECT -37.565 -117.125 -37.235 -116.795 ;
        RECT -37.565 -118.485 -37.235 -118.155 ;
        RECT -37.565 -119.79 -37.235 -119.46 ;
        RECT -37.565 -121.205 -37.235 -120.875 ;
        RECT -37.565 -122.565 -37.235 -122.235 ;
        RECT -37.565 -123.925 -37.235 -123.595 ;
        RECT -37.565 -126.645 -37.235 -126.315 ;
        RECT -37.565 -128.43 -37.235 -128.1 ;
        RECT -37.565 -129.365 -37.235 -129.035 ;
        RECT -37.565 -130.725 -37.235 -130.395 ;
        RECT -37.565 -133.445 -37.235 -133.115 ;
        RECT -37.565 -134.805 -37.235 -134.475 ;
        RECT -37.565 -136.165 -37.235 -135.835 ;
        RECT -37.565 -137.525 -37.235 -137.195 ;
        RECT -37.565 -140.245 -37.235 -139.915 ;
        RECT -37.565 -142.965 -37.235 -142.635 ;
        RECT -37.565 -144.325 -37.235 -143.995 ;
        RECT -37.565 -145.685 -37.235 -145.355 ;
        RECT -37.565 -147.045 -37.235 -146.715 ;
        RECT -37.565 -148.405 -37.235 -148.075 ;
        RECT -37.565 -149.765 -37.235 -149.435 ;
        RECT -37.565 -151.125 -37.235 -150.795 ;
        RECT -37.565 -152.485 -37.235 -152.155 ;
        RECT -37.565 -153.845 -37.235 -153.515 ;
        RECT -37.565 -155.205 -37.235 -154.875 ;
        RECT -37.565 -156.565 -37.235 -156.235 ;
        RECT -37.565 -157.925 -37.235 -157.595 ;
        RECT -37.565 -159.285 -37.235 -158.955 ;
        RECT -37.565 -160.645 -37.235 -160.315 ;
        RECT -37.565 -162.005 -37.235 -161.675 ;
        RECT -37.565 -163.365 -37.235 -163.035 ;
        RECT -37.565 -164.725 -37.235 -164.395 ;
        RECT -37.565 -166.085 -37.235 -165.755 ;
        RECT -37.565 -167.445 -37.235 -167.115 ;
        RECT -37.565 -168.805 -37.235 -168.475 ;
        RECT -37.565 -170.165 -37.235 -169.835 ;
        RECT -37.565 -171.525 -37.235 -171.195 ;
        RECT -37.565 -172.885 -37.235 -172.555 ;
        RECT -37.565 -174.245 -37.235 -173.915 ;
        RECT -37.565 -175.605 -37.235 -175.275 ;
        RECT -37.565 -176.965 -37.235 -176.635 ;
        RECT -37.565 -178.325 -37.235 -177.995 ;
        RECT -37.565 -179.685 -37.235 -179.355 ;
        RECT -37.565 -181.045 -37.235 -180.715 ;
        RECT -37.565 -182.405 -37.235 -182.075 ;
        RECT -37.565 -183.765 -37.235 -183.435 ;
        RECT -37.565 -185.125 -37.235 -184.795 ;
        RECT -37.565 -186.485 -37.235 -186.155 ;
        RECT -37.565 -187.845 -37.235 -187.515 ;
        RECT -37.565 -189.205 -37.235 -188.875 ;
        RECT -37.565 -190.565 -37.235 -190.235 ;
        RECT -37.565 -191.925 -37.235 -191.595 ;
        RECT -37.565 -193.285 -37.235 -192.955 ;
        RECT -37.565 -194.645 -37.235 -194.315 ;
        RECT -37.565 -196.005 -37.235 -195.675 ;
        RECT -37.565 -197.365 -37.235 -197.035 ;
        RECT -37.565 -198.725 -37.235 -198.395 ;
        RECT -37.565 -200.085 -37.235 -199.755 ;
        RECT -37.565 -201.445 -37.235 -201.115 ;
        RECT -37.565 -202.805 -37.235 -202.475 ;
        RECT -37.565 -204.165 -37.235 -203.835 ;
        RECT -37.565 -205.525 -37.235 -205.195 ;
        RECT -37.565 -208.245 -37.235 -207.915 ;
        RECT -37.565 -210.965 -37.235 -210.635 ;
        RECT -37.565 -212.325 -37.235 -211.995 ;
        RECT -37.565 -213.625 -37.235 -213.295 ;
        RECT -37.565 -215.045 -37.235 -214.715 ;
        RECT -37.565 -216.405 -37.235 -216.075 ;
        RECT -37.565 -217.765 -37.235 -217.435 ;
        RECT -37.565 -219.125 -37.235 -218.795 ;
        RECT -37.565 -221.37 -37.235 -220.24 ;
        RECT -37.56 -221.485 -37.24 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.205 129.8 -35.875 130.93 ;
        RECT -36.205 127.675 -35.875 128.005 ;
        RECT -36.205 126.315 -35.875 126.645 ;
        RECT -36.205 124.955 -35.875 125.285 ;
        RECT -36.205 123.595 -35.875 123.925 ;
        RECT -36.205 122.235 -35.875 122.565 ;
        RECT -36.205 120.875 -35.875 121.205 ;
        RECT -36.205 119.515 -35.875 119.845 ;
        RECT -36.205 118.155 -35.875 118.485 ;
        RECT -36.205 116.795 -35.875 117.125 ;
        RECT -36.205 115.435 -35.875 115.765 ;
        RECT -36.205 114.075 -35.875 114.405 ;
        RECT -36.205 112.715 -35.875 113.045 ;
        RECT -36.205 111.355 -35.875 111.685 ;
        RECT -36.205 109.995 -35.875 110.325 ;
        RECT -36.205 108.635 -35.875 108.965 ;
        RECT -36.205 107.275 -35.875 107.605 ;
        RECT -36.205 105.915 -35.875 106.245 ;
        RECT -36.205 104.555 -35.875 104.885 ;
        RECT -36.205 103.195 -35.875 103.525 ;
        RECT -36.205 101.835 -35.875 102.165 ;
        RECT -36.205 100.475 -35.875 100.805 ;
        RECT -36.205 99.115 -35.875 99.445 ;
        RECT -36.205 97.755 -35.875 98.085 ;
        RECT -36.205 96.395 -35.875 96.725 ;
        RECT -36.205 95.035 -35.875 95.365 ;
        RECT -36.205 93.675 -35.875 94.005 ;
        RECT -36.205 92.315 -35.875 92.645 ;
        RECT -36.205 90.955 -35.875 91.285 ;
        RECT -36.205 89.595 -35.875 89.925 ;
        RECT -36.205 88.235 -35.875 88.565 ;
        RECT -36.205 86.875 -35.875 87.205 ;
        RECT -36.205 85.515 -35.875 85.845 ;
        RECT -36.205 84.155 -35.875 84.485 ;
        RECT -36.205 82.795 -35.875 83.125 ;
        RECT -36.205 81.435 -35.875 81.765 ;
        RECT -36.205 80.075 -35.875 80.405 ;
        RECT -36.205 78.715 -35.875 79.045 ;
        RECT -36.205 77.355 -35.875 77.685 ;
        RECT -36.205 75.995 -35.875 76.325 ;
        RECT -36.205 74.635 -35.875 74.965 ;
        RECT -36.205 73.275 -35.875 73.605 ;
        RECT -36.205 71.915 -35.875 72.245 ;
        RECT -36.205 70.555 -35.875 70.885 ;
        RECT -36.205 69.195 -35.875 69.525 ;
        RECT -36.205 67.835 -35.875 68.165 ;
        RECT -36.205 66.475 -35.875 66.805 ;
        RECT -36.205 65.115 -35.875 65.445 ;
        RECT -36.205 63.755 -35.875 64.085 ;
        RECT -36.205 62.395 -35.875 62.725 ;
        RECT -36.205 61.035 -35.875 61.365 ;
        RECT -36.205 59.675 -35.875 60.005 ;
        RECT -36.205 58.315 -35.875 58.645 ;
        RECT -36.205 56.955 -35.875 57.285 ;
        RECT -36.205 55.595 -35.875 55.925 ;
        RECT -36.205 54.235 -35.875 54.565 ;
        RECT -36.205 52.875 -35.875 53.205 ;
        RECT -36.205 51.515 -35.875 51.845 ;
        RECT -36.205 50.155 -35.875 50.485 ;
        RECT -36.205 48.795 -35.875 49.125 ;
        RECT -36.205 47.435 -35.875 47.765 ;
        RECT -36.205 46.075 -35.875 46.405 ;
        RECT -36.205 44.715 -35.875 45.045 ;
        RECT -36.205 43.355 -35.875 43.685 ;
        RECT -36.205 41.995 -35.875 42.325 ;
        RECT -36.205 40.635 -35.875 40.965 ;
        RECT -36.205 39.275 -35.875 39.605 ;
        RECT -36.205 37.915 -35.875 38.245 ;
        RECT -36.205 36.555 -35.875 36.885 ;
        RECT -36.205 35.195 -35.875 35.525 ;
        RECT -36.205 33.835 -35.875 34.165 ;
        RECT -36.205 32.475 -35.875 32.805 ;
        RECT -36.205 31.115 -35.875 31.445 ;
        RECT -36.205 29.755 -35.875 30.085 ;
        RECT -36.205 28.395 -35.875 28.725 ;
        RECT -36.205 27.035 -35.875 27.365 ;
        RECT -36.205 25.675 -35.875 26.005 ;
        RECT -36.205 24.315 -35.875 24.645 ;
        RECT -36.205 22.955 -35.875 23.285 ;
        RECT -36.205 21.595 -35.875 21.925 ;
        RECT -36.205 20.235 -35.875 20.565 ;
        RECT -36.205 18.875 -35.875 19.205 ;
        RECT -36.205 17.515 -35.875 17.845 ;
        RECT -36.205 16.155 -35.875 16.485 ;
        RECT -36.205 14.795 -35.875 15.125 ;
        RECT -36.205 13.435 -35.875 13.765 ;
        RECT -36.205 12.075 -35.875 12.405 ;
        RECT -36.205 10.715 -35.875 11.045 ;
        RECT -36.205 9.355 -35.875 9.685 ;
        RECT -36.205 7.995 -35.875 8.325 ;
        RECT -36.205 6.635 -35.875 6.965 ;
        RECT -36.205 5.275 -35.875 5.605 ;
        RECT -36.205 3.915 -35.875 4.245 ;
        RECT -36.205 2.555 -35.875 2.885 ;
        RECT -36.205 1.195 -35.875 1.525 ;
        RECT -36.205 -0.165 -35.875 0.165 ;
        RECT -36.205 -1.525 -35.875 -1.195 ;
        RECT -36.205 -2.885 -35.875 -2.555 ;
        RECT -36.205 -6.965 -35.875 -6.635 ;
        RECT -36.205 -8.325 -35.875 -7.995 ;
        RECT -36.205 -9.685 -35.875 -9.355 ;
        RECT -36.205 -11.045 -35.875 -10.715 ;
        RECT -36.205 -12.405 -35.875 -12.075 ;
        RECT -36.205 -13.765 -35.875 -13.435 ;
        RECT -36.205 -15.125 -35.875 -14.795 ;
        RECT -36.205 -16.485 -35.875 -16.155 ;
        RECT -36.205 -17.845 -35.875 -17.515 ;
        RECT -36.205 -19.205 -35.875 -18.875 ;
        RECT -36.205 -20.565 -35.875 -20.235 ;
        RECT -36.205 -27.365 -35.875 -27.035 ;
        RECT -36.205 -28.725 -35.875 -28.395 ;
        RECT -36.205 -30.085 -35.875 -29.755 ;
        RECT -36.205 -32.805 -35.875 -32.475 ;
        RECT -36.205 -35.525 -35.875 -35.195 ;
        RECT -36.205 -36.885 -35.875 -36.555 ;
        RECT -36.205 -39.605 -35.875 -39.275 ;
        RECT -36.205 -40.965 -35.875 -40.635 ;
        RECT -36.205 -42.325 -35.875 -41.995 ;
        RECT -36.205 -43.685 -35.875 -43.355 ;
        RECT -36.205 -45.045 -35.875 -44.715 ;
        RECT -36.205 -46.405 -35.875 -46.075 ;
        RECT -36.205 -47.765 -35.875 -47.435 ;
        RECT -36.205 -49.125 -35.875 -48.795 ;
        RECT -36.205 -50.485 -35.875 -50.155 ;
        RECT -36.205 -51.845 -35.875 -51.515 ;
        RECT -36.205 -53.205 -35.875 -52.875 ;
        RECT -36.205 -54.565 -35.875 -54.235 ;
        RECT -36.205 -55.925 -35.875 -55.595 ;
        RECT -36.205 -57.285 -35.875 -56.955 ;
        RECT -36.205 -58.645 -35.875 -58.315 ;
        RECT -36.205 -60.005 -35.875 -59.675 ;
        RECT -36.205 -61.365 -35.875 -61.035 ;
        RECT -36.205 -62.725 -35.875 -62.395 ;
        RECT -36.205 -64.085 -35.875 -63.755 ;
        RECT -36.205 -65.445 -35.875 -65.115 ;
        RECT -36.205 -66.805 -35.875 -66.475 ;
        RECT -36.205 -68.165 -35.875 -67.835 ;
        RECT -36.205 -69.525 -35.875 -69.195 ;
        RECT -36.205 -70.885 -35.875 -70.555 ;
        RECT -36.205 -72.245 -35.875 -71.915 ;
        RECT -36.205 -73.605 -35.875 -73.275 ;
        RECT -36.205 -74.965 -35.875 -74.635 ;
        RECT -36.205 -76.325 -35.875 -75.995 ;
        RECT -36.205 -77.685 -35.875 -77.355 ;
        RECT -36.205 -79.045 -35.875 -78.715 ;
        RECT -36.205 -80.405 -35.875 -80.075 ;
        RECT -36.205 -81.765 -35.875 -81.435 ;
        RECT -36.205 -83.125 -35.875 -82.795 ;
        RECT -36.205 -84.485 -35.875 -84.155 ;
        RECT -36.205 -85.845 -35.875 -85.515 ;
        RECT -36.205 -87.205 -35.875 -86.875 ;
        RECT -36.205 -88.565 -35.875 -88.235 ;
        RECT -36.205 -89.925 -35.875 -89.595 ;
        RECT -36.205 -91.285 -35.875 -90.955 ;
        RECT -36.205 -92.645 -35.875 -92.315 ;
        RECT -36.205 -94.005 -35.875 -93.675 ;
        RECT -36.205 -95.365 -35.875 -95.035 ;
        RECT -36.205 -96.725 -35.875 -96.395 ;
        RECT -36.205 -98.085 -35.875 -97.755 ;
        RECT -36.205 -99.445 -35.875 -99.115 ;
        RECT -36.205 -100.805 -35.875 -100.475 ;
        RECT -36.205 -102.165 -35.875 -101.835 ;
        RECT -36.205 -103.525 -35.875 -103.195 ;
        RECT -36.205 -104.885 -35.875 -104.555 ;
        RECT -36.205 -106.245 -35.875 -105.915 ;
        RECT -36.205 -108.965 -35.875 -108.635 ;
        RECT -36.205 -110.325 -35.875 -109.995 ;
        RECT -36.205 -113.045 -35.875 -112.715 ;
        RECT -36.205 -114.405 -35.875 -114.075 ;
        RECT -36.205 -115.765 -35.875 -115.435 ;
        RECT -36.205 -117.125 -35.875 -116.795 ;
        RECT -36.205 -118.485 -35.875 -118.155 ;
        RECT -36.205 -119.79 -35.875 -119.46 ;
        RECT -36.205 -121.205 -35.875 -120.875 ;
        RECT -36.205 -122.565 -35.875 -122.235 ;
        RECT -36.205 -123.925 -35.875 -123.595 ;
        RECT -36.205 -126.645 -35.875 -126.315 ;
        RECT -36.205 -128.43 -35.875 -128.1 ;
        RECT -36.205 -129.365 -35.875 -129.035 ;
        RECT -36.205 -130.725 -35.875 -130.395 ;
        RECT -36.205 -133.445 -35.875 -133.115 ;
        RECT -36.205 -134.805 -35.875 -134.475 ;
        RECT -36.205 -136.165 -35.875 -135.835 ;
        RECT -36.205 -137.525 -35.875 -137.195 ;
        RECT -36.205 -140.245 -35.875 -139.915 ;
        RECT -36.205 -142.965 -35.875 -142.635 ;
        RECT -36.205 -144.325 -35.875 -143.995 ;
        RECT -36.205 -145.685 -35.875 -145.355 ;
        RECT -36.205 -147.045 -35.875 -146.715 ;
        RECT -36.205 -148.405 -35.875 -148.075 ;
        RECT -36.205 -149.765 -35.875 -149.435 ;
        RECT -36.205 -151.125 -35.875 -150.795 ;
        RECT -36.205 -152.485 -35.875 -152.155 ;
        RECT -36.205 -153.845 -35.875 -153.515 ;
        RECT -36.205 -155.205 -35.875 -154.875 ;
        RECT -36.205 -156.565 -35.875 -156.235 ;
        RECT -36.205 -157.925 -35.875 -157.595 ;
        RECT -36.205 -159.285 -35.875 -158.955 ;
        RECT -36.205 -160.645 -35.875 -160.315 ;
        RECT -36.205 -162.005 -35.875 -161.675 ;
        RECT -36.205 -163.365 -35.875 -163.035 ;
        RECT -36.205 -164.725 -35.875 -164.395 ;
        RECT -36.205 -166.085 -35.875 -165.755 ;
        RECT -36.205 -167.445 -35.875 -167.115 ;
        RECT -36.205 -168.805 -35.875 -168.475 ;
        RECT -36.205 -170.165 -35.875 -169.835 ;
        RECT -36.205 -171.525 -35.875 -171.195 ;
        RECT -36.205 -172.885 -35.875 -172.555 ;
        RECT -36.205 -174.245 -35.875 -173.915 ;
        RECT -36.205 -175.605 -35.875 -175.275 ;
        RECT -36.205 -176.965 -35.875 -176.635 ;
        RECT -36.205 -178.325 -35.875 -177.995 ;
        RECT -36.205 -179.685 -35.875 -179.355 ;
        RECT -36.205 -181.045 -35.875 -180.715 ;
        RECT -36.205 -182.405 -35.875 -182.075 ;
        RECT -36.205 -183.765 -35.875 -183.435 ;
        RECT -36.205 -185.125 -35.875 -184.795 ;
        RECT -36.205 -186.485 -35.875 -186.155 ;
        RECT -36.205 -187.845 -35.875 -187.515 ;
        RECT -36.205 -189.205 -35.875 -188.875 ;
        RECT -36.205 -190.565 -35.875 -190.235 ;
        RECT -36.205 -191.925 -35.875 -191.595 ;
        RECT -36.205 -193.285 -35.875 -192.955 ;
        RECT -36.205 -194.645 -35.875 -194.315 ;
        RECT -36.205 -196.005 -35.875 -195.675 ;
        RECT -36.205 -197.365 -35.875 -197.035 ;
        RECT -36.205 -198.725 -35.875 -198.395 ;
        RECT -36.205 -200.085 -35.875 -199.755 ;
        RECT -36.205 -201.445 -35.875 -201.115 ;
        RECT -36.205 -202.805 -35.875 -202.475 ;
        RECT -36.205 -204.165 -35.875 -203.835 ;
        RECT -36.205 -205.525 -35.875 -205.195 ;
        RECT -36.205 -208.245 -35.875 -207.915 ;
        RECT -36.205 -212.325 -35.875 -211.995 ;
        RECT -36.205 -213.625 -35.875 -213.295 ;
        RECT -36.205 -215.045 -35.875 -214.715 ;
        RECT -36.205 -216.405 -35.875 -216.075 ;
        RECT -36.205 -217.765 -35.875 -217.435 ;
        RECT -36.205 -219.125 -35.875 -218.795 ;
        RECT -36.205 -221.37 -35.875 -220.24 ;
        RECT -36.2 -221.485 -35.88 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -34.845 48.795 -34.515 49.125 ;
        RECT -34.845 47.435 -34.515 47.765 ;
        RECT -34.845 46.075 -34.515 46.405 ;
        RECT -34.845 44.715 -34.515 45.045 ;
        RECT -34.845 43.355 -34.515 43.685 ;
        RECT -34.845 41.995 -34.515 42.325 ;
        RECT -34.845 40.635 -34.515 40.965 ;
        RECT -34.845 39.275 -34.515 39.605 ;
        RECT -34.845 37.915 -34.515 38.245 ;
        RECT -34.845 36.555 -34.515 36.885 ;
        RECT -34.845 35.195 -34.515 35.525 ;
        RECT -34.845 33.835 -34.515 34.165 ;
        RECT -34.845 32.475 -34.515 32.805 ;
        RECT -34.845 31.115 -34.515 31.445 ;
        RECT -34.845 29.755 -34.515 30.085 ;
        RECT -34.845 28.395 -34.515 28.725 ;
        RECT -34.845 27.035 -34.515 27.365 ;
        RECT -34.845 25.675 -34.515 26.005 ;
        RECT -34.845 24.315 -34.515 24.645 ;
        RECT -34.845 22.955 -34.515 23.285 ;
        RECT -34.845 21.595 -34.515 21.925 ;
        RECT -34.845 20.235 -34.515 20.565 ;
        RECT -34.845 18.875 -34.515 19.205 ;
        RECT -34.845 17.515 -34.515 17.845 ;
        RECT -34.845 16.155 -34.515 16.485 ;
        RECT -34.845 14.795 -34.515 15.125 ;
        RECT -34.845 13.435 -34.515 13.765 ;
        RECT -34.845 12.075 -34.515 12.405 ;
        RECT -34.845 10.715 -34.515 11.045 ;
        RECT -34.845 9.355 -34.515 9.685 ;
        RECT -34.845 7.995 -34.515 8.325 ;
        RECT -34.845 6.635 -34.515 6.965 ;
        RECT -34.845 5.275 -34.515 5.605 ;
        RECT -34.845 3.915 -34.515 4.245 ;
        RECT -34.845 2.555 -34.515 2.885 ;
        RECT -34.845 1.195 -34.515 1.525 ;
        RECT -34.845 -0.165 -34.515 0.165 ;
        RECT -34.845 -1.525 -34.515 -1.195 ;
        RECT -34.845 -6.965 -34.515 -6.635 ;
        RECT -34.845 -8.325 -34.515 -7.995 ;
        RECT -34.845 -9.685 -34.515 -9.355 ;
        RECT -34.845 -11.045 -34.515 -10.715 ;
        RECT -34.845 -12.405 -34.515 -12.075 ;
        RECT -34.845 -13.765 -34.515 -13.435 ;
        RECT -34.845 -15.125 -34.515 -14.795 ;
        RECT -34.845 -16.485 -34.515 -16.155 ;
        RECT -34.845 -17.845 -34.515 -17.515 ;
        RECT -34.845 -19.205 -34.515 -18.875 ;
        RECT -34.845 -20.565 -34.515 -20.235 ;
        RECT -34.845 -27.365 -34.515 -27.035 ;
        RECT -34.845 -28.725 -34.515 -28.395 ;
        RECT -34.845 -30.085 -34.515 -29.755 ;
        RECT -34.845 -32.805 -34.515 -32.475 ;
        RECT -34.845 -35.525 -34.515 -35.195 ;
        RECT -34.845 -36.885 -34.515 -36.555 ;
        RECT -34.845 -39.605 -34.515 -39.275 ;
        RECT -34.845 -40.965 -34.515 -40.635 ;
        RECT -34.845 -42.325 -34.515 -41.995 ;
        RECT -34.845 -43.685 -34.515 -43.355 ;
        RECT -34.845 -45.045 -34.515 -44.715 ;
        RECT -34.845 -46.405 -34.515 -46.075 ;
        RECT -34.845 -47.765 -34.515 -47.435 ;
        RECT -34.845 -49.125 -34.515 -48.795 ;
        RECT -34.845 -50.485 -34.515 -50.155 ;
        RECT -34.845 -51.845 -34.515 -51.515 ;
        RECT -34.845 -53.205 -34.515 -52.875 ;
        RECT -34.845 -54.565 -34.515 -54.235 ;
        RECT -34.845 -55.925 -34.515 -55.595 ;
        RECT -34.845 -57.285 -34.515 -56.955 ;
        RECT -34.845 -58.645 -34.515 -58.315 ;
        RECT -34.845 -60.005 -34.515 -59.675 ;
        RECT -34.845 -61.365 -34.515 -61.035 ;
        RECT -34.845 -62.725 -34.515 -62.395 ;
        RECT -34.845 -64.085 -34.515 -63.755 ;
        RECT -34.845 -65.445 -34.515 -65.115 ;
        RECT -34.845 -66.805 -34.515 -66.475 ;
        RECT -34.845 -68.165 -34.515 -67.835 ;
        RECT -34.845 -69.525 -34.515 -69.195 ;
        RECT -34.845 -70.885 -34.515 -70.555 ;
        RECT -34.845 -72.245 -34.515 -71.915 ;
        RECT -34.845 -73.605 -34.515 -73.275 ;
        RECT -34.845 -74.965 -34.515 -74.635 ;
        RECT -34.845 -76.325 -34.515 -75.995 ;
        RECT -34.845 -77.685 -34.515 -77.355 ;
        RECT -34.845 -79.045 -34.515 -78.715 ;
        RECT -34.845 -80.405 -34.515 -80.075 ;
        RECT -34.845 -81.765 -34.515 -81.435 ;
        RECT -34.845 -83.125 -34.515 -82.795 ;
        RECT -34.845 -84.485 -34.515 -84.155 ;
        RECT -34.845 -85.845 -34.515 -85.515 ;
        RECT -34.845 -87.205 -34.515 -86.875 ;
        RECT -34.845 -88.565 -34.515 -88.235 ;
        RECT -34.845 -89.925 -34.515 -89.595 ;
        RECT -34.845 -91.285 -34.515 -90.955 ;
        RECT -34.845 -92.645 -34.515 -92.315 ;
        RECT -34.845 -94.005 -34.515 -93.675 ;
        RECT -34.845 -95.365 -34.515 -95.035 ;
        RECT -34.845 -96.725 -34.515 -96.395 ;
        RECT -34.845 -98.085 -34.515 -97.755 ;
        RECT -34.845 -99.445 -34.515 -99.115 ;
        RECT -34.845 -100.805 -34.515 -100.475 ;
        RECT -34.845 -102.165 -34.515 -101.835 ;
        RECT -34.845 -103.525 -34.515 -103.195 ;
        RECT -34.845 -104.885 -34.515 -104.555 ;
        RECT -34.845 -106.245 -34.515 -105.915 ;
        RECT -34.845 -108.965 -34.515 -108.635 ;
        RECT -34.845 -110.325 -34.515 -109.995 ;
        RECT -34.845 -113.045 -34.515 -112.715 ;
        RECT -34.845 -114.405 -34.515 -114.075 ;
        RECT -34.845 -115.765 -34.515 -115.435 ;
        RECT -34.845 -117.125 -34.515 -116.795 ;
        RECT -34.845 -118.485 -34.515 -118.155 ;
        RECT -34.845 -119.79 -34.515 -119.46 ;
        RECT -34.845 -121.205 -34.515 -120.875 ;
        RECT -34.845 -122.565 -34.515 -122.235 ;
        RECT -34.845 -123.925 -34.515 -123.595 ;
        RECT -34.845 -126.645 -34.515 -126.315 ;
        RECT -34.845 -128.43 -34.515 -128.1 ;
        RECT -34.845 -129.365 -34.515 -129.035 ;
        RECT -34.845 -130.725 -34.515 -130.395 ;
        RECT -34.84 -132.76 -34.52 131.045 ;
        RECT -34.845 129.8 -34.515 130.93 ;
        RECT -34.845 127.675 -34.515 128.005 ;
        RECT -34.845 126.315 -34.515 126.645 ;
        RECT -34.845 124.955 -34.515 125.285 ;
        RECT -34.845 123.595 -34.515 123.925 ;
        RECT -34.845 122.235 -34.515 122.565 ;
        RECT -34.845 120.875 -34.515 121.205 ;
        RECT -34.845 119.515 -34.515 119.845 ;
        RECT -34.845 118.155 -34.515 118.485 ;
        RECT -34.845 116.795 -34.515 117.125 ;
        RECT -34.845 115.435 -34.515 115.765 ;
        RECT -34.845 114.075 -34.515 114.405 ;
        RECT -34.845 112.715 -34.515 113.045 ;
        RECT -34.845 111.355 -34.515 111.685 ;
        RECT -34.845 109.995 -34.515 110.325 ;
        RECT -34.845 108.635 -34.515 108.965 ;
        RECT -34.845 107.275 -34.515 107.605 ;
        RECT -34.845 105.915 -34.515 106.245 ;
        RECT -34.845 104.555 -34.515 104.885 ;
        RECT -34.845 103.195 -34.515 103.525 ;
        RECT -34.845 101.835 -34.515 102.165 ;
        RECT -34.845 100.475 -34.515 100.805 ;
        RECT -34.845 99.115 -34.515 99.445 ;
        RECT -34.845 97.755 -34.515 98.085 ;
        RECT -34.845 96.395 -34.515 96.725 ;
        RECT -34.845 95.035 -34.515 95.365 ;
        RECT -34.845 93.675 -34.515 94.005 ;
        RECT -34.845 92.315 -34.515 92.645 ;
        RECT -34.845 90.955 -34.515 91.285 ;
        RECT -34.845 89.595 -34.515 89.925 ;
        RECT -34.845 88.235 -34.515 88.565 ;
        RECT -34.845 86.875 -34.515 87.205 ;
        RECT -34.845 85.515 -34.515 85.845 ;
        RECT -34.845 84.155 -34.515 84.485 ;
        RECT -34.845 82.795 -34.515 83.125 ;
        RECT -34.845 81.435 -34.515 81.765 ;
        RECT -34.845 80.075 -34.515 80.405 ;
        RECT -34.845 78.715 -34.515 79.045 ;
        RECT -34.845 77.355 -34.515 77.685 ;
        RECT -34.845 75.995 -34.515 76.325 ;
        RECT -34.845 74.635 -34.515 74.965 ;
        RECT -34.845 73.275 -34.515 73.605 ;
        RECT -34.845 71.915 -34.515 72.245 ;
        RECT -34.845 70.555 -34.515 70.885 ;
        RECT -34.845 69.195 -34.515 69.525 ;
        RECT -34.845 67.835 -34.515 68.165 ;
        RECT -34.845 66.475 -34.515 66.805 ;
        RECT -34.845 65.115 -34.515 65.445 ;
        RECT -34.845 63.755 -34.515 64.085 ;
        RECT -34.845 62.395 -34.515 62.725 ;
        RECT -34.845 61.035 -34.515 61.365 ;
        RECT -34.845 59.675 -34.515 60.005 ;
        RECT -34.845 58.315 -34.515 58.645 ;
        RECT -34.845 56.955 -34.515 57.285 ;
        RECT -34.845 55.595 -34.515 55.925 ;
        RECT -34.845 54.235 -34.515 54.565 ;
        RECT -34.845 52.875 -34.515 53.205 ;
        RECT -34.845 51.515 -34.515 51.845 ;
        RECT -34.845 50.155 -34.515 50.485 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.085 -212.325 -46.755 -211.995 ;
        RECT -47.085 -215.045 -46.755 -214.715 ;
        RECT -47.085 -216.405 -46.755 -216.075 ;
        RECT -47.085 -217.765 -46.755 -217.435 ;
        RECT -47.085 -219.125 -46.755 -218.795 ;
        RECT -47.085 -221.37 -46.755 -220.24 ;
        RECT -47.08 -221.485 -46.76 -210.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.725 129.8 -45.395 130.93 ;
        RECT -45.725 127.675 -45.395 128.005 ;
        RECT -45.725 126.315 -45.395 126.645 ;
        RECT -45.725 124.955 -45.395 125.285 ;
        RECT -45.725 123.595 -45.395 123.925 ;
        RECT -45.725 122.235 -45.395 122.565 ;
        RECT -45.725 120.875 -45.395 121.205 ;
        RECT -45.725 119.515 -45.395 119.845 ;
        RECT -45.725 118.155 -45.395 118.485 ;
        RECT -45.725 116.795 -45.395 117.125 ;
        RECT -45.725 115.435 -45.395 115.765 ;
        RECT -45.725 114.075 -45.395 114.405 ;
        RECT -45.725 112.715 -45.395 113.045 ;
        RECT -45.725 111.355 -45.395 111.685 ;
        RECT -45.725 109.995 -45.395 110.325 ;
        RECT -45.725 108.635 -45.395 108.965 ;
        RECT -45.725 107.275 -45.395 107.605 ;
        RECT -45.725 105.915 -45.395 106.245 ;
        RECT -45.725 104.555 -45.395 104.885 ;
        RECT -45.725 103.195 -45.395 103.525 ;
        RECT -45.725 101.835 -45.395 102.165 ;
        RECT -45.725 100.475 -45.395 100.805 ;
        RECT -45.725 99.115 -45.395 99.445 ;
        RECT -45.725 97.755 -45.395 98.085 ;
        RECT -45.725 96.395 -45.395 96.725 ;
        RECT -45.725 95.035 -45.395 95.365 ;
        RECT -45.725 93.675 -45.395 94.005 ;
        RECT -45.725 92.315 -45.395 92.645 ;
        RECT -45.725 90.955 -45.395 91.285 ;
        RECT -45.725 89.595 -45.395 89.925 ;
        RECT -45.725 88.235 -45.395 88.565 ;
        RECT -45.725 86.875 -45.395 87.205 ;
        RECT -45.725 85.515 -45.395 85.845 ;
        RECT -45.725 84.155 -45.395 84.485 ;
        RECT -45.725 82.795 -45.395 83.125 ;
        RECT -45.725 81.435 -45.395 81.765 ;
        RECT -45.725 80.075 -45.395 80.405 ;
        RECT -45.725 78.715 -45.395 79.045 ;
        RECT -45.725 77.355 -45.395 77.685 ;
        RECT -45.725 75.995 -45.395 76.325 ;
        RECT -45.725 74.635 -45.395 74.965 ;
        RECT -45.725 73.275 -45.395 73.605 ;
        RECT -45.72 73.275 -45.4 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.725 48.795 -45.395 49.125 ;
        RECT -45.725 47.435 -45.395 47.765 ;
        RECT -45.725 46.075 -45.395 46.405 ;
        RECT -45.725 44.715 -45.395 45.045 ;
        RECT -45.725 43.355 -45.395 43.685 ;
        RECT -45.725 40.635 -45.395 40.965 ;
        RECT -45.725 39.275 -45.395 39.605 ;
        RECT -45.725 35.195 -45.395 35.525 ;
        RECT -45.725 33.835 -45.395 34.165 ;
        RECT -45.725 32.475 -45.395 32.805 ;
        RECT -45.725 31.115 -45.395 31.445 ;
        RECT -45.725 29.755 -45.395 30.085 ;
        RECT -45.725 28.395 -45.395 28.725 ;
        RECT -45.725 27.035 -45.395 27.365 ;
        RECT -45.725 25.675 -45.395 26.005 ;
        RECT -45.725 24.315 -45.395 24.645 ;
        RECT -45.725 22.955 -45.395 23.285 ;
        RECT -45.725 21.595 -45.395 21.925 ;
        RECT -45.725 20.235 -45.395 20.565 ;
        RECT -45.725 18.875 -45.395 19.205 ;
        RECT -45.725 17.515 -45.395 17.845 ;
        RECT -45.725 16.155 -45.395 16.485 ;
        RECT -45.725 14.795 -45.395 15.125 ;
        RECT -45.725 13.435 -45.395 13.765 ;
        RECT -45.725 12.075 -45.395 12.405 ;
        RECT -45.725 10.715 -45.395 11.045 ;
        RECT -45.725 9.355 -45.395 9.685 ;
        RECT -45.725 7.995 -45.395 8.325 ;
        RECT -45.725 6.635 -45.395 6.965 ;
        RECT -45.725 5.275 -45.395 5.605 ;
        RECT -45.725 3.915 -45.395 4.245 ;
        RECT -45.725 2.555 -45.395 2.885 ;
        RECT -45.725 1.195 -45.395 1.525 ;
        RECT -45.725 -0.165 -45.395 0.165 ;
        RECT -45.725 -1.525 -45.395 -1.195 ;
        RECT -45.725 -2.885 -45.395 -2.555 ;
        RECT -45.725 -4.245 -45.395 -3.915 ;
        RECT -45.725 -5.605 -45.395 -5.275 ;
        RECT -45.725 -6.965 -45.395 -6.635 ;
        RECT -45.725 -8.325 -45.395 -7.995 ;
        RECT -45.725 -9.685 -45.395 -9.355 ;
        RECT -45.725 -11.045 -45.395 -10.715 ;
        RECT -45.725 -12.405 -45.395 -12.075 ;
        RECT -45.725 -13.765 -45.395 -13.435 ;
        RECT -45.725 -15.125 -45.395 -14.795 ;
        RECT -45.725 -16.485 -45.395 -16.155 ;
        RECT -45.725 -17.845 -45.395 -17.515 ;
        RECT -45.725 -19.205 -45.395 -18.875 ;
        RECT -45.725 -20.565 -45.395 -20.235 ;
        RECT -45.725 -21.925 -45.395 -21.595 ;
        RECT -45.725 -23.285 -45.395 -22.955 ;
        RECT -45.725 -24.645 -45.395 -24.315 ;
        RECT -45.725 -26.005 -45.395 -25.675 ;
        RECT -45.725 -27.365 -45.395 -27.035 ;
        RECT -45.725 -28.725 -45.395 -28.395 ;
        RECT -45.725 -30.085 -45.395 -29.755 ;
        RECT -45.725 -31.445 -45.395 -31.115 ;
        RECT -45.725 -32.805 -45.395 -32.475 ;
        RECT -45.725 -35.525 -45.395 -35.195 ;
        RECT -45.725 -36.885 -45.395 -36.555 ;
        RECT -45.725 -39.605 -45.395 -39.275 ;
        RECT -45.725 -40.965 -45.395 -40.635 ;
        RECT -45.725 -42.325 -45.395 -41.995 ;
        RECT -45.725 -43.685 -45.395 -43.355 ;
        RECT -45.725 -45.045 -45.395 -44.715 ;
        RECT -45.725 -46.405 -45.395 -46.075 ;
        RECT -45.725 -47.765 -45.395 -47.435 ;
        RECT -45.725 -49.125 -45.395 -48.795 ;
        RECT -45.725 -50.485 -45.395 -50.155 ;
        RECT -45.725 -51.845 -45.395 -51.515 ;
        RECT -45.725 -53.205 -45.395 -52.875 ;
        RECT -45.725 -54.565 -45.395 -54.235 ;
        RECT -45.725 -55.925 -45.395 -55.595 ;
        RECT -45.725 -57.285 -45.395 -56.955 ;
        RECT -45.725 -58.645 -45.395 -58.315 ;
        RECT -45.725 -60.005 -45.395 -59.675 ;
        RECT -45.725 -61.365 -45.395 -61.035 ;
        RECT -45.725 -62.725 -45.395 -62.395 ;
        RECT -45.725 -64.085 -45.395 -63.755 ;
        RECT -45.725 -65.445 -45.395 -65.115 ;
        RECT -45.725 -66.805 -45.395 -66.475 ;
        RECT -45.725 -68.165 -45.395 -67.835 ;
        RECT -45.725 -69.525 -45.395 -69.195 ;
        RECT -45.725 -70.885 -45.395 -70.555 ;
        RECT -45.725 -72.245 -45.395 -71.915 ;
        RECT -45.725 -73.605 -45.395 -73.275 ;
        RECT -45.725 -74.965 -45.395 -74.635 ;
        RECT -45.725 -76.325 -45.395 -75.995 ;
        RECT -45.725 -77.685 -45.395 -77.355 ;
        RECT -45.725 -79.045 -45.395 -78.715 ;
        RECT -45.725 -80.405 -45.395 -80.075 ;
        RECT -45.725 -81.765 -45.395 -81.435 ;
        RECT -45.725 -83.125 -45.395 -82.795 ;
        RECT -45.725 -84.485 -45.395 -84.155 ;
        RECT -45.725 -85.845 -45.395 -85.515 ;
        RECT -45.725 -87.205 -45.395 -86.875 ;
        RECT -45.725 -88.565 -45.395 -88.235 ;
        RECT -45.725 -89.925 -45.395 -89.595 ;
        RECT -45.725 -91.285 -45.395 -90.955 ;
        RECT -45.725 -92.645 -45.395 -92.315 ;
        RECT -45.725 -94.005 -45.395 -93.675 ;
        RECT -45.725 -95.365 -45.395 -95.035 ;
        RECT -45.725 -96.725 -45.395 -96.395 ;
        RECT -45.725 -98.085 -45.395 -97.755 ;
        RECT -45.725 -99.445 -45.395 -99.115 ;
        RECT -45.725 -100.805 -45.395 -100.475 ;
        RECT -45.725 -102.165 -45.395 -101.835 ;
        RECT -45.725 -103.525 -45.395 -103.195 ;
        RECT -45.725 -104.885 -45.395 -104.555 ;
        RECT -45.725 -106.245 -45.395 -105.915 ;
        RECT -45.725 -107.605 -45.395 -107.275 ;
        RECT -45.725 -108.965 -45.395 -108.635 ;
        RECT -45.725 -110.325 -45.395 -109.995 ;
        RECT -45.725 -113.045 -45.395 -112.715 ;
        RECT -45.725 -114.405 -45.395 -114.075 ;
        RECT -45.725 -115.765 -45.395 -115.435 ;
        RECT -45.725 -117.125 -45.395 -116.795 ;
        RECT -45.725 -118.485 -45.395 -118.155 ;
        RECT -45.725 -119.79 -45.395 -119.46 ;
        RECT -45.725 -121.205 -45.395 -120.875 ;
        RECT -45.725 -122.565 -45.395 -122.235 ;
        RECT -45.725 -123.925 -45.395 -123.595 ;
        RECT -45.725 -126.645 -45.395 -126.315 ;
        RECT -45.725 -128.43 -45.395 -128.1 ;
        RECT -45.725 -129.365 -45.395 -129.035 ;
        RECT -45.725 -130.725 -45.395 -130.395 ;
        RECT -45.725 -134.805 -45.395 -134.475 ;
        RECT -45.725 -136.165 -45.395 -135.835 ;
        RECT -45.725 -137.525 -45.395 -137.195 ;
        RECT -45.725 -138.885 -45.395 -138.555 ;
        RECT -45.725 -140.245 -45.395 -139.915 ;
        RECT -45.725 -142.965 -45.395 -142.635 ;
        RECT -45.725 -144.325 -45.395 -143.995 ;
        RECT -45.725 -145.685 -45.395 -145.355 ;
        RECT -45.725 -147.045 -45.395 -146.715 ;
        RECT -45.725 -148.405 -45.395 -148.075 ;
        RECT -45.725 -149.765 -45.395 -149.435 ;
        RECT -45.725 -151.125 -45.395 -150.795 ;
        RECT -45.725 -152.485 -45.395 -152.155 ;
        RECT -45.725 -153.845 -45.395 -153.515 ;
        RECT -45.725 -155.205 -45.395 -154.875 ;
        RECT -45.725 -156.565 -45.395 -156.235 ;
        RECT -45.725 -157.925 -45.395 -157.595 ;
        RECT -45.725 -159.285 -45.395 -158.955 ;
        RECT -45.725 -160.645 -45.395 -160.315 ;
        RECT -45.725 -162.005 -45.395 -161.675 ;
        RECT -45.725 -163.365 -45.395 -163.035 ;
        RECT -45.725 -164.725 -45.395 -164.395 ;
        RECT -45.725 -166.085 -45.395 -165.755 ;
        RECT -45.725 -167.445 -45.395 -167.115 ;
        RECT -45.725 -168.805 -45.395 -168.475 ;
        RECT -45.725 -170.165 -45.395 -169.835 ;
        RECT -45.725 -171.525 -45.395 -171.195 ;
        RECT -45.725 -172.885 -45.395 -172.555 ;
        RECT -45.725 -174.245 -45.395 -173.915 ;
        RECT -45.725 -175.605 -45.395 -175.275 ;
        RECT -45.725 -176.965 -45.395 -176.635 ;
        RECT -45.725 -178.325 -45.395 -177.995 ;
        RECT -45.725 -179.685 -45.395 -179.355 ;
        RECT -45.725 -181.045 -45.395 -180.715 ;
        RECT -45.725 -182.405 -45.395 -182.075 ;
        RECT -45.725 -183.765 -45.395 -183.435 ;
        RECT -45.725 -185.125 -45.395 -184.795 ;
        RECT -45.725 -186.485 -45.395 -186.155 ;
        RECT -45.725 -187.845 -45.395 -187.515 ;
        RECT -45.725 -189.205 -45.395 -188.875 ;
        RECT -45.725 -190.565 -45.395 -190.235 ;
        RECT -45.725 -191.925 -45.395 -191.595 ;
        RECT -45.725 -193.285 -45.395 -192.955 ;
        RECT -45.725 -194.645 -45.395 -194.315 ;
        RECT -45.725 -196.005 -45.395 -195.675 ;
        RECT -45.725 -197.365 -45.395 -197.035 ;
        RECT -45.725 -198.725 -45.395 -198.395 ;
        RECT -45.725 -200.085 -45.395 -199.755 ;
        RECT -45.725 -201.445 -45.395 -201.115 ;
        RECT -45.725 -202.805 -45.395 -202.475 ;
        RECT -45.725 -204.165 -45.395 -203.835 ;
        RECT -45.725 -205.525 -45.395 -205.195 ;
        RECT -45.725 -208.245 -45.395 -207.915 ;
        RECT -45.725 -212.325 -45.395 -211.995 ;
        RECT -45.725 -213.625 -45.395 -213.295 ;
        RECT -45.725 -215.045 -45.395 -214.715 ;
        RECT -45.725 -216.405 -45.395 -216.075 ;
        RECT -45.725 -217.765 -45.395 -217.435 ;
        RECT -45.725 -219.125 -45.395 -218.795 ;
        RECT -45.725 -221.37 -45.395 -220.24 ;
        RECT -45.72 -221.485 -45.4 49.125 ;
    END
    PORT
      LAYER met3 ;
        RECT -44.365 129.8 -44.035 130.93 ;
        RECT -44.365 127.675 -44.035 128.005 ;
        RECT -44.365 126.315 -44.035 126.645 ;
        RECT -44.365 124.955 -44.035 125.285 ;
        RECT -44.365 123.595 -44.035 123.925 ;
        RECT -44.365 122.235 -44.035 122.565 ;
        RECT -44.365 120.875 -44.035 121.205 ;
        RECT -44.365 119.515 -44.035 119.845 ;
        RECT -44.365 118.155 -44.035 118.485 ;
        RECT -44.365 116.795 -44.035 117.125 ;
        RECT -44.365 115.435 -44.035 115.765 ;
        RECT -44.365 114.075 -44.035 114.405 ;
        RECT -44.365 112.715 -44.035 113.045 ;
        RECT -44.365 111.355 -44.035 111.685 ;
        RECT -44.365 109.995 -44.035 110.325 ;
        RECT -44.365 108.635 -44.035 108.965 ;
        RECT -44.365 107.275 -44.035 107.605 ;
        RECT -44.365 105.915 -44.035 106.245 ;
        RECT -44.365 104.555 -44.035 104.885 ;
        RECT -44.365 103.195 -44.035 103.525 ;
        RECT -44.365 101.835 -44.035 102.165 ;
        RECT -44.365 100.475 -44.035 100.805 ;
        RECT -44.365 99.115 -44.035 99.445 ;
        RECT -44.365 97.755 -44.035 98.085 ;
        RECT -44.365 96.395 -44.035 96.725 ;
        RECT -44.365 95.035 -44.035 95.365 ;
        RECT -44.365 93.675 -44.035 94.005 ;
        RECT -44.365 92.315 -44.035 92.645 ;
        RECT -44.365 90.955 -44.035 91.285 ;
        RECT -44.365 89.595 -44.035 89.925 ;
        RECT -44.365 88.235 -44.035 88.565 ;
        RECT -44.365 86.875 -44.035 87.205 ;
        RECT -44.365 85.515 -44.035 85.845 ;
        RECT -44.365 84.155 -44.035 84.485 ;
        RECT -44.365 82.795 -44.035 83.125 ;
        RECT -44.365 81.435 -44.035 81.765 ;
        RECT -44.365 80.075 -44.035 80.405 ;
        RECT -44.365 78.715 -44.035 79.045 ;
        RECT -44.365 77.355 -44.035 77.685 ;
        RECT -44.365 75.995 -44.035 76.325 ;
        RECT -44.365 74.635 -44.035 74.965 ;
        RECT -44.365 73.275 -44.035 73.605 ;
        RECT -44.365 72.445 -44.035 72.775 ;
        RECT -44.365 70.395 -44.035 70.725 ;
        RECT -44.365 68.035 -44.035 68.365 ;
        RECT -44.365 66.885 -44.035 67.215 ;
        RECT -44.365 64.875 -44.035 65.205 ;
        RECT -44.365 63.725 -44.035 64.055 ;
        RECT -44.365 61.715 -44.035 62.045 ;
        RECT -44.365 60.395 -44.035 60.725 ;
        RECT -44.365 58.555 -44.035 58.885 ;
        RECT -44.365 57.405 -44.035 57.735 ;
        RECT -44.365 55.395 -44.035 55.725 ;
        RECT -44.365 54.245 -44.035 54.575 ;
        RECT -44.365 51.885 -44.035 52.215 ;
        RECT -44.365 49.83 -44.035 50.16 ;
        RECT -44.365 48.795 -44.035 49.125 ;
        RECT -44.365 47.435 -44.035 47.765 ;
        RECT -44.365 46.075 -44.035 46.405 ;
        RECT -44.365 44.715 -44.035 45.045 ;
        RECT -44.365 43.355 -44.035 43.685 ;
        RECT -44.365 41.995 -44.035 42.325 ;
        RECT -44.365 40.635 -44.035 40.965 ;
        RECT -44.365 39.275 -44.035 39.605 ;
        RECT -44.365 37.915 -44.035 38.245 ;
        RECT -44.365 36.555 -44.035 36.885 ;
        RECT -44.365 35.195 -44.035 35.525 ;
        RECT -44.365 33.835 -44.035 34.165 ;
        RECT -44.365 32.475 -44.035 32.805 ;
        RECT -44.365 31.115 -44.035 31.445 ;
        RECT -44.365 29.755 -44.035 30.085 ;
        RECT -44.365 28.395 -44.035 28.725 ;
        RECT -44.365 27.035 -44.035 27.365 ;
        RECT -44.365 25.675 -44.035 26.005 ;
        RECT -44.365 24.315 -44.035 24.645 ;
        RECT -44.365 22.955 -44.035 23.285 ;
        RECT -44.365 21.595 -44.035 21.925 ;
        RECT -44.365 20.235 -44.035 20.565 ;
        RECT -44.365 18.875 -44.035 19.205 ;
        RECT -44.365 17.515 -44.035 17.845 ;
        RECT -44.365 16.155 -44.035 16.485 ;
        RECT -44.365 14.795 -44.035 15.125 ;
        RECT -44.365 13.435 -44.035 13.765 ;
        RECT -44.365 12.075 -44.035 12.405 ;
        RECT -44.365 10.715 -44.035 11.045 ;
        RECT -44.365 9.355 -44.035 9.685 ;
        RECT -44.365 7.995 -44.035 8.325 ;
        RECT -44.365 6.635 -44.035 6.965 ;
        RECT -44.365 5.275 -44.035 5.605 ;
        RECT -44.365 3.915 -44.035 4.245 ;
        RECT -44.365 2.555 -44.035 2.885 ;
        RECT -44.365 1.195 -44.035 1.525 ;
        RECT -44.365 -0.165 -44.035 0.165 ;
        RECT -44.365 -1.525 -44.035 -1.195 ;
        RECT -44.365 -2.885 -44.035 -2.555 ;
        RECT -44.365 -4.245 -44.035 -3.915 ;
        RECT -44.365 -5.605 -44.035 -5.275 ;
        RECT -44.365 -6.965 -44.035 -6.635 ;
        RECT -44.365 -8.325 -44.035 -7.995 ;
        RECT -44.365 -9.685 -44.035 -9.355 ;
        RECT -44.365 -11.045 -44.035 -10.715 ;
        RECT -44.365 -12.405 -44.035 -12.075 ;
        RECT -44.365 -13.765 -44.035 -13.435 ;
        RECT -44.365 -15.125 -44.035 -14.795 ;
        RECT -44.365 -16.485 -44.035 -16.155 ;
        RECT -44.365 -17.845 -44.035 -17.515 ;
        RECT -44.365 -19.205 -44.035 -18.875 ;
        RECT -44.365 -20.565 -44.035 -20.235 ;
        RECT -44.365 -21.925 -44.035 -21.595 ;
        RECT -44.365 -23.285 -44.035 -22.955 ;
        RECT -44.365 -24.645 -44.035 -24.315 ;
        RECT -44.365 -26.005 -44.035 -25.675 ;
        RECT -44.365 -27.365 -44.035 -27.035 ;
        RECT -44.365 -28.725 -44.035 -28.395 ;
        RECT -44.365 -30.085 -44.035 -29.755 ;
        RECT -44.365 -32.805 -44.035 -32.475 ;
        RECT -44.365 -35.525 -44.035 -35.195 ;
        RECT -44.365 -36.885 -44.035 -36.555 ;
        RECT -44.365 -39.605 -44.035 -39.275 ;
        RECT -44.365 -40.965 -44.035 -40.635 ;
        RECT -44.365 -42.325 -44.035 -41.995 ;
        RECT -44.365 -43.685 -44.035 -43.355 ;
        RECT -44.365 -45.045 -44.035 -44.715 ;
        RECT -44.365 -46.405 -44.035 -46.075 ;
        RECT -44.365 -47.765 -44.035 -47.435 ;
        RECT -44.365 -49.125 -44.035 -48.795 ;
        RECT -44.365 -50.485 -44.035 -50.155 ;
        RECT -44.365 -51.845 -44.035 -51.515 ;
        RECT -44.365 -53.205 -44.035 -52.875 ;
        RECT -44.365 -54.565 -44.035 -54.235 ;
        RECT -44.365 -55.925 -44.035 -55.595 ;
        RECT -44.365 -57.285 -44.035 -56.955 ;
        RECT -44.365 -58.645 -44.035 -58.315 ;
        RECT -44.365 -60.005 -44.035 -59.675 ;
        RECT -44.365 -61.365 -44.035 -61.035 ;
        RECT -44.365 -62.725 -44.035 -62.395 ;
        RECT -44.365 -64.085 -44.035 -63.755 ;
        RECT -44.365 -65.445 -44.035 -65.115 ;
        RECT -44.365 -66.805 -44.035 -66.475 ;
        RECT -44.365 -68.165 -44.035 -67.835 ;
        RECT -44.365 -69.525 -44.035 -69.195 ;
        RECT -44.365 -70.885 -44.035 -70.555 ;
        RECT -44.365 -72.245 -44.035 -71.915 ;
        RECT -44.365 -73.605 -44.035 -73.275 ;
        RECT -44.365 -74.965 -44.035 -74.635 ;
        RECT -44.365 -76.325 -44.035 -75.995 ;
        RECT -44.365 -77.685 -44.035 -77.355 ;
        RECT -44.365 -79.045 -44.035 -78.715 ;
        RECT -44.365 -80.405 -44.035 -80.075 ;
        RECT -44.365 -81.765 -44.035 -81.435 ;
        RECT -44.365 -83.125 -44.035 -82.795 ;
        RECT -44.365 -84.485 -44.035 -84.155 ;
        RECT -44.365 -85.845 -44.035 -85.515 ;
        RECT -44.365 -87.205 -44.035 -86.875 ;
        RECT -44.365 -88.565 -44.035 -88.235 ;
        RECT -44.365 -89.925 -44.035 -89.595 ;
        RECT -44.365 -91.285 -44.035 -90.955 ;
        RECT -44.365 -92.645 -44.035 -92.315 ;
        RECT -44.365 -94.005 -44.035 -93.675 ;
        RECT -44.365 -95.365 -44.035 -95.035 ;
        RECT -44.365 -96.725 -44.035 -96.395 ;
        RECT -44.365 -98.085 -44.035 -97.755 ;
        RECT -44.365 -99.445 -44.035 -99.115 ;
        RECT -44.365 -100.805 -44.035 -100.475 ;
        RECT -44.365 -102.165 -44.035 -101.835 ;
        RECT -44.365 -103.525 -44.035 -103.195 ;
        RECT -44.365 -104.885 -44.035 -104.555 ;
        RECT -44.365 -106.245 -44.035 -105.915 ;
        RECT -44.365 -107.605 -44.035 -107.275 ;
        RECT -44.365 -108.965 -44.035 -108.635 ;
        RECT -44.365 -110.325 -44.035 -109.995 ;
        RECT -44.365 -113.045 -44.035 -112.715 ;
        RECT -44.365 -114.405 -44.035 -114.075 ;
        RECT -44.365 -115.765 -44.035 -115.435 ;
        RECT -44.365 -117.125 -44.035 -116.795 ;
        RECT -44.365 -118.485 -44.035 -118.155 ;
        RECT -44.365 -119.79 -44.035 -119.46 ;
        RECT -44.365 -121.205 -44.035 -120.875 ;
        RECT -44.365 -122.565 -44.035 -122.235 ;
        RECT -44.365 -123.925 -44.035 -123.595 ;
        RECT -44.365 -126.645 -44.035 -126.315 ;
        RECT -44.365 -128.43 -44.035 -128.1 ;
        RECT -44.365 -129.365 -44.035 -129.035 ;
        RECT -44.365 -130.725 -44.035 -130.395 ;
        RECT -44.365 -134.805 -44.035 -134.475 ;
        RECT -44.365 -136.165 -44.035 -135.835 ;
        RECT -44.365 -137.525 -44.035 -137.195 ;
        RECT -44.365 -140.245 -44.035 -139.915 ;
        RECT -44.365 -142.965 -44.035 -142.635 ;
        RECT -44.365 -144.325 -44.035 -143.995 ;
        RECT -44.365 -145.685 -44.035 -145.355 ;
        RECT -44.365 -147.045 -44.035 -146.715 ;
        RECT -44.365 -148.405 -44.035 -148.075 ;
        RECT -44.365 -149.765 -44.035 -149.435 ;
        RECT -44.365 -151.125 -44.035 -150.795 ;
        RECT -44.365 -152.485 -44.035 -152.155 ;
        RECT -44.365 -153.845 -44.035 -153.515 ;
        RECT -44.365 -155.205 -44.035 -154.875 ;
        RECT -44.365 -156.565 -44.035 -156.235 ;
        RECT -44.365 -157.925 -44.035 -157.595 ;
        RECT -44.365 -159.285 -44.035 -158.955 ;
        RECT -44.365 -160.645 -44.035 -160.315 ;
        RECT -44.365 -162.005 -44.035 -161.675 ;
        RECT -44.365 -163.365 -44.035 -163.035 ;
        RECT -44.365 -164.725 -44.035 -164.395 ;
        RECT -44.365 -166.085 -44.035 -165.755 ;
        RECT -44.365 -167.445 -44.035 -167.115 ;
        RECT -44.365 -168.805 -44.035 -168.475 ;
        RECT -44.365 -170.165 -44.035 -169.835 ;
        RECT -44.365 -171.525 -44.035 -171.195 ;
        RECT -44.365 -172.885 -44.035 -172.555 ;
        RECT -44.365 -174.245 -44.035 -173.915 ;
        RECT -44.365 -175.605 -44.035 -175.275 ;
        RECT -44.365 -176.965 -44.035 -176.635 ;
        RECT -44.365 -178.325 -44.035 -177.995 ;
        RECT -44.365 -179.685 -44.035 -179.355 ;
        RECT -44.365 -181.045 -44.035 -180.715 ;
        RECT -44.365 -182.405 -44.035 -182.075 ;
        RECT -44.365 -183.765 -44.035 -183.435 ;
        RECT -44.365 -185.125 -44.035 -184.795 ;
        RECT -44.365 -186.485 -44.035 -186.155 ;
        RECT -44.365 -187.845 -44.035 -187.515 ;
        RECT -44.365 -189.205 -44.035 -188.875 ;
        RECT -44.365 -190.565 -44.035 -190.235 ;
        RECT -44.365 -191.925 -44.035 -191.595 ;
        RECT -44.365 -193.285 -44.035 -192.955 ;
        RECT -44.365 -194.645 -44.035 -194.315 ;
        RECT -44.365 -196.005 -44.035 -195.675 ;
        RECT -44.365 -197.365 -44.035 -197.035 ;
        RECT -44.365 -198.725 -44.035 -198.395 ;
        RECT -44.365 -200.085 -44.035 -199.755 ;
        RECT -44.365 -201.445 -44.035 -201.115 ;
        RECT -44.365 -202.805 -44.035 -202.475 ;
        RECT -44.365 -204.165 -44.035 -203.835 ;
        RECT -44.365 -205.525 -44.035 -205.195 ;
        RECT -44.365 -208.245 -44.035 -207.915 ;
        RECT -44.365 -210.965 -44.035 -210.635 ;
        RECT -44.365 -212.325 -44.035 -211.995 ;
        RECT -44.365 -213.625 -44.035 -213.295 ;
        RECT -44.365 -215.045 -44.035 -214.715 ;
        RECT -44.365 -216.405 -44.035 -216.075 ;
        RECT -44.365 -217.765 -44.035 -217.435 ;
        RECT -44.365 -219.125 -44.035 -218.795 ;
        RECT -44.365 -221.37 -44.035 -220.24 ;
        RECT -44.36 -221.485 -44.04 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.005 129.8 -42.675 130.93 ;
        RECT -43.005 127.675 -42.675 128.005 ;
        RECT -43.005 126.315 -42.675 126.645 ;
        RECT -43.005 124.955 -42.675 125.285 ;
        RECT -43.005 123.595 -42.675 123.925 ;
        RECT -43.005 122.235 -42.675 122.565 ;
        RECT -43.005 120.875 -42.675 121.205 ;
        RECT -43.005 119.515 -42.675 119.845 ;
        RECT -43.005 118.155 -42.675 118.485 ;
        RECT -43.005 116.795 -42.675 117.125 ;
        RECT -43.005 115.435 -42.675 115.765 ;
        RECT -43.005 114.075 -42.675 114.405 ;
        RECT -43.005 112.715 -42.675 113.045 ;
        RECT -43.005 111.355 -42.675 111.685 ;
        RECT -43.005 109.995 -42.675 110.325 ;
        RECT -43.005 108.635 -42.675 108.965 ;
        RECT -43.005 107.275 -42.675 107.605 ;
        RECT -43.005 105.915 -42.675 106.245 ;
        RECT -43.005 104.555 -42.675 104.885 ;
        RECT -43.005 103.195 -42.675 103.525 ;
        RECT -43.005 101.835 -42.675 102.165 ;
        RECT -43.005 100.475 -42.675 100.805 ;
        RECT -43.005 99.115 -42.675 99.445 ;
        RECT -43.005 97.755 -42.675 98.085 ;
        RECT -43.005 96.395 -42.675 96.725 ;
        RECT -43.005 95.035 -42.675 95.365 ;
        RECT -43.005 93.675 -42.675 94.005 ;
        RECT -43.005 92.315 -42.675 92.645 ;
        RECT -43.005 90.955 -42.675 91.285 ;
        RECT -43.005 89.595 -42.675 89.925 ;
        RECT -43.005 88.235 -42.675 88.565 ;
        RECT -43.005 86.875 -42.675 87.205 ;
        RECT -43.005 85.515 -42.675 85.845 ;
        RECT -43.005 84.155 -42.675 84.485 ;
        RECT -43.005 82.795 -42.675 83.125 ;
        RECT -43.005 81.435 -42.675 81.765 ;
        RECT -43.005 80.075 -42.675 80.405 ;
        RECT -43.005 78.715 -42.675 79.045 ;
        RECT -43.005 77.355 -42.675 77.685 ;
        RECT -43.005 75.995 -42.675 76.325 ;
        RECT -43.005 74.635 -42.675 74.965 ;
        RECT -43.005 73.275 -42.675 73.605 ;
        RECT -43.005 72.445 -42.675 72.775 ;
        RECT -43.005 70.395 -42.675 70.725 ;
        RECT -43.005 68.035 -42.675 68.365 ;
        RECT -43.005 66.885 -42.675 67.215 ;
        RECT -43.005 64.875 -42.675 65.205 ;
        RECT -43.005 63.725 -42.675 64.055 ;
        RECT -43.005 61.715 -42.675 62.045 ;
        RECT -43.005 60.395 -42.675 60.725 ;
        RECT -43.005 58.555 -42.675 58.885 ;
        RECT -43.005 57.405 -42.675 57.735 ;
        RECT -43.005 55.395 -42.675 55.725 ;
        RECT -43.005 54.245 -42.675 54.575 ;
        RECT -43.005 51.885 -42.675 52.215 ;
        RECT -43.005 49.83 -42.675 50.16 ;
        RECT -43.005 48.795 -42.675 49.125 ;
        RECT -43.005 47.435 -42.675 47.765 ;
        RECT -43.005 46.075 -42.675 46.405 ;
        RECT -43.005 44.715 -42.675 45.045 ;
        RECT -43.005 43.355 -42.675 43.685 ;
        RECT -43.005 41.995 -42.675 42.325 ;
        RECT -43.005 40.635 -42.675 40.965 ;
        RECT -43.005 39.275 -42.675 39.605 ;
        RECT -43.005 37.915 -42.675 38.245 ;
        RECT -43.005 36.555 -42.675 36.885 ;
        RECT -43.005 35.195 -42.675 35.525 ;
        RECT -43.005 33.835 -42.675 34.165 ;
        RECT -43.005 32.475 -42.675 32.805 ;
        RECT -43.005 31.115 -42.675 31.445 ;
        RECT -43.005 29.755 -42.675 30.085 ;
        RECT -43.005 28.395 -42.675 28.725 ;
        RECT -43.005 27.035 -42.675 27.365 ;
        RECT -43.005 25.675 -42.675 26.005 ;
        RECT -43.005 24.315 -42.675 24.645 ;
        RECT -43.005 22.955 -42.675 23.285 ;
        RECT -43.005 21.595 -42.675 21.925 ;
        RECT -43.005 20.235 -42.675 20.565 ;
        RECT -43.005 18.875 -42.675 19.205 ;
        RECT -43.005 17.515 -42.675 17.845 ;
        RECT -43.005 16.155 -42.675 16.485 ;
        RECT -43.005 14.795 -42.675 15.125 ;
        RECT -43.005 13.435 -42.675 13.765 ;
        RECT -43.005 12.075 -42.675 12.405 ;
        RECT -43.005 10.715 -42.675 11.045 ;
        RECT -43.005 9.355 -42.675 9.685 ;
        RECT -43.005 7.995 -42.675 8.325 ;
        RECT -43.005 6.635 -42.675 6.965 ;
        RECT -43.005 5.275 -42.675 5.605 ;
        RECT -43.005 3.915 -42.675 4.245 ;
        RECT -43.005 2.555 -42.675 2.885 ;
        RECT -43.005 1.195 -42.675 1.525 ;
        RECT -43.005 -0.165 -42.675 0.165 ;
        RECT -43.005 -1.525 -42.675 -1.195 ;
        RECT -43.005 -2.885 -42.675 -2.555 ;
        RECT -43.005 -4.245 -42.675 -3.915 ;
        RECT -43.005 -5.605 -42.675 -5.275 ;
        RECT -43.005 -6.965 -42.675 -6.635 ;
        RECT -43.005 -8.325 -42.675 -7.995 ;
        RECT -43.005 -9.685 -42.675 -9.355 ;
        RECT -43.005 -11.045 -42.675 -10.715 ;
        RECT -43.005 -12.405 -42.675 -12.075 ;
        RECT -43.005 -13.765 -42.675 -13.435 ;
        RECT -43.005 -15.125 -42.675 -14.795 ;
        RECT -43.005 -16.485 -42.675 -16.155 ;
        RECT -43.005 -17.845 -42.675 -17.515 ;
        RECT -43.005 -19.205 -42.675 -18.875 ;
        RECT -43.005 -20.565 -42.675 -20.235 ;
        RECT -43.005 -21.925 -42.675 -21.595 ;
        RECT -43.005 -23.285 -42.675 -22.955 ;
        RECT -43.005 -24.645 -42.675 -24.315 ;
        RECT -43.005 -27.365 -42.675 -27.035 ;
        RECT -43.005 -28.725 -42.675 -28.395 ;
        RECT -43.005 -30.085 -42.675 -29.755 ;
        RECT -43.005 -32.805 -42.675 -32.475 ;
        RECT -43.005 -35.525 -42.675 -35.195 ;
        RECT -43.005 -36.885 -42.675 -36.555 ;
        RECT -43.005 -39.605 -42.675 -39.275 ;
        RECT -43.005 -40.965 -42.675 -40.635 ;
        RECT -43.005 -42.325 -42.675 -41.995 ;
        RECT -43.005 -43.685 -42.675 -43.355 ;
        RECT -43.005 -45.045 -42.675 -44.715 ;
        RECT -43.005 -46.405 -42.675 -46.075 ;
        RECT -43.005 -47.765 -42.675 -47.435 ;
        RECT -43.005 -49.125 -42.675 -48.795 ;
        RECT -43.005 -50.485 -42.675 -50.155 ;
        RECT -43.005 -51.845 -42.675 -51.515 ;
        RECT -43.005 -53.205 -42.675 -52.875 ;
        RECT -43.005 -54.565 -42.675 -54.235 ;
        RECT -43.005 -55.925 -42.675 -55.595 ;
        RECT -43.005 -57.285 -42.675 -56.955 ;
        RECT -43.005 -58.645 -42.675 -58.315 ;
        RECT -43.005 -60.005 -42.675 -59.675 ;
        RECT -43.005 -61.365 -42.675 -61.035 ;
        RECT -43.005 -62.725 -42.675 -62.395 ;
        RECT -43.005 -64.085 -42.675 -63.755 ;
        RECT -43.005 -65.445 -42.675 -65.115 ;
        RECT -43.005 -66.805 -42.675 -66.475 ;
        RECT -43.005 -68.165 -42.675 -67.835 ;
        RECT -43.005 -69.525 -42.675 -69.195 ;
        RECT -43.005 -70.885 -42.675 -70.555 ;
        RECT -43.005 -72.245 -42.675 -71.915 ;
        RECT -43.005 -73.605 -42.675 -73.275 ;
        RECT -43.005 -74.965 -42.675 -74.635 ;
        RECT -43.005 -76.325 -42.675 -75.995 ;
        RECT -43.005 -77.685 -42.675 -77.355 ;
        RECT -43.005 -79.045 -42.675 -78.715 ;
        RECT -43.005 -80.405 -42.675 -80.075 ;
        RECT -43.005 -81.765 -42.675 -81.435 ;
        RECT -43.005 -83.125 -42.675 -82.795 ;
        RECT -43.005 -84.485 -42.675 -84.155 ;
        RECT -43.005 -85.845 -42.675 -85.515 ;
        RECT -43.005 -87.205 -42.675 -86.875 ;
        RECT -43.005 -88.565 -42.675 -88.235 ;
        RECT -43.005 -89.925 -42.675 -89.595 ;
        RECT -43.005 -91.285 -42.675 -90.955 ;
        RECT -43.005 -92.645 -42.675 -92.315 ;
        RECT -43.005 -94.005 -42.675 -93.675 ;
        RECT -43.005 -95.365 -42.675 -95.035 ;
        RECT -43.005 -96.725 -42.675 -96.395 ;
        RECT -43.005 -98.085 -42.675 -97.755 ;
        RECT -43.005 -99.445 -42.675 -99.115 ;
        RECT -43.005 -100.805 -42.675 -100.475 ;
        RECT -43.005 -102.165 -42.675 -101.835 ;
        RECT -43.005 -103.525 -42.675 -103.195 ;
        RECT -43.005 -104.885 -42.675 -104.555 ;
        RECT -43.005 -106.245 -42.675 -105.915 ;
        RECT -43.005 -107.605 -42.675 -107.275 ;
        RECT -43.005 -108.965 -42.675 -108.635 ;
        RECT -43.005 -110.325 -42.675 -109.995 ;
        RECT -43.005 -113.045 -42.675 -112.715 ;
        RECT -43.005 -114.405 -42.675 -114.075 ;
        RECT -43.005 -115.765 -42.675 -115.435 ;
        RECT -43.005 -117.125 -42.675 -116.795 ;
        RECT -43.005 -118.485 -42.675 -118.155 ;
        RECT -43.005 -119.79 -42.675 -119.46 ;
        RECT -43.005 -121.205 -42.675 -120.875 ;
        RECT -43.005 -122.565 -42.675 -122.235 ;
        RECT -43.005 -123.925 -42.675 -123.595 ;
        RECT -43.005 -126.645 -42.675 -126.315 ;
        RECT -43.005 -128.43 -42.675 -128.1 ;
        RECT -43.005 -129.365 -42.675 -129.035 ;
        RECT -43.005 -130.725 -42.675 -130.395 ;
        RECT -43.005 -133.445 -42.675 -133.115 ;
        RECT -43.005 -134.805 -42.675 -134.475 ;
        RECT -43.005 -136.165 -42.675 -135.835 ;
        RECT -43.005 -137.525 -42.675 -137.195 ;
        RECT -43.005 -140.245 -42.675 -139.915 ;
        RECT -43.005 -142.965 -42.675 -142.635 ;
        RECT -43.005 -144.325 -42.675 -143.995 ;
        RECT -43.005 -145.685 -42.675 -145.355 ;
        RECT -43.005 -147.045 -42.675 -146.715 ;
        RECT -43.005 -148.405 -42.675 -148.075 ;
        RECT -43.005 -149.765 -42.675 -149.435 ;
        RECT -43.005 -151.125 -42.675 -150.795 ;
        RECT -43.005 -152.485 -42.675 -152.155 ;
        RECT -43.005 -153.845 -42.675 -153.515 ;
        RECT -43.005 -155.205 -42.675 -154.875 ;
        RECT -43.005 -156.565 -42.675 -156.235 ;
        RECT -43.005 -157.925 -42.675 -157.595 ;
        RECT -43.005 -159.285 -42.675 -158.955 ;
        RECT -43.005 -160.645 -42.675 -160.315 ;
        RECT -43.005 -162.005 -42.675 -161.675 ;
        RECT -43.005 -163.365 -42.675 -163.035 ;
        RECT -43.005 -164.725 -42.675 -164.395 ;
        RECT -43.005 -166.085 -42.675 -165.755 ;
        RECT -43.005 -167.445 -42.675 -167.115 ;
        RECT -43.005 -168.805 -42.675 -168.475 ;
        RECT -43.005 -170.165 -42.675 -169.835 ;
        RECT -43.005 -171.525 -42.675 -171.195 ;
        RECT -43.005 -172.885 -42.675 -172.555 ;
        RECT -43.005 -174.245 -42.675 -173.915 ;
        RECT -43.005 -175.605 -42.675 -175.275 ;
        RECT -43.005 -176.965 -42.675 -176.635 ;
        RECT -43.005 -178.325 -42.675 -177.995 ;
        RECT -43.005 -179.685 -42.675 -179.355 ;
        RECT -43.005 -181.045 -42.675 -180.715 ;
        RECT -43.005 -182.405 -42.675 -182.075 ;
        RECT -43.005 -183.765 -42.675 -183.435 ;
        RECT -43.005 -185.125 -42.675 -184.795 ;
        RECT -43.005 -186.485 -42.675 -186.155 ;
        RECT -43.005 -187.845 -42.675 -187.515 ;
        RECT -43.005 -189.205 -42.675 -188.875 ;
        RECT -43.005 -190.565 -42.675 -190.235 ;
        RECT -43.005 -191.925 -42.675 -191.595 ;
        RECT -43.005 -193.285 -42.675 -192.955 ;
        RECT -43.005 -194.645 -42.675 -194.315 ;
        RECT -43.005 -196.005 -42.675 -195.675 ;
        RECT -43.005 -197.365 -42.675 -197.035 ;
        RECT -43.005 -198.725 -42.675 -198.395 ;
        RECT -43.005 -200.085 -42.675 -199.755 ;
        RECT -43.005 -201.445 -42.675 -201.115 ;
        RECT -43.005 -202.805 -42.675 -202.475 ;
        RECT -43.005 -204.165 -42.675 -203.835 ;
        RECT -43.005 -205.525 -42.675 -205.195 ;
        RECT -43.005 -208.245 -42.675 -207.915 ;
        RECT -43.005 -210.965 -42.675 -210.635 ;
        RECT -43.005 -212.325 -42.675 -211.995 ;
        RECT -43.005 -213.625 -42.675 -213.295 ;
        RECT -43.005 -215.045 -42.675 -214.715 ;
        RECT -43.005 -216.405 -42.675 -216.075 ;
        RECT -43.005 -217.765 -42.675 -217.435 ;
        RECT -43.005 -219.125 -42.675 -218.795 ;
        RECT -43.005 -221.37 -42.675 -220.24 ;
        RECT -43 -221.485 -42.68 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -41.645 129.8 -41.315 130.93 ;
        RECT -41.645 127.675 -41.315 128.005 ;
        RECT -41.645 126.315 -41.315 126.645 ;
        RECT -41.645 124.955 -41.315 125.285 ;
        RECT -41.645 123.595 -41.315 123.925 ;
        RECT -41.645 122.235 -41.315 122.565 ;
        RECT -41.645 120.875 -41.315 121.205 ;
        RECT -41.645 119.515 -41.315 119.845 ;
        RECT -41.645 118.155 -41.315 118.485 ;
        RECT -41.645 116.795 -41.315 117.125 ;
        RECT -41.645 115.435 -41.315 115.765 ;
        RECT -41.645 114.075 -41.315 114.405 ;
        RECT -41.645 112.715 -41.315 113.045 ;
        RECT -41.645 111.355 -41.315 111.685 ;
        RECT -41.645 109.995 -41.315 110.325 ;
        RECT -41.645 108.635 -41.315 108.965 ;
        RECT -41.645 107.275 -41.315 107.605 ;
        RECT -41.645 105.915 -41.315 106.245 ;
        RECT -41.645 104.555 -41.315 104.885 ;
        RECT -41.645 103.195 -41.315 103.525 ;
        RECT -41.645 101.835 -41.315 102.165 ;
        RECT -41.645 100.475 -41.315 100.805 ;
        RECT -41.645 99.115 -41.315 99.445 ;
        RECT -41.645 97.755 -41.315 98.085 ;
        RECT -41.645 96.395 -41.315 96.725 ;
        RECT -41.645 95.035 -41.315 95.365 ;
        RECT -41.645 93.675 -41.315 94.005 ;
        RECT -41.645 92.315 -41.315 92.645 ;
        RECT -41.645 90.955 -41.315 91.285 ;
        RECT -41.645 89.595 -41.315 89.925 ;
        RECT -41.645 88.235 -41.315 88.565 ;
        RECT -41.645 86.875 -41.315 87.205 ;
        RECT -41.645 85.515 -41.315 85.845 ;
        RECT -41.645 84.155 -41.315 84.485 ;
        RECT -41.645 82.795 -41.315 83.125 ;
        RECT -41.645 81.435 -41.315 81.765 ;
        RECT -41.645 80.075 -41.315 80.405 ;
        RECT -41.645 78.715 -41.315 79.045 ;
        RECT -41.645 77.355 -41.315 77.685 ;
        RECT -41.645 75.995 -41.315 76.325 ;
        RECT -41.645 74.635 -41.315 74.965 ;
        RECT -41.645 73.275 -41.315 73.605 ;
        RECT -41.645 72.445 -41.315 72.775 ;
        RECT -41.645 70.395 -41.315 70.725 ;
        RECT -41.645 68.035 -41.315 68.365 ;
        RECT -41.645 66.885 -41.315 67.215 ;
        RECT -41.645 64.875 -41.315 65.205 ;
        RECT -41.645 63.725 -41.315 64.055 ;
        RECT -41.645 61.715 -41.315 62.045 ;
        RECT -41.645 60.395 -41.315 60.725 ;
        RECT -41.645 58.555 -41.315 58.885 ;
        RECT -41.645 57.405 -41.315 57.735 ;
        RECT -41.645 55.395 -41.315 55.725 ;
        RECT -41.645 54.245 -41.315 54.575 ;
        RECT -41.645 51.885 -41.315 52.215 ;
        RECT -41.645 49.83 -41.315 50.16 ;
        RECT -41.645 48.795 -41.315 49.125 ;
        RECT -41.645 47.435 -41.315 47.765 ;
        RECT -41.645 46.075 -41.315 46.405 ;
        RECT -41.645 44.715 -41.315 45.045 ;
        RECT -41.645 43.355 -41.315 43.685 ;
        RECT -41.645 41.995 -41.315 42.325 ;
        RECT -41.645 40.635 -41.315 40.965 ;
        RECT -41.645 39.275 -41.315 39.605 ;
        RECT -41.645 37.915 -41.315 38.245 ;
        RECT -41.645 36.555 -41.315 36.885 ;
        RECT -41.645 35.195 -41.315 35.525 ;
        RECT -41.645 33.835 -41.315 34.165 ;
        RECT -41.645 32.475 -41.315 32.805 ;
        RECT -41.645 31.115 -41.315 31.445 ;
        RECT -41.645 29.755 -41.315 30.085 ;
        RECT -41.645 28.395 -41.315 28.725 ;
        RECT -41.645 27.035 -41.315 27.365 ;
        RECT -41.645 25.675 -41.315 26.005 ;
        RECT -41.645 24.315 -41.315 24.645 ;
        RECT -41.645 22.955 -41.315 23.285 ;
        RECT -41.645 21.595 -41.315 21.925 ;
        RECT -41.645 20.235 -41.315 20.565 ;
        RECT -41.645 18.875 -41.315 19.205 ;
        RECT -41.645 17.515 -41.315 17.845 ;
        RECT -41.645 16.155 -41.315 16.485 ;
        RECT -41.645 14.795 -41.315 15.125 ;
        RECT -41.645 13.435 -41.315 13.765 ;
        RECT -41.645 12.075 -41.315 12.405 ;
        RECT -41.645 10.715 -41.315 11.045 ;
        RECT -41.645 9.355 -41.315 9.685 ;
        RECT -41.645 7.995 -41.315 8.325 ;
        RECT -41.645 6.635 -41.315 6.965 ;
        RECT -41.645 5.275 -41.315 5.605 ;
        RECT -41.645 3.915 -41.315 4.245 ;
        RECT -41.645 2.555 -41.315 2.885 ;
        RECT -41.645 1.195 -41.315 1.525 ;
        RECT -41.645 -0.165 -41.315 0.165 ;
        RECT -41.645 -1.525 -41.315 -1.195 ;
        RECT -41.645 -2.885 -41.315 -2.555 ;
        RECT -41.645 -4.245 -41.315 -3.915 ;
        RECT -41.645 -5.605 -41.315 -5.275 ;
        RECT -41.645 -6.965 -41.315 -6.635 ;
        RECT -41.645 -8.325 -41.315 -7.995 ;
        RECT -41.645 -9.685 -41.315 -9.355 ;
        RECT -41.645 -11.045 -41.315 -10.715 ;
        RECT -41.645 -12.405 -41.315 -12.075 ;
        RECT -41.645 -13.765 -41.315 -13.435 ;
        RECT -41.645 -15.125 -41.315 -14.795 ;
        RECT -41.645 -16.485 -41.315 -16.155 ;
        RECT -41.645 -17.845 -41.315 -17.515 ;
        RECT -41.645 -19.205 -41.315 -18.875 ;
        RECT -41.645 -20.565 -41.315 -20.235 ;
        RECT -41.645 -21.925 -41.315 -21.595 ;
        RECT -41.645 -23.285 -41.315 -22.955 ;
        RECT -41.645 -27.365 -41.315 -27.035 ;
        RECT -41.645 -28.725 -41.315 -28.395 ;
        RECT -41.645 -30.085 -41.315 -29.755 ;
        RECT -41.645 -32.805 -41.315 -32.475 ;
        RECT -41.645 -35.525 -41.315 -35.195 ;
        RECT -41.645 -36.885 -41.315 -36.555 ;
        RECT -41.645 -39.605 -41.315 -39.275 ;
        RECT -41.645 -40.965 -41.315 -40.635 ;
        RECT -41.645 -42.325 -41.315 -41.995 ;
        RECT -41.645 -43.685 -41.315 -43.355 ;
        RECT -41.645 -45.045 -41.315 -44.715 ;
        RECT -41.645 -46.405 -41.315 -46.075 ;
        RECT -41.645 -47.765 -41.315 -47.435 ;
        RECT -41.645 -49.125 -41.315 -48.795 ;
        RECT -41.645 -50.485 -41.315 -50.155 ;
        RECT -41.645 -51.845 -41.315 -51.515 ;
        RECT -41.645 -53.205 -41.315 -52.875 ;
        RECT -41.645 -54.565 -41.315 -54.235 ;
        RECT -41.645 -55.925 -41.315 -55.595 ;
        RECT -41.645 -57.285 -41.315 -56.955 ;
        RECT -41.645 -58.645 -41.315 -58.315 ;
        RECT -41.645 -60.005 -41.315 -59.675 ;
        RECT -41.645 -61.365 -41.315 -61.035 ;
        RECT -41.645 -62.725 -41.315 -62.395 ;
        RECT -41.645 -64.085 -41.315 -63.755 ;
        RECT -41.645 -65.445 -41.315 -65.115 ;
        RECT -41.645 -66.805 -41.315 -66.475 ;
        RECT -41.645 -68.165 -41.315 -67.835 ;
        RECT -41.645 -69.525 -41.315 -69.195 ;
        RECT -41.645 -70.885 -41.315 -70.555 ;
        RECT -41.645 -72.245 -41.315 -71.915 ;
        RECT -41.645 -73.605 -41.315 -73.275 ;
        RECT -41.645 -74.965 -41.315 -74.635 ;
        RECT -41.645 -76.325 -41.315 -75.995 ;
        RECT -41.645 -77.685 -41.315 -77.355 ;
        RECT -41.645 -79.045 -41.315 -78.715 ;
        RECT -41.645 -80.405 -41.315 -80.075 ;
        RECT -41.645 -81.765 -41.315 -81.435 ;
        RECT -41.645 -83.125 -41.315 -82.795 ;
        RECT -41.645 -84.485 -41.315 -84.155 ;
        RECT -41.645 -85.845 -41.315 -85.515 ;
        RECT -41.645 -87.205 -41.315 -86.875 ;
        RECT -41.645 -88.565 -41.315 -88.235 ;
        RECT -41.645 -89.925 -41.315 -89.595 ;
        RECT -41.645 -91.285 -41.315 -90.955 ;
        RECT -41.645 -92.645 -41.315 -92.315 ;
        RECT -41.645 -94.005 -41.315 -93.675 ;
        RECT -41.645 -95.365 -41.315 -95.035 ;
        RECT -41.645 -96.725 -41.315 -96.395 ;
        RECT -41.645 -98.085 -41.315 -97.755 ;
        RECT -41.645 -99.445 -41.315 -99.115 ;
        RECT -41.645 -100.805 -41.315 -100.475 ;
        RECT -41.645 -102.165 -41.315 -101.835 ;
        RECT -41.645 -103.525 -41.315 -103.195 ;
        RECT -41.645 -104.885 -41.315 -104.555 ;
        RECT -41.645 -106.245 -41.315 -105.915 ;
        RECT -41.645 -107.605 -41.315 -107.275 ;
        RECT -41.645 -108.965 -41.315 -108.635 ;
        RECT -41.645 -110.325 -41.315 -109.995 ;
        RECT -41.645 -113.045 -41.315 -112.715 ;
        RECT -41.645 -114.405 -41.315 -114.075 ;
        RECT -41.645 -115.765 -41.315 -115.435 ;
        RECT -41.645 -117.125 -41.315 -116.795 ;
        RECT -41.645 -118.485 -41.315 -118.155 ;
        RECT -41.645 -119.79 -41.315 -119.46 ;
        RECT -41.645 -121.205 -41.315 -120.875 ;
        RECT -41.645 -122.565 -41.315 -122.235 ;
        RECT -41.645 -123.925 -41.315 -123.595 ;
        RECT -41.645 -126.645 -41.315 -126.315 ;
        RECT -41.645 -128.43 -41.315 -128.1 ;
        RECT -41.645 -129.365 -41.315 -129.035 ;
        RECT -41.645 -130.725 -41.315 -130.395 ;
        RECT -41.64 -132.08 -41.32 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -41.645 -212.325 -41.315 -211.995 ;
        RECT -41.645 -213.625 -41.315 -213.295 ;
        RECT -41.645 -215.045 -41.315 -214.715 ;
        RECT -41.645 -216.405 -41.315 -216.075 ;
        RECT -41.645 -217.765 -41.315 -217.435 ;
        RECT -41.645 -219.125 -41.315 -218.795 ;
        RECT -41.645 -221.37 -41.315 -220.24 ;
        RECT -41.64 -221.485 -41.32 -210.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -40.285 -186.485 -39.955 -186.155 ;
        RECT -40.285 -187.845 -39.955 -187.515 ;
        RECT -40.285 -189.205 -39.955 -188.875 ;
        RECT -40.285 -190.565 -39.955 -190.235 ;
        RECT -40.285 -191.925 -39.955 -191.595 ;
        RECT -40.285 -193.285 -39.955 -192.955 ;
        RECT -40.285 -194.645 -39.955 -194.315 ;
        RECT -40.285 -196.005 -39.955 -195.675 ;
        RECT -40.285 -197.365 -39.955 -197.035 ;
        RECT -40.285 -198.725 -39.955 -198.395 ;
        RECT -40.285 -200.085 -39.955 -199.755 ;
        RECT -40.285 -201.445 -39.955 -201.115 ;
        RECT -40.285 -202.805 -39.955 -202.475 ;
        RECT -40.285 -204.165 -39.955 -203.835 ;
        RECT -40.285 -205.525 -39.955 -205.195 ;
        RECT -40.285 -208.245 -39.955 -207.915 ;
        RECT -40.28 -209.6 -39.96 131.045 ;
        RECT -40.285 129.8 -39.955 130.93 ;
        RECT -40.285 127.675 -39.955 128.005 ;
        RECT -40.285 126.315 -39.955 126.645 ;
        RECT -40.285 124.955 -39.955 125.285 ;
        RECT -40.285 123.595 -39.955 123.925 ;
        RECT -40.285 122.235 -39.955 122.565 ;
        RECT -40.285 120.875 -39.955 121.205 ;
        RECT -40.285 119.515 -39.955 119.845 ;
        RECT -40.285 118.155 -39.955 118.485 ;
        RECT -40.285 116.795 -39.955 117.125 ;
        RECT -40.285 115.435 -39.955 115.765 ;
        RECT -40.285 114.075 -39.955 114.405 ;
        RECT -40.285 112.715 -39.955 113.045 ;
        RECT -40.285 111.355 -39.955 111.685 ;
        RECT -40.285 109.995 -39.955 110.325 ;
        RECT -40.285 108.635 -39.955 108.965 ;
        RECT -40.285 107.275 -39.955 107.605 ;
        RECT -40.285 105.915 -39.955 106.245 ;
        RECT -40.285 104.555 -39.955 104.885 ;
        RECT -40.285 103.195 -39.955 103.525 ;
        RECT -40.285 101.835 -39.955 102.165 ;
        RECT -40.285 100.475 -39.955 100.805 ;
        RECT -40.285 99.115 -39.955 99.445 ;
        RECT -40.285 97.755 -39.955 98.085 ;
        RECT -40.285 96.395 -39.955 96.725 ;
        RECT -40.285 95.035 -39.955 95.365 ;
        RECT -40.285 93.675 -39.955 94.005 ;
        RECT -40.285 92.315 -39.955 92.645 ;
        RECT -40.285 90.955 -39.955 91.285 ;
        RECT -40.285 89.595 -39.955 89.925 ;
        RECT -40.285 88.235 -39.955 88.565 ;
        RECT -40.285 86.875 -39.955 87.205 ;
        RECT -40.285 85.515 -39.955 85.845 ;
        RECT -40.285 84.155 -39.955 84.485 ;
        RECT -40.285 82.795 -39.955 83.125 ;
        RECT -40.285 81.435 -39.955 81.765 ;
        RECT -40.285 80.075 -39.955 80.405 ;
        RECT -40.285 78.715 -39.955 79.045 ;
        RECT -40.285 77.355 -39.955 77.685 ;
        RECT -40.285 75.995 -39.955 76.325 ;
        RECT -40.285 74.635 -39.955 74.965 ;
        RECT -40.285 73.275 -39.955 73.605 ;
        RECT -40.285 48.795 -39.955 49.125 ;
        RECT -40.285 47.435 -39.955 47.765 ;
        RECT -40.285 46.075 -39.955 46.405 ;
        RECT -40.285 44.715 -39.955 45.045 ;
        RECT -40.285 43.355 -39.955 43.685 ;
        RECT -40.285 41.995 -39.955 42.325 ;
        RECT -40.285 40.635 -39.955 40.965 ;
        RECT -40.285 39.275 -39.955 39.605 ;
        RECT -40.285 37.915 -39.955 38.245 ;
        RECT -40.285 36.555 -39.955 36.885 ;
        RECT -40.285 35.195 -39.955 35.525 ;
        RECT -40.285 33.835 -39.955 34.165 ;
        RECT -40.285 32.475 -39.955 32.805 ;
        RECT -40.285 31.115 -39.955 31.445 ;
        RECT -40.285 29.755 -39.955 30.085 ;
        RECT -40.285 28.395 -39.955 28.725 ;
        RECT -40.285 27.035 -39.955 27.365 ;
        RECT -40.285 25.675 -39.955 26.005 ;
        RECT -40.285 24.315 -39.955 24.645 ;
        RECT -40.285 22.955 -39.955 23.285 ;
        RECT -40.285 21.595 -39.955 21.925 ;
        RECT -40.285 20.235 -39.955 20.565 ;
        RECT -40.285 18.875 -39.955 19.205 ;
        RECT -40.285 17.515 -39.955 17.845 ;
        RECT -40.285 16.155 -39.955 16.485 ;
        RECT -40.285 14.795 -39.955 15.125 ;
        RECT -40.285 13.435 -39.955 13.765 ;
        RECT -40.285 12.075 -39.955 12.405 ;
        RECT -40.285 10.715 -39.955 11.045 ;
        RECT -40.285 9.355 -39.955 9.685 ;
        RECT -40.285 7.995 -39.955 8.325 ;
        RECT -40.285 6.635 -39.955 6.965 ;
        RECT -40.285 5.275 -39.955 5.605 ;
        RECT -40.285 3.915 -39.955 4.245 ;
        RECT -40.285 2.555 -39.955 2.885 ;
        RECT -40.285 1.195 -39.955 1.525 ;
        RECT -40.285 -0.165 -39.955 0.165 ;
        RECT -40.285 -1.525 -39.955 -1.195 ;
        RECT -40.285 -2.885 -39.955 -2.555 ;
        RECT -40.285 -4.245 -39.955 -3.915 ;
        RECT -40.285 -5.605 -39.955 -5.275 ;
        RECT -40.285 -6.965 -39.955 -6.635 ;
        RECT -40.285 -8.325 -39.955 -7.995 ;
        RECT -40.285 -9.685 -39.955 -9.355 ;
        RECT -40.285 -11.045 -39.955 -10.715 ;
        RECT -40.285 -12.405 -39.955 -12.075 ;
        RECT -40.285 -13.765 -39.955 -13.435 ;
        RECT -40.285 -15.125 -39.955 -14.795 ;
        RECT -40.285 -16.485 -39.955 -16.155 ;
        RECT -40.285 -17.845 -39.955 -17.515 ;
        RECT -40.285 -19.205 -39.955 -18.875 ;
        RECT -40.285 -20.565 -39.955 -20.235 ;
        RECT -40.285 -21.925 -39.955 -21.595 ;
        RECT -40.285 -27.365 -39.955 -27.035 ;
        RECT -40.285 -28.725 -39.955 -28.395 ;
        RECT -40.285 -30.085 -39.955 -29.755 ;
        RECT -40.285 -32.805 -39.955 -32.475 ;
        RECT -40.285 -35.525 -39.955 -35.195 ;
        RECT -40.285 -36.885 -39.955 -36.555 ;
        RECT -40.285 -39.605 -39.955 -39.275 ;
        RECT -40.285 -40.965 -39.955 -40.635 ;
        RECT -40.285 -42.325 -39.955 -41.995 ;
        RECT -40.285 -43.685 -39.955 -43.355 ;
        RECT -40.285 -45.045 -39.955 -44.715 ;
        RECT -40.285 -46.405 -39.955 -46.075 ;
        RECT -40.285 -47.765 -39.955 -47.435 ;
        RECT -40.285 -49.125 -39.955 -48.795 ;
        RECT -40.285 -50.485 -39.955 -50.155 ;
        RECT -40.285 -51.845 -39.955 -51.515 ;
        RECT -40.285 -53.205 -39.955 -52.875 ;
        RECT -40.285 -54.565 -39.955 -54.235 ;
        RECT -40.285 -55.925 -39.955 -55.595 ;
        RECT -40.285 -57.285 -39.955 -56.955 ;
        RECT -40.285 -58.645 -39.955 -58.315 ;
        RECT -40.285 -60.005 -39.955 -59.675 ;
        RECT -40.285 -61.365 -39.955 -61.035 ;
        RECT -40.285 -62.725 -39.955 -62.395 ;
        RECT -40.285 -64.085 -39.955 -63.755 ;
        RECT -40.285 -65.445 -39.955 -65.115 ;
        RECT -40.285 -66.805 -39.955 -66.475 ;
        RECT -40.285 -68.165 -39.955 -67.835 ;
        RECT -40.285 -69.525 -39.955 -69.195 ;
        RECT -40.285 -70.885 -39.955 -70.555 ;
        RECT -40.285 -72.245 -39.955 -71.915 ;
        RECT -40.285 -73.605 -39.955 -73.275 ;
        RECT -40.285 -74.965 -39.955 -74.635 ;
        RECT -40.285 -76.325 -39.955 -75.995 ;
        RECT -40.285 -77.685 -39.955 -77.355 ;
        RECT -40.285 -79.045 -39.955 -78.715 ;
        RECT -40.285 -80.405 -39.955 -80.075 ;
        RECT -40.285 -81.765 -39.955 -81.435 ;
        RECT -40.285 -83.125 -39.955 -82.795 ;
        RECT -40.285 -84.485 -39.955 -84.155 ;
        RECT -40.285 -85.845 -39.955 -85.515 ;
        RECT -40.285 -87.205 -39.955 -86.875 ;
        RECT -40.285 -88.565 -39.955 -88.235 ;
        RECT -40.285 -89.925 -39.955 -89.595 ;
        RECT -40.285 -91.285 -39.955 -90.955 ;
        RECT -40.285 -92.645 -39.955 -92.315 ;
        RECT -40.285 -94.005 -39.955 -93.675 ;
        RECT -40.285 -95.365 -39.955 -95.035 ;
        RECT -40.285 -96.725 -39.955 -96.395 ;
        RECT -40.285 -98.085 -39.955 -97.755 ;
        RECT -40.285 -99.445 -39.955 -99.115 ;
        RECT -40.285 -100.805 -39.955 -100.475 ;
        RECT -40.285 -102.165 -39.955 -101.835 ;
        RECT -40.285 -103.525 -39.955 -103.195 ;
        RECT -40.285 -104.885 -39.955 -104.555 ;
        RECT -40.285 -106.245 -39.955 -105.915 ;
        RECT -40.285 -107.605 -39.955 -107.275 ;
        RECT -40.285 -108.965 -39.955 -108.635 ;
        RECT -40.285 -110.325 -39.955 -109.995 ;
        RECT -40.285 -113.045 -39.955 -112.715 ;
        RECT -40.285 -114.405 -39.955 -114.075 ;
        RECT -40.285 -115.765 -39.955 -115.435 ;
        RECT -40.285 -117.125 -39.955 -116.795 ;
        RECT -40.285 -118.485 -39.955 -118.155 ;
        RECT -40.285 -119.79 -39.955 -119.46 ;
        RECT -40.285 -121.205 -39.955 -120.875 ;
        RECT -40.285 -122.565 -39.955 -122.235 ;
        RECT -40.285 -123.925 -39.955 -123.595 ;
        RECT -40.285 -126.645 -39.955 -126.315 ;
        RECT -40.285 -128.43 -39.955 -128.1 ;
        RECT -40.285 -129.365 -39.955 -129.035 ;
        RECT -40.285 -130.725 -39.955 -130.395 ;
        RECT -40.285 -133.445 -39.955 -133.115 ;
        RECT -40.285 -134.805 -39.955 -134.475 ;
        RECT -40.285 -136.165 -39.955 -135.835 ;
        RECT -40.285 -137.525 -39.955 -137.195 ;
        RECT -40.285 -140.245 -39.955 -139.915 ;
        RECT -40.285 -142.965 -39.955 -142.635 ;
        RECT -40.285 -144.325 -39.955 -143.995 ;
        RECT -40.285 -145.685 -39.955 -145.355 ;
        RECT -40.285 -147.045 -39.955 -146.715 ;
        RECT -40.285 -148.405 -39.955 -148.075 ;
        RECT -40.285 -149.765 -39.955 -149.435 ;
        RECT -40.285 -151.125 -39.955 -150.795 ;
        RECT -40.285 -152.485 -39.955 -152.155 ;
        RECT -40.285 -153.845 -39.955 -153.515 ;
        RECT -40.285 -155.205 -39.955 -154.875 ;
        RECT -40.285 -156.565 -39.955 -156.235 ;
        RECT -40.285 -157.925 -39.955 -157.595 ;
        RECT -40.285 -159.285 -39.955 -158.955 ;
        RECT -40.285 -160.645 -39.955 -160.315 ;
        RECT -40.285 -162.005 -39.955 -161.675 ;
        RECT -40.285 -163.365 -39.955 -163.035 ;
        RECT -40.285 -164.725 -39.955 -164.395 ;
        RECT -40.285 -166.085 -39.955 -165.755 ;
        RECT -40.285 -167.445 -39.955 -167.115 ;
        RECT -40.285 -168.805 -39.955 -168.475 ;
        RECT -40.285 -170.165 -39.955 -169.835 ;
        RECT -40.285 -171.525 -39.955 -171.195 ;
        RECT -40.285 -172.885 -39.955 -172.555 ;
        RECT -40.285 -174.245 -39.955 -173.915 ;
        RECT -40.285 -175.605 -39.955 -175.275 ;
        RECT -40.285 -176.965 -39.955 -176.635 ;
        RECT -40.285 -178.325 -39.955 -177.995 ;
        RECT -40.285 -179.685 -39.955 -179.355 ;
        RECT -40.285 -181.045 -39.955 -180.715 ;
        RECT -40.285 -182.405 -39.955 -182.075 ;
        RECT -40.285 -183.765 -39.955 -183.435 ;
        RECT -40.285 -185.125 -39.955 -184.795 ;
    END
    PORT
      LAYER met3 ;
        RECT -52.525 129.8 -52.195 130.93 ;
        RECT -52.525 127.675 -52.195 128.005 ;
        RECT -52.525 126.315 -52.195 126.645 ;
        RECT -52.525 124.955 -52.195 125.285 ;
        RECT -52.525 123.595 -52.195 123.925 ;
        RECT -52.525 122.235 -52.195 122.565 ;
        RECT -52.525 120.875 -52.195 121.205 ;
        RECT -52.525 119.515 -52.195 119.845 ;
        RECT -52.525 118.155 -52.195 118.485 ;
        RECT -52.525 116.795 -52.195 117.125 ;
        RECT -52.525 115.435 -52.195 115.765 ;
        RECT -52.525 114.075 -52.195 114.405 ;
        RECT -52.525 112.715 -52.195 113.045 ;
        RECT -52.525 111.355 -52.195 111.685 ;
        RECT -52.525 109.995 -52.195 110.325 ;
        RECT -52.525 108.635 -52.195 108.965 ;
        RECT -52.525 107.275 -52.195 107.605 ;
        RECT -52.525 105.915 -52.195 106.245 ;
        RECT -52.525 104.555 -52.195 104.885 ;
        RECT -52.525 103.195 -52.195 103.525 ;
        RECT -52.525 101.835 -52.195 102.165 ;
        RECT -52.525 100.475 -52.195 100.805 ;
        RECT -52.525 99.115 -52.195 99.445 ;
        RECT -52.525 97.755 -52.195 98.085 ;
        RECT -52.525 96.395 -52.195 96.725 ;
        RECT -52.525 95.035 -52.195 95.365 ;
        RECT -52.525 93.675 -52.195 94.005 ;
        RECT -52.525 92.315 -52.195 92.645 ;
        RECT -52.525 90.955 -52.195 91.285 ;
        RECT -52.525 89.595 -52.195 89.925 ;
        RECT -52.525 88.235 -52.195 88.565 ;
        RECT -52.525 86.875 -52.195 87.205 ;
        RECT -52.525 85.515 -52.195 85.845 ;
        RECT -52.525 84.155 -52.195 84.485 ;
        RECT -52.525 82.795 -52.195 83.125 ;
        RECT -52.525 81.435 -52.195 81.765 ;
        RECT -52.525 80.075 -52.195 80.405 ;
        RECT -52.525 78.715 -52.195 79.045 ;
        RECT -52.525 77.355 -52.195 77.685 ;
        RECT -52.525 75.995 -52.195 76.325 ;
        RECT -52.525 74.635 -52.195 74.965 ;
        RECT -52.525 73.275 -52.195 73.605 ;
        RECT -52.525 72.445 -52.195 72.775 ;
        RECT -52.525 70.395 -52.195 70.725 ;
        RECT -52.525 68.035 -52.195 68.365 ;
        RECT -52.525 66.885 -52.195 67.215 ;
        RECT -52.525 64.875 -52.195 65.205 ;
        RECT -52.525 63.725 -52.195 64.055 ;
        RECT -52.525 61.715 -52.195 62.045 ;
        RECT -52.525 60.395 -52.195 60.725 ;
        RECT -52.525 58.555 -52.195 58.885 ;
        RECT -52.525 57.405 -52.195 57.735 ;
        RECT -52.525 55.395 -52.195 55.725 ;
        RECT -52.525 54.245 -52.195 54.575 ;
        RECT -52.525 51.885 -52.195 52.215 ;
        RECT -52.525 49.83 -52.195 50.16 ;
        RECT -52.525 48.795 -52.195 49.125 ;
        RECT -52.525 47.435 -52.195 47.765 ;
        RECT -52.525 46.075 -52.195 46.405 ;
        RECT -52.525 44.715 -52.195 45.045 ;
        RECT -52.525 43.355 -52.195 43.685 ;
        RECT -52.525 41.995 -52.195 42.325 ;
        RECT -52.525 40.635 -52.195 40.965 ;
        RECT -52.525 39.275 -52.195 39.605 ;
        RECT -52.52 37.92 -52.2 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -52.525 -142.965 -52.195 -142.635 ;
        RECT -52.525 -144.325 -52.195 -143.995 ;
        RECT -52.525 -145.685 -52.195 -145.355 ;
        RECT -52.525 -147.045 -52.195 -146.715 ;
        RECT -52.525 -148.405 -52.195 -148.075 ;
        RECT -52.525 -149.765 -52.195 -149.435 ;
        RECT -52.525 -151.125 -52.195 -150.795 ;
        RECT -52.525 -152.485 -52.195 -152.155 ;
        RECT -52.525 -153.845 -52.195 -153.515 ;
        RECT -52.525 -155.205 -52.195 -154.875 ;
        RECT -52.525 -156.565 -52.195 -156.235 ;
        RECT -52.525 -157.925 -52.195 -157.595 ;
        RECT -52.525 -159.285 -52.195 -158.955 ;
        RECT -52.525 -160.645 -52.195 -160.315 ;
        RECT -52.525 -162.005 -52.195 -161.675 ;
        RECT -52.525 -163.365 -52.195 -163.035 ;
        RECT -52.525 -164.725 -52.195 -164.395 ;
        RECT -52.525 -166.085 -52.195 -165.755 ;
        RECT -52.525 -167.445 -52.195 -167.115 ;
        RECT -52.525 -168.805 -52.195 -168.475 ;
        RECT -52.525 -170.165 -52.195 -169.835 ;
        RECT -52.525 -171.525 -52.195 -171.195 ;
        RECT -52.525 -172.885 -52.195 -172.555 ;
        RECT -52.525 -174.245 -52.195 -173.915 ;
        RECT -52.525 -175.605 -52.195 -175.275 ;
        RECT -52.525 -176.965 -52.195 -176.635 ;
        RECT -52.525 -178.325 -52.195 -177.995 ;
        RECT -52.525 -179.685 -52.195 -179.355 ;
        RECT -52.525 -181.045 -52.195 -180.715 ;
        RECT -52.525 -182.405 -52.195 -182.075 ;
        RECT -52.525 -183.765 -52.195 -183.435 ;
        RECT -52.525 -185.125 -52.195 -184.795 ;
        RECT -52.525 -186.485 -52.195 -186.155 ;
        RECT -52.525 -187.845 -52.195 -187.515 ;
        RECT -52.525 -189.205 -52.195 -188.875 ;
        RECT -52.525 -190.565 -52.195 -190.235 ;
        RECT -52.525 -191.925 -52.195 -191.595 ;
        RECT -52.525 -193.285 -52.195 -192.955 ;
        RECT -52.525 -194.645 -52.195 -194.315 ;
        RECT -52.525 -196.005 -52.195 -195.675 ;
        RECT -52.525 -197.365 -52.195 -197.035 ;
        RECT -52.525 -198.725 -52.195 -198.395 ;
        RECT -52.525 -200.085 -52.195 -199.755 ;
        RECT -52.525 -201.445 -52.195 -201.115 ;
        RECT -52.525 -202.805 -52.195 -202.475 ;
        RECT -52.525 -204.165 -52.195 -203.835 ;
        RECT -52.525 -205.525 -52.195 -205.195 ;
        RECT -52.525 -208.245 -52.195 -207.915 ;
        RECT -52.52 -209.6 -52.2 -141.96 ;
    END
    PORT
      LAYER met3 ;
        RECT -51.165 129.8 -50.835 130.93 ;
        RECT -51.165 127.675 -50.835 128.005 ;
        RECT -51.165 126.315 -50.835 126.645 ;
        RECT -51.165 124.955 -50.835 125.285 ;
        RECT -51.165 123.595 -50.835 123.925 ;
        RECT -51.165 122.235 -50.835 122.565 ;
        RECT -51.165 120.875 -50.835 121.205 ;
        RECT -51.165 119.515 -50.835 119.845 ;
        RECT -51.165 118.155 -50.835 118.485 ;
        RECT -51.165 116.795 -50.835 117.125 ;
        RECT -51.165 115.435 -50.835 115.765 ;
        RECT -51.165 114.075 -50.835 114.405 ;
        RECT -51.165 112.715 -50.835 113.045 ;
        RECT -51.165 111.355 -50.835 111.685 ;
        RECT -51.165 109.995 -50.835 110.325 ;
        RECT -51.165 108.635 -50.835 108.965 ;
        RECT -51.165 107.275 -50.835 107.605 ;
        RECT -51.165 105.915 -50.835 106.245 ;
        RECT -51.165 104.555 -50.835 104.885 ;
        RECT -51.165 103.195 -50.835 103.525 ;
        RECT -51.165 101.835 -50.835 102.165 ;
        RECT -51.165 100.475 -50.835 100.805 ;
        RECT -51.165 99.115 -50.835 99.445 ;
        RECT -51.165 97.755 -50.835 98.085 ;
        RECT -51.165 96.395 -50.835 96.725 ;
        RECT -51.165 95.035 -50.835 95.365 ;
        RECT -51.165 93.675 -50.835 94.005 ;
        RECT -51.165 92.315 -50.835 92.645 ;
        RECT -51.165 90.955 -50.835 91.285 ;
        RECT -51.165 89.595 -50.835 89.925 ;
        RECT -51.165 88.235 -50.835 88.565 ;
        RECT -51.165 86.875 -50.835 87.205 ;
        RECT -51.165 85.515 -50.835 85.845 ;
        RECT -51.165 84.155 -50.835 84.485 ;
        RECT -51.165 82.795 -50.835 83.125 ;
        RECT -51.165 81.435 -50.835 81.765 ;
        RECT -51.165 80.075 -50.835 80.405 ;
        RECT -51.165 78.715 -50.835 79.045 ;
        RECT -51.165 77.355 -50.835 77.685 ;
        RECT -51.165 75.995 -50.835 76.325 ;
        RECT -51.165 74.635 -50.835 74.965 ;
        RECT -51.165 73.275 -50.835 73.605 ;
        RECT -51.16 73.275 -50.84 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -51.165 48.795 -50.835 49.125 ;
        RECT -51.165 47.435 -50.835 47.765 ;
        RECT -51.165 46.075 -50.835 46.405 ;
        RECT -51.165 44.715 -50.835 45.045 ;
        RECT -51.165 43.355 -50.835 43.685 ;
        RECT -51.165 40.635 -50.835 40.965 ;
        RECT -51.165 39.275 -50.835 39.605 ;
        RECT -51.165 35.195 -50.835 35.525 ;
        RECT -51.165 33.835 -50.835 34.165 ;
        RECT -51.165 32.475 -50.835 32.805 ;
        RECT -51.165 31.115 -50.835 31.445 ;
        RECT -51.165 29.755 -50.835 30.085 ;
        RECT -51.165 28.395 -50.835 28.725 ;
        RECT -51.165 27.035 -50.835 27.365 ;
        RECT -51.165 25.675 -50.835 26.005 ;
        RECT -51.165 24.315 -50.835 24.645 ;
        RECT -51.165 22.955 -50.835 23.285 ;
        RECT -51.165 21.595 -50.835 21.925 ;
        RECT -51.165 20.235 -50.835 20.565 ;
        RECT -51.165 18.875 -50.835 19.205 ;
        RECT -51.165 17.515 -50.835 17.845 ;
        RECT -51.165 16.155 -50.835 16.485 ;
        RECT -51.165 14.795 -50.835 15.125 ;
        RECT -51.165 13.435 -50.835 13.765 ;
        RECT -51.165 12.075 -50.835 12.405 ;
        RECT -51.165 10.715 -50.835 11.045 ;
        RECT -51.165 9.355 -50.835 9.685 ;
        RECT -51.165 7.995 -50.835 8.325 ;
        RECT -51.165 6.635 -50.835 6.965 ;
        RECT -51.165 5.275 -50.835 5.605 ;
        RECT -51.165 3.915 -50.835 4.245 ;
        RECT -51.165 2.555 -50.835 2.885 ;
        RECT -51.165 1.195 -50.835 1.525 ;
        RECT -51.165 -0.165 -50.835 0.165 ;
        RECT -51.165 -1.525 -50.835 -1.195 ;
        RECT -51.165 -2.885 -50.835 -2.555 ;
        RECT -51.165 -4.245 -50.835 -3.915 ;
        RECT -51.165 -5.605 -50.835 -5.275 ;
        RECT -51.165 -6.965 -50.835 -6.635 ;
        RECT -51.165 -8.325 -50.835 -7.995 ;
        RECT -51.165 -9.685 -50.835 -9.355 ;
        RECT -51.165 -11.045 -50.835 -10.715 ;
        RECT -51.165 -12.405 -50.835 -12.075 ;
        RECT -51.165 -13.765 -50.835 -13.435 ;
        RECT -51.165 -15.125 -50.835 -14.795 ;
        RECT -51.165 -16.485 -50.835 -16.155 ;
        RECT -51.165 -17.845 -50.835 -17.515 ;
        RECT -51.165 -19.205 -50.835 -18.875 ;
        RECT -51.165 -20.565 -50.835 -20.235 ;
        RECT -51.165 -21.925 -50.835 -21.595 ;
        RECT -51.165 -23.285 -50.835 -22.955 ;
        RECT -51.165 -24.645 -50.835 -24.315 ;
        RECT -51.165 -26.005 -50.835 -25.675 ;
        RECT -51.165 -27.365 -50.835 -27.035 ;
        RECT -51.165 -28.725 -50.835 -28.395 ;
        RECT -51.165 -30.085 -50.835 -29.755 ;
        RECT -51.165 -31.445 -50.835 -31.115 ;
        RECT -51.165 -32.805 -50.835 -32.475 ;
        RECT -51.165 -34.165 -50.835 -33.835 ;
        RECT -51.165 -35.525 -50.835 -35.195 ;
        RECT -51.165 -36.885 -50.835 -36.555 ;
        RECT -51.165 -39.605 -50.835 -39.275 ;
        RECT -51.165 -40.965 -50.835 -40.635 ;
        RECT -51.165 -42.325 -50.835 -41.995 ;
        RECT -51.165 -43.685 -50.835 -43.355 ;
        RECT -51.165 -45.045 -50.835 -44.715 ;
        RECT -51.165 -46.405 -50.835 -46.075 ;
        RECT -51.165 -47.765 -50.835 -47.435 ;
        RECT -51.165 -49.125 -50.835 -48.795 ;
        RECT -51.165 -50.485 -50.835 -50.155 ;
        RECT -51.165 -51.845 -50.835 -51.515 ;
        RECT -51.165 -53.205 -50.835 -52.875 ;
        RECT -51.165 -54.565 -50.835 -54.235 ;
        RECT -51.165 -55.925 -50.835 -55.595 ;
        RECT -51.165 -57.285 -50.835 -56.955 ;
        RECT -51.165 -58.645 -50.835 -58.315 ;
        RECT -51.165 -60.005 -50.835 -59.675 ;
        RECT -51.165 -61.365 -50.835 -61.035 ;
        RECT -51.165 -62.725 -50.835 -62.395 ;
        RECT -51.165 -64.085 -50.835 -63.755 ;
        RECT -51.165 -65.445 -50.835 -65.115 ;
        RECT -51.165 -66.805 -50.835 -66.475 ;
        RECT -51.165 -68.165 -50.835 -67.835 ;
        RECT -51.165 -69.525 -50.835 -69.195 ;
        RECT -51.165 -70.885 -50.835 -70.555 ;
        RECT -51.165 -72.245 -50.835 -71.915 ;
        RECT -51.165 -73.605 -50.835 -73.275 ;
        RECT -51.165 -74.965 -50.835 -74.635 ;
        RECT -51.165 -76.325 -50.835 -75.995 ;
        RECT -51.165 -77.685 -50.835 -77.355 ;
        RECT -51.165 -79.045 -50.835 -78.715 ;
        RECT -51.165 -80.405 -50.835 -80.075 ;
        RECT -51.165 -81.765 -50.835 -81.435 ;
        RECT -51.165 -83.125 -50.835 -82.795 ;
        RECT -51.165 -84.485 -50.835 -84.155 ;
        RECT -51.165 -85.845 -50.835 -85.515 ;
        RECT -51.165 -87.205 -50.835 -86.875 ;
        RECT -51.165 -88.565 -50.835 -88.235 ;
        RECT -51.165 -89.925 -50.835 -89.595 ;
        RECT -51.165 -91.285 -50.835 -90.955 ;
        RECT -51.165 -92.645 -50.835 -92.315 ;
        RECT -51.165 -94.005 -50.835 -93.675 ;
        RECT -51.165 -95.365 -50.835 -95.035 ;
        RECT -51.165 -96.725 -50.835 -96.395 ;
        RECT -51.165 -98.085 -50.835 -97.755 ;
        RECT -51.165 -99.445 -50.835 -99.115 ;
        RECT -51.165 -100.805 -50.835 -100.475 ;
        RECT -51.165 -102.165 -50.835 -101.835 ;
        RECT -51.165 -103.525 -50.835 -103.195 ;
        RECT -51.165 -104.885 -50.835 -104.555 ;
        RECT -51.165 -106.245 -50.835 -105.915 ;
        RECT -51.165 -107.605 -50.835 -107.275 ;
        RECT -51.165 -108.965 -50.835 -108.635 ;
        RECT -51.165 -110.325 -50.835 -109.995 ;
        RECT -51.165 -113.045 -50.835 -112.715 ;
        RECT -51.165 -114.405 -50.835 -114.075 ;
        RECT -51.165 -115.765 -50.835 -115.435 ;
        RECT -51.165 -117.125 -50.835 -116.795 ;
        RECT -51.165 -118.485 -50.835 -118.155 ;
        RECT -51.165 -119.79 -50.835 -119.46 ;
        RECT -51.165 -121.205 -50.835 -120.875 ;
        RECT -51.165 -122.565 -50.835 -122.235 ;
        RECT -51.165 -123.925 -50.835 -123.595 ;
        RECT -51.165 -126.645 -50.835 -126.315 ;
        RECT -51.165 -128.43 -50.835 -128.1 ;
        RECT -51.165 -129.365 -50.835 -129.035 ;
        RECT -51.165 -130.725 -50.835 -130.395 ;
        RECT -51.165 -133.445 -50.835 -133.115 ;
        RECT -51.165 -134.805 -50.835 -134.475 ;
        RECT -51.165 -136.165 -50.835 -135.835 ;
        RECT -51.165 -137.525 -50.835 -137.195 ;
        RECT -51.165 -138.885 -50.835 -138.555 ;
        RECT -51.165 -140.245 -50.835 -139.915 ;
        RECT -51.165 -142.965 -50.835 -142.635 ;
        RECT -51.165 -144.325 -50.835 -143.995 ;
        RECT -51.165 -145.685 -50.835 -145.355 ;
        RECT -51.165 -147.045 -50.835 -146.715 ;
        RECT -51.165 -148.405 -50.835 -148.075 ;
        RECT -51.165 -149.765 -50.835 -149.435 ;
        RECT -51.165 -151.125 -50.835 -150.795 ;
        RECT -51.165 -152.485 -50.835 -152.155 ;
        RECT -51.165 -153.845 -50.835 -153.515 ;
        RECT -51.165 -155.205 -50.835 -154.875 ;
        RECT -51.165 -156.565 -50.835 -156.235 ;
        RECT -51.165 -157.925 -50.835 -157.595 ;
        RECT -51.165 -159.285 -50.835 -158.955 ;
        RECT -51.165 -160.645 -50.835 -160.315 ;
        RECT -51.165 -162.005 -50.835 -161.675 ;
        RECT -51.165 -163.365 -50.835 -163.035 ;
        RECT -51.165 -164.725 -50.835 -164.395 ;
        RECT -51.165 -166.085 -50.835 -165.755 ;
        RECT -51.165 -167.445 -50.835 -167.115 ;
        RECT -51.165 -168.805 -50.835 -168.475 ;
        RECT -51.165 -170.165 -50.835 -169.835 ;
        RECT -51.165 -171.525 -50.835 -171.195 ;
        RECT -51.165 -172.885 -50.835 -172.555 ;
        RECT -51.165 -174.245 -50.835 -173.915 ;
        RECT -51.165 -175.605 -50.835 -175.275 ;
        RECT -51.165 -176.965 -50.835 -176.635 ;
        RECT -51.165 -178.325 -50.835 -177.995 ;
        RECT -51.165 -179.685 -50.835 -179.355 ;
        RECT -51.165 -181.045 -50.835 -180.715 ;
        RECT -51.165 -182.405 -50.835 -182.075 ;
        RECT -51.165 -183.765 -50.835 -183.435 ;
        RECT -51.165 -185.125 -50.835 -184.795 ;
        RECT -51.165 -186.485 -50.835 -186.155 ;
        RECT -51.165 -187.845 -50.835 -187.515 ;
        RECT -51.165 -189.205 -50.835 -188.875 ;
        RECT -51.165 -190.565 -50.835 -190.235 ;
        RECT -51.165 -191.925 -50.835 -191.595 ;
        RECT -51.165 -193.285 -50.835 -192.955 ;
        RECT -51.165 -194.645 -50.835 -194.315 ;
        RECT -51.165 -196.005 -50.835 -195.675 ;
        RECT -51.165 -197.365 -50.835 -197.035 ;
        RECT -51.165 -198.725 -50.835 -198.395 ;
        RECT -51.165 -200.085 -50.835 -199.755 ;
        RECT -51.165 -201.445 -50.835 -201.115 ;
        RECT -51.165 -202.805 -50.835 -202.475 ;
        RECT -51.165 -204.165 -50.835 -203.835 ;
        RECT -51.165 -205.525 -50.835 -205.195 ;
        RECT -51.165 -208.245 -50.835 -207.915 ;
        RECT -51.165 -210.965 -50.835 -210.635 ;
        RECT -51.165 -212.325 -50.835 -211.995 ;
        RECT -51.165 -213.625 -50.835 -213.295 ;
        RECT -51.165 -215.045 -50.835 -214.715 ;
        RECT -51.165 -216.405 -50.835 -216.075 ;
        RECT -51.165 -217.765 -50.835 -217.435 ;
        RECT -51.165 -219.125 -50.835 -218.795 ;
        RECT -51.165 -221.37 -50.835 -220.24 ;
        RECT -51.16 -221.485 -50.84 49.125 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.805 129.8 -49.475 130.93 ;
        RECT -49.805 127.675 -49.475 128.005 ;
        RECT -49.805 126.315 -49.475 126.645 ;
        RECT -49.805 124.955 -49.475 125.285 ;
        RECT -49.805 123.595 -49.475 123.925 ;
        RECT -49.805 122.235 -49.475 122.565 ;
        RECT -49.805 120.875 -49.475 121.205 ;
        RECT -49.805 119.515 -49.475 119.845 ;
        RECT -49.805 118.155 -49.475 118.485 ;
        RECT -49.805 116.795 -49.475 117.125 ;
        RECT -49.805 115.435 -49.475 115.765 ;
        RECT -49.805 114.075 -49.475 114.405 ;
        RECT -49.805 112.715 -49.475 113.045 ;
        RECT -49.805 111.355 -49.475 111.685 ;
        RECT -49.805 109.995 -49.475 110.325 ;
        RECT -49.805 108.635 -49.475 108.965 ;
        RECT -49.805 107.275 -49.475 107.605 ;
        RECT -49.805 105.915 -49.475 106.245 ;
        RECT -49.805 104.555 -49.475 104.885 ;
        RECT -49.805 103.195 -49.475 103.525 ;
        RECT -49.805 101.835 -49.475 102.165 ;
        RECT -49.805 100.475 -49.475 100.805 ;
        RECT -49.805 99.115 -49.475 99.445 ;
        RECT -49.805 97.755 -49.475 98.085 ;
        RECT -49.805 96.395 -49.475 96.725 ;
        RECT -49.805 95.035 -49.475 95.365 ;
        RECT -49.805 93.675 -49.475 94.005 ;
        RECT -49.805 92.315 -49.475 92.645 ;
        RECT -49.805 90.955 -49.475 91.285 ;
        RECT -49.805 89.595 -49.475 89.925 ;
        RECT -49.805 88.235 -49.475 88.565 ;
        RECT -49.805 86.875 -49.475 87.205 ;
        RECT -49.805 85.515 -49.475 85.845 ;
        RECT -49.805 84.155 -49.475 84.485 ;
        RECT -49.805 82.795 -49.475 83.125 ;
        RECT -49.805 81.435 -49.475 81.765 ;
        RECT -49.805 80.075 -49.475 80.405 ;
        RECT -49.805 78.715 -49.475 79.045 ;
        RECT -49.805 77.355 -49.475 77.685 ;
        RECT -49.805 75.995 -49.475 76.325 ;
        RECT -49.805 74.635 -49.475 74.965 ;
        RECT -49.805 73.275 -49.475 73.605 ;
        RECT -49.8 73.275 -49.48 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.805 48.795 -49.475 49.125 ;
        RECT -49.805 47.435 -49.475 47.765 ;
        RECT -49.805 46.075 -49.475 46.405 ;
        RECT -49.805 44.715 -49.475 45.045 ;
        RECT -49.805 43.355 -49.475 43.685 ;
        RECT -49.805 40.635 -49.475 40.965 ;
        RECT -49.805 39.275 -49.475 39.605 ;
        RECT -49.805 35.195 -49.475 35.525 ;
        RECT -49.805 33.835 -49.475 34.165 ;
        RECT -49.805 32.475 -49.475 32.805 ;
        RECT -49.805 31.115 -49.475 31.445 ;
        RECT -49.805 29.755 -49.475 30.085 ;
        RECT -49.805 28.395 -49.475 28.725 ;
        RECT -49.805 27.035 -49.475 27.365 ;
        RECT -49.805 25.675 -49.475 26.005 ;
        RECT -49.805 24.315 -49.475 24.645 ;
        RECT -49.805 22.955 -49.475 23.285 ;
        RECT -49.805 21.595 -49.475 21.925 ;
        RECT -49.805 20.235 -49.475 20.565 ;
        RECT -49.805 18.875 -49.475 19.205 ;
        RECT -49.805 17.515 -49.475 17.845 ;
        RECT -49.805 16.155 -49.475 16.485 ;
        RECT -49.805 14.795 -49.475 15.125 ;
        RECT -49.805 13.435 -49.475 13.765 ;
        RECT -49.805 12.075 -49.475 12.405 ;
        RECT -49.805 10.715 -49.475 11.045 ;
        RECT -49.805 9.355 -49.475 9.685 ;
        RECT -49.805 7.995 -49.475 8.325 ;
        RECT -49.805 6.635 -49.475 6.965 ;
        RECT -49.805 5.275 -49.475 5.605 ;
        RECT -49.805 3.915 -49.475 4.245 ;
        RECT -49.805 2.555 -49.475 2.885 ;
        RECT -49.805 1.195 -49.475 1.525 ;
        RECT -49.805 -0.165 -49.475 0.165 ;
        RECT -49.805 -1.525 -49.475 -1.195 ;
        RECT -49.805 -2.885 -49.475 -2.555 ;
        RECT -49.805 -4.245 -49.475 -3.915 ;
        RECT -49.805 -5.605 -49.475 -5.275 ;
        RECT -49.805 -6.965 -49.475 -6.635 ;
        RECT -49.805 -8.325 -49.475 -7.995 ;
        RECT -49.805 -9.685 -49.475 -9.355 ;
        RECT -49.805 -11.045 -49.475 -10.715 ;
        RECT -49.805 -12.405 -49.475 -12.075 ;
        RECT -49.805 -13.765 -49.475 -13.435 ;
        RECT -49.805 -15.125 -49.475 -14.795 ;
        RECT -49.805 -16.485 -49.475 -16.155 ;
        RECT -49.805 -17.845 -49.475 -17.515 ;
        RECT -49.805 -19.205 -49.475 -18.875 ;
        RECT -49.805 -20.565 -49.475 -20.235 ;
        RECT -49.805 -21.925 -49.475 -21.595 ;
        RECT -49.805 -23.285 -49.475 -22.955 ;
        RECT -49.805 -24.645 -49.475 -24.315 ;
        RECT -49.805 -26.005 -49.475 -25.675 ;
        RECT -49.805 -27.365 -49.475 -27.035 ;
        RECT -49.805 -28.725 -49.475 -28.395 ;
        RECT -49.805 -30.085 -49.475 -29.755 ;
        RECT -49.805 -31.445 -49.475 -31.115 ;
        RECT -49.805 -32.805 -49.475 -32.475 ;
        RECT -49.805 -34.165 -49.475 -33.835 ;
        RECT -49.805 -35.525 -49.475 -35.195 ;
        RECT -49.805 -36.885 -49.475 -36.555 ;
        RECT -49.805 -39.605 -49.475 -39.275 ;
        RECT -49.805 -40.965 -49.475 -40.635 ;
        RECT -49.805 -42.325 -49.475 -41.995 ;
        RECT -49.805 -43.685 -49.475 -43.355 ;
        RECT -49.805 -45.045 -49.475 -44.715 ;
        RECT -49.805 -46.405 -49.475 -46.075 ;
        RECT -49.805 -47.765 -49.475 -47.435 ;
        RECT -49.805 -49.125 -49.475 -48.795 ;
        RECT -49.805 -50.485 -49.475 -50.155 ;
        RECT -49.805 -51.845 -49.475 -51.515 ;
        RECT -49.805 -53.205 -49.475 -52.875 ;
        RECT -49.805 -54.565 -49.475 -54.235 ;
        RECT -49.805 -55.925 -49.475 -55.595 ;
        RECT -49.805 -57.285 -49.475 -56.955 ;
        RECT -49.805 -58.645 -49.475 -58.315 ;
        RECT -49.805 -60.005 -49.475 -59.675 ;
        RECT -49.805 -61.365 -49.475 -61.035 ;
        RECT -49.805 -62.725 -49.475 -62.395 ;
        RECT -49.805 -64.085 -49.475 -63.755 ;
        RECT -49.805 -65.445 -49.475 -65.115 ;
        RECT -49.805 -66.805 -49.475 -66.475 ;
        RECT -49.805 -68.165 -49.475 -67.835 ;
        RECT -49.805 -69.525 -49.475 -69.195 ;
        RECT -49.805 -70.885 -49.475 -70.555 ;
        RECT -49.805 -72.245 -49.475 -71.915 ;
        RECT -49.805 -73.605 -49.475 -73.275 ;
        RECT -49.805 -74.965 -49.475 -74.635 ;
        RECT -49.805 -76.325 -49.475 -75.995 ;
        RECT -49.805 -77.685 -49.475 -77.355 ;
        RECT -49.805 -79.045 -49.475 -78.715 ;
        RECT -49.805 -80.405 -49.475 -80.075 ;
        RECT -49.805 -81.765 -49.475 -81.435 ;
        RECT -49.805 -83.125 -49.475 -82.795 ;
        RECT -49.805 -84.485 -49.475 -84.155 ;
        RECT -49.805 -85.845 -49.475 -85.515 ;
        RECT -49.805 -87.205 -49.475 -86.875 ;
        RECT -49.805 -88.565 -49.475 -88.235 ;
        RECT -49.805 -89.925 -49.475 -89.595 ;
        RECT -49.805 -91.285 -49.475 -90.955 ;
        RECT -49.805 -92.645 -49.475 -92.315 ;
        RECT -49.805 -94.005 -49.475 -93.675 ;
        RECT -49.805 -95.365 -49.475 -95.035 ;
        RECT -49.805 -96.725 -49.475 -96.395 ;
        RECT -49.805 -98.085 -49.475 -97.755 ;
        RECT -49.805 -99.445 -49.475 -99.115 ;
        RECT -49.805 -100.805 -49.475 -100.475 ;
        RECT -49.805 -102.165 -49.475 -101.835 ;
        RECT -49.805 -103.525 -49.475 -103.195 ;
        RECT -49.805 -104.885 -49.475 -104.555 ;
        RECT -49.805 -106.245 -49.475 -105.915 ;
        RECT -49.805 -107.605 -49.475 -107.275 ;
        RECT -49.805 -108.965 -49.475 -108.635 ;
        RECT -49.805 -110.325 -49.475 -109.995 ;
        RECT -49.805 -113.045 -49.475 -112.715 ;
        RECT -49.805 -114.405 -49.475 -114.075 ;
        RECT -49.805 -115.765 -49.475 -115.435 ;
        RECT -49.805 -117.125 -49.475 -116.795 ;
        RECT -49.805 -118.485 -49.475 -118.155 ;
        RECT -49.805 -119.79 -49.475 -119.46 ;
        RECT -49.805 -121.205 -49.475 -120.875 ;
        RECT -49.805 -122.565 -49.475 -122.235 ;
        RECT -49.805 -123.925 -49.475 -123.595 ;
        RECT -49.805 -126.645 -49.475 -126.315 ;
        RECT -49.805 -128.43 -49.475 -128.1 ;
        RECT -49.805 -129.365 -49.475 -129.035 ;
        RECT -49.805 -130.725 -49.475 -130.395 ;
        RECT -49.805 -133.445 -49.475 -133.115 ;
        RECT -49.805 -134.805 -49.475 -134.475 ;
        RECT -49.805 -136.165 -49.475 -135.835 ;
        RECT -49.805 -137.525 -49.475 -137.195 ;
        RECT -49.805 -138.885 -49.475 -138.555 ;
        RECT -49.805 -140.245 -49.475 -139.915 ;
        RECT -49.805 -142.965 -49.475 -142.635 ;
        RECT -49.805 -144.325 -49.475 -143.995 ;
        RECT -49.805 -145.685 -49.475 -145.355 ;
        RECT -49.805 -147.045 -49.475 -146.715 ;
        RECT -49.805 -148.405 -49.475 -148.075 ;
        RECT -49.805 -149.765 -49.475 -149.435 ;
        RECT -49.805 -151.125 -49.475 -150.795 ;
        RECT -49.805 -152.485 -49.475 -152.155 ;
        RECT -49.805 -153.845 -49.475 -153.515 ;
        RECT -49.805 -155.205 -49.475 -154.875 ;
        RECT -49.805 -156.565 -49.475 -156.235 ;
        RECT -49.805 -157.925 -49.475 -157.595 ;
        RECT -49.805 -159.285 -49.475 -158.955 ;
        RECT -49.805 -160.645 -49.475 -160.315 ;
        RECT -49.805 -162.005 -49.475 -161.675 ;
        RECT -49.805 -163.365 -49.475 -163.035 ;
        RECT -49.805 -164.725 -49.475 -164.395 ;
        RECT -49.805 -166.085 -49.475 -165.755 ;
        RECT -49.805 -167.445 -49.475 -167.115 ;
        RECT -49.805 -168.805 -49.475 -168.475 ;
        RECT -49.805 -170.165 -49.475 -169.835 ;
        RECT -49.805 -171.525 -49.475 -171.195 ;
        RECT -49.805 -172.885 -49.475 -172.555 ;
        RECT -49.805 -174.245 -49.475 -173.915 ;
        RECT -49.805 -175.605 -49.475 -175.275 ;
        RECT -49.805 -176.965 -49.475 -176.635 ;
        RECT -49.805 -178.325 -49.475 -177.995 ;
        RECT -49.805 -179.685 -49.475 -179.355 ;
        RECT -49.805 -181.045 -49.475 -180.715 ;
        RECT -49.805 -182.405 -49.475 -182.075 ;
        RECT -49.805 -183.765 -49.475 -183.435 ;
        RECT -49.805 -185.125 -49.475 -184.795 ;
        RECT -49.805 -186.485 -49.475 -186.155 ;
        RECT -49.805 -187.845 -49.475 -187.515 ;
        RECT -49.805 -189.205 -49.475 -188.875 ;
        RECT -49.805 -190.565 -49.475 -190.235 ;
        RECT -49.805 -191.925 -49.475 -191.595 ;
        RECT -49.805 -193.285 -49.475 -192.955 ;
        RECT -49.805 -194.645 -49.475 -194.315 ;
        RECT -49.805 -196.005 -49.475 -195.675 ;
        RECT -49.805 -197.365 -49.475 -197.035 ;
        RECT -49.805 -198.725 -49.475 -198.395 ;
        RECT -49.805 -200.085 -49.475 -199.755 ;
        RECT -49.805 -201.445 -49.475 -201.115 ;
        RECT -49.805 -202.805 -49.475 -202.475 ;
        RECT -49.805 -204.165 -49.475 -203.835 ;
        RECT -49.805 -205.525 -49.475 -205.195 ;
        RECT -49.805 -208.245 -49.475 -207.915 ;
        RECT -49.805 -210.965 -49.475 -210.635 ;
        RECT -49.805 -212.325 -49.475 -211.995 ;
        RECT -49.805 -213.625 -49.475 -213.295 ;
        RECT -49.805 -215.045 -49.475 -214.715 ;
        RECT -49.805 -216.405 -49.475 -216.075 ;
        RECT -49.805 -217.765 -49.475 -217.435 ;
        RECT -49.805 -219.125 -49.475 -218.795 ;
        RECT -49.805 -221.37 -49.475 -220.24 ;
        RECT -49.8 -221.485 -49.48 49.125 ;
    END
    PORT
      LAYER met3 ;
        RECT -48.445 129.8 -48.115 130.93 ;
        RECT -48.445 127.675 -48.115 128.005 ;
        RECT -48.445 126.315 -48.115 126.645 ;
        RECT -48.445 124.955 -48.115 125.285 ;
        RECT -48.445 123.595 -48.115 123.925 ;
        RECT -48.445 122.235 -48.115 122.565 ;
        RECT -48.445 120.875 -48.115 121.205 ;
        RECT -48.445 119.515 -48.115 119.845 ;
        RECT -48.445 118.155 -48.115 118.485 ;
        RECT -48.445 116.795 -48.115 117.125 ;
        RECT -48.445 115.435 -48.115 115.765 ;
        RECT -48.445 114.075 -48.115 114.405 ;
        RECT -48.445 112.715 -48.115 113.045 ;
        RECT -48.445 111.355 -48.115 111.685 ;
        RECT -48.445 109.995 -48.115 110.325 ;
        RECT -48.445 108.635 -48.115 108.965 ;
        RECT -48.445 107.275 -48.115 107.605 ;
        RECT -48.445 105.915 -48.115 106.245 ;
        RECT -48.445 104.555 -48.115 104.885 ;
        RECT -48.445 103.195 -48.115 103.525 ;
        RECT -48.445 101.835 -48.115 102.165 ;
        RECT -48.445 100.475 -48.115 100.805 ;
        RECT -48.445 99.115 -48.115 99.445 ;
        RECT -48.445 97.755 -48.115 98.085 ;
        RECT -48.445 96.395 -48.115 96.725 ;
        RECT -48.445 95.035 -48.115 95.365 ;
        RECT -48.445 93.675 -48.115 94.005 ;
        RECT -48.445 92.315 -48.115 92.645 ;
        RECT -48.445 90.955 -48.115 91.285 ;
        RECT -48.445 89.595 -48.115 89.925 ;
        RECT -48.445 88.235 -48.115 88.565 ;
        RECT -48.445 86.875 -48.115 87.205 ;
        RECT -48.445 85.515 -48.115 85.845 ;
        RECT -48.445 84.155 -48.115 84.485 ;
        RECT -48.445 82.795 -48.115 83.125 ;
        RECT -48.445 81.435 -48.115 81.765 ;
        RECT -48.445 80.075 -48.115 80.405 ;
        RECT -48.445 78.715 -48.115 79.045 ;
        RECT -48.445 77.355 -48.115 77.685 ;
        RECT -48.445 75.995 -48.115 76.325 ;
        RECT -48.445 74.635 -48.115 74.965 ;
        RECT -48.445 73.275 -48.115 73.605 ;
        RECT -48.44 73.275 -48.12 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -48.445 48.795 -48.115 49.125 ;
        RECT -48.445 47.435 -48.115 47.765 ;
        RECT -48.445 46.075 -48.115 46.405 ;
        RECT -48.445 44.715 -48.115 45.045 ;
        RECT -48.445 43.355 -48.115 43.685 ;
        RECT -48.445 40.635 -48.115 40.965 ;
        RECT -48.445 39.275 -48.115 39.605 ;
        RECT -48.445 35.195 -48.115 35.525 ;
        RECT -48.445 33.835 -48.115 34.165 ;
        RECT -48.445 32.475 -48.115 32.805 ;
        RECT -48.445 31.115 -48.115 31.445 ;
        RECT -48.445 29.755 -48.115 30.085 ;
        RECT -48.445 28.395 -48.115 28.725 ;
        RECT -48.445 27.035 -48.115 27.365 ;
        RECT -48.445 25.675 -48.115 26.005 ;
        RECT -48.445 24.315 -48.115 24.645 ;
        RECT -48.445 22.955 -48.115 23.285 ;
        RECT -48.445 21.595 -48.115 21.925 ;
        RECT -48.445 20.235 -48.115 20.565 ;
        RECT -48.445 18.875 -48.115 19.205 ;
        RECT -48.445 17.515 -48.115 17.845 ;
        RECT -48.445 16.155 -48.115 16.485 ;
        RECT -48.445 14.795 -48.115 15.125 ;
        RECT -48.445 13.435 -48.115 13.765 ;
        RECT -48.445 12.075 -48.115 12.405 ;
        RECT -48.445 10.715 -48.115 11.045 ;
        RECT -48.445 9.355 -48.115 9.685 ;
        RECT -48.445 7.995 -48.115 8.325 ;
        RECT -48.445 6.635 -48.115 6.965 ;
        RECT -48.445 5.275 -48.115 5.605 ;
        RECT -48.445 3.915 -48.115 4.245 ;
        RECT -48.445 2.555 -48.115 2.885 ;
        RECT -48.445 1.195 -48.115 1.525 ;
        RECT -48.445 -0.165 -48.115 0.165 ;
        RECT -48.445 -1.525 -48.115 -1.195 ;
        RECT -48.445 -2.885 -48.115 -2.555 ;
        RECT -48.445 -4.245 -48.115 -3.915 ;
        RECT -48.445 -5.605 -48.115 -5.275 ;
        RECT -48.445 -6.965 -48.115 -6.635 ;
        RECT -48.445 -8.325 -48.115 -7.995 ;
        RECT -48.445 -9.685 -48.115 -9.355 ;
        RECT -48.445 -11.045 -48.115 -10.715 ;
        RECT -48.445 -12.405 -48.115 -12.075 ;
        RECT -48.445 -13.765 -48.115 -13.435 ;
        RECT -48.445 -15.125 -48.115 -14.795 ;
        RECT -48.445 -16.485 -48.115 -16.155 ;
        RECT -48.445 -17.845 -48.115 -17.515 ;
        RECT -48.445 -19.205 -48.115 -18.875 ;
        RECT -48.445 -20.565 -48.115 -20.235 ;
        RECT -48.445 -21.925 -48.115 -21.595 ;
        RECT -48.445 -23.285 -48.115 -22.955 ;
        RECT -48.445 -24.645 -48.115 -24.315 ;
        RECT -48.445 -26.005 -48.115 -25.675 ;
        RECT -48.445 -27.365 -48.115 -27.035 ;
        RECT -48.445 -28.725 -48.115 -28.395 ;
        RECT -48.445 -30.085 -48.115 -29.755 ;
        RECT -48.445 -31.445 -48.115 -31.115 ;
        RECT -48.445 -32.805 -48.115 -32.475 ;
        RECT -48.445 -35.525 -48.115 -35.195 ;
        RECT -48.445 -36.885 -48.115 -36.555 ;
        RECT -48.445 -39.605 -48.115 -39.275 ;
        RECT -48.445 -40.965 -48.115 -40.635 ;
        RECT -48.445 -42.325 -48.115 -41.995 ;
        RECT -48.445 -43.685 -48.115 -43.355 ;
        RECT -48.445 -45.045 -48.115 -44.715 ;
        RECT -48.445 -46.405 -48.115 -46.075 ;
        RECT -48.445 -47.765 -48.115 -47.435 ;
        RECT -48.445 -49.125 -48.115 -48.795 ;
        RECT -48.445 -50.485 -48.115 -50.155 ;
        RECT -48.445 -51.845 -48.115 -51.515 ;
        RECT -48.445 -53.205 -48.115 -52.875 ;
        RECT -48.445 -54.565 -48.115 -54.235 ;
        RECT -48.445 -55.925 -48.115 -55.595 ;
        RECT -48.445 -57.285 -48.115 -56.955 ;
        RECT -48.445 -58.645 -48.115 -58.315 ;
        RECT -48.445 -60.005 -48.115 -59.675 ;
        RECT -48.445 -61.365 -48.115 -61.035 ;
        RECT -48.445 -62.725 -48.115 -62.395 ;
        RECT -48.445 -64.085 -48.115 -63.755 ;
        RECT -48.445 -65.445 -48.115 -65.115 ;
        RECT -48.445 -66.805 -48.115 -66.475 ;
        RECT -48.445 -68.165 -48.115 -67.835 ;
        RECT -48.445 -69.525 -48.115 -69.195 ;
        RECT -48.445 -70.885 -48.115 -70.555 ;
        RECT -48.445 -72.245 -48.115 -71.915 ;
        RECT -48.445 -73.605 -48.115 -73.275 ;
        RECT -48.445 -74.965 -48.115 -74.635 ;
        RECT -48.445 -76.325 -48.115 -75.995 ;
        RECT -48.445 -77.685 -48.115 -77.355 ;
        RECT -48.445 -79.045 -48.115 -78.715 ;
        RECT -48.445 -80.405 -48.115 -80.075 ;
        RECT -48.445 -81.765 -48.115 -81.435 ;
        RECT -48.445 -83.125 -48.115 -82.795 ;
        RECT -48.445 -84.485 -48.115 -84.155 ;
        RECT -48.445 -85.845 -48.115 -85.515 ;
        RECT -48.445 -87.205 -48.115 -86.875 ;
        RECT -48.445 -88.565 -48.115 -88.235 ;
        RECT -48.445 -89.925 -48.115 -89.595 ;
        RECT -48.445 -91.285 -48.115 -90.955 ;
        RECT -48.445 -92.645 -48.115 -92.315 ;
        RECT -48.445 -94.005 -48.115 -93.675 ;
        RECT -48.445 -95.365 -48.115 -95.035 ;
        RECT -48.445 -96.725 -48.115 -96.395 ;
        RECT -48.445 -98.085 -48.115 -97.755 ;
        RECT -48.445 -99.445 -48.115 -99.115 ;
        RECT -48.445 -100.805 -48.115 -100.475 ;
        RECT -48.445 -102.165 -48.115 -101.835 ;
        RECT -48.445 -103.525 -48.115 -103.195 ;
        RECT -48.445 -104.885 -48.115 -104.555 ;
        RECT -48.445 -106.245 -48.115 -105.915 ;
        RECT -48.445 -107.605 -48.115 -107.275 ;
        RECT -48.445 -108.965 -48.115 -108.635 ;
        RECT -48.445 -110.325 -48.115 -109.995 ;
        RECT -48.445 -113.045 -48.115 -112.715 ;
        RECT -48.445 -114.405 -48.115 -114.075 ;
        RECT -48.445 -115.765 -48.115 -115.435 ;
        RECT -48.445 -117.125 -48.115 -116.795 ;
        RECT -48.445 -118.485 -48.115 -118.155 ;
        RECT -48.445 -119.79 -48.115 -119.46 ;
        RECT -48.445 -121.205 -48.115 -120.875 ;
        RECT -48.445 -122.565 -48.115 -122.235 ;
        RECT -48.445 -123.925 -48.115 -123.595 ;
        RECT -48.445 -126.645 -48.115 -126.315 ;
        RECT -48.445 -128.43 -48.115 -128.1 ;
        RECT -48.445 -129.365 -48.115 -129.035 ;
        RECT -48.445 -130.725 -48.115 -130.395 ;
        RECT -48.44 -132.76 -48.12 49.125 ;
    END
    PORT
      LAYER met3 ;
        RECT -48.445 -212.325 -48.115 -211.995 ;
        RECT -48.445 -213.625 -48.115 -213.295 ;
        RECT -48.445 -215.045 -48.115 -214.715 ;
        RECT -48.445 -216.405 -48.115 -216.075 ;
        RECT -48.445 -217.765 -48.115 -217.435 ;
        RECT -48.445 -219.125 -48.115 -218.795 ;
        RECT -48.445 -221.37 -48.115 -220.24 ;
        RECT -48.44 -221.485 -48.12 -211.995 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.085 129.8 -46.755 130.93 ;
        RECT -47.085 127.675 -46.755 128.005 ;
        RECT -47.085 126.315 -46.755 126.645 ;
        RECT -47.085 124.955 -46.755 125.285 ;
        RECT -47.085 123.595 -46.755 123.925 ;
        RECT -47.085 122.235 -46.755 122.565 ;
        RECT -47.085 120.875 -46.755 121.205 ;
        RECT -47.085 119.515 -46.755 119.845 ;
        RECT -47.085 118.155 -46.755 118.485 ;
        RECT -47.085 116.795 -46.755 117.125 ;
        RECT -47.085 115.435 -46.755 115.765 ;
        RECT -47.085 114.075 -46.755 114.405 ;
        RECT -47.085 112.715 -46.755 113.045 ;
        RECT -47.085 111.355 -46.755 111.685 ;
        RECT -47.085 109.995 -46.755 110.325 ;
        RECT -47.085 108.635 -46.755 108.965 ;
        RECT -47.085 107.275 -46.755 107.605 ;
        RECT -47.085 105.915 -46.755 106.245 ;
        RECT -47.085 104.555 -46.755 104.885 ;
        RECT -47.085 103.195 -46.755 103.525 ;
        RECT -47.085 101.835 -46.755 102.165 ;
        RECT -47.085 100.475 -46.755 100.805 ;
        RECT -47.085 99.115 -46.755 99.445 ;
        RECT -47.085 97.755 -46.755 98.085 ;
        RECT -47.085 96.395 -46.755 96.725 ;
        RECT -47.085 95.035 -46.755 95.365 ;
        RECT -47.085 93.675 -46.755 94.005 ;
        RECT -47.085 92.315 -46.755 92.645 ;
        RECT -47.085 90.955 -46.755 91.285 ;
        RECT -47.085 89.595 -46.755 89.925 ;
        RECT -47.085 88.235 -46.755 88.565 ;
        RECT -47.085 86.875 -46.755 87.205 ;
        RECT -47.085 85.515 -46.755 85.845 ;
        RECT -47.085 84.155 -46.755 84.485 ;
        RECT -47.085 82.795 -46.755 83.125 ;
        RECT -47.085 81.435 -46.755 81.765 ;
        RECT -47.085 80.075 -46.755 80.405 ;
        RECT -47.085 78.715 -46.755 79.045 ;
        RECT -47.085 77.355 -46.755 77.685 ;
        RECT -47.085 75.995 -46.755 76.325 ;
        RECT -47.085 74.635 -46.755 74.965 ;
        RECT -47.085 73.275 -46.755 73.605 ;
        RECT -47.08 73.275 -46.76 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.085 -46.405 -46.755 -46.075 ;
        RECT -47.085 -47.765 -46.755 -47.435 ;
        RECT -47.085 -49.125 -46.755 -48.795 ;
        RECT -47.085 -50.485 -46.755 -50.155 ;
        RECT -47.085 -51.845 -46.755 -51.515 ;
        RECT -47.085 -53.205 -46.755 -52.875 ;
        RECT -47.085 -54.565 -46.755 -54.235 ;
        RECT -47.085 -55.925 -46.755 -55.595 ;
        RECT -47.085 -57.285 -46.755 -56.955 ;
        RECT -47.085 -58.645 -46.755 -58.315 ;
        RECT -47.085 -60.005 -46.755 -59.675 ;
        RECT -47.085 -61.365 -46.755 -61.035 ;
        RECT -47.085 -62.725 -46.755 -62.395 ;
        RECT -47.085 -64.085 -46.755 -63.755 ;
        RECT -47.085 -65.445 -46.755 -65.115 ;
        RECT -47.085 -66.805 -46.755 -66.475 ;
        RECT -47.085 -68.165 -46.755 -67.835 ;
        RECT -47.085 -69.525 -46.755 -69.195 ;
        RECT -47.085 -70.885 -46.755 -70.555 ;
        RECT -47.085 -72.245 -46.755 -71.915 ;
        RECT -47.085 -73.605 -46.755 -73.275 ;
        RECT -47.085 -74.965 -46.755 -74.635 ;
        RECT -47.085 -76.325 -46.755 -75.995 ;
        RECT -47.085 -77.685 -46.755 -77.355 ;
        RECT -47.085 -79.045 -46.755 -78.715 ;
        RECT -47.085 -80.405 -46.755 -80.075 ;
        RECT -47.085 -81.765 -46.755 -81.435 ;
        RECT -47.085 -83.125 -46.755 -82.795 ;
        RECT -47.085 -84.485 -46.755 -84.155 ;
        RECT -47.085 -85.845 -46.755 -85.515 ;
        RECT -47.085 -87.205 -46.755 -86.875 ;
        RECT -47.085 -88.565 -46.755 -88.235 ;
        RECT -47.085 -89.925 -46.755 -89.595 ;
        RECT -47.085 -91.285 -46.755 -90.955 ;
        RECT -47.085 -92.645 -46.755 -92.315 ;
        RECT -47.085 -94.005 -46.755 -93.675 ;
        RECT -47.085 -95.365 -46.755 -95.035 ;
        RECT -47.085 -96.725 -46.755 -96.395 ;
        RECT -47.085 -98.085 -46.755 -97.755 ;
        RECT -47.085 -99.445 -46.755 -99.115 ;
        RECT -47.085 -100.805 -46.755 -100.475 ;
        RECT -47.085 -102.165 -46.755 -101.835 ;
        RECT -47.085 -103.525 -46.755 -103.195 ;
        RECT -47.085 -104.885 -46.755 -104.555 ;
        RECT -47.085 -106.245 -46.755 -105.915 ;
        RECT -47.085 -107.605 -46.755 -107.275 ;
        RECT -47.085 -108.965 -46.755 -108.635 ;
        RECT -47.085 -110.325 -46.755 -109.995 ;
        RECT -47.085 -113.045 -46.755 -112.715 ;
        RECT -47.085 -114.405 -46.755 -114.075 ;
        RECT -47.085 -115.765 -46.755 -115.435 ;
        RECT -47.085 -117.125 -46.755 -116.795 ;
        RECT -47.085 -118.485 -46.755 -118.155 ;
        RECT -47.085 -119.79 -46.755 -119.46 ;
        RECT -47.085 -121.205 -46.755 -120.875 ;
        RECT -47.085 -122.565 -46.755 -122.235 ;
        RECT -47.085 -123.925 -46.755 -123.595 ;
        RECT -47.085 -126.645 -46.755 -126.315 ;
        RECT -47.085 -128.43 -46.755 -128.1 ;
        RECT -47.085 -129.365 -46.755 -129.035 ;
        RECT -47.085 -130.725 -46.755 -130.395 ;
        RECT -47.08 -132.08 -46.76 49.125 ;
        RECT -47.085 48.795 -46.755 49.125 ;
        RECT -47.085 47.435 -46.755 47.765 ;
        RECT -47.085 46.075 -46.755 46.405 ;
        RECT -47.085 44.715 -46.755 45.045 ;
        RECT -47.085 43.355 -46.755 43.685 ;
        RECT -47.085 40.635 -46.755 40.965 ;
        RECT -47.085 39.275 -46.755 39.605 ;
        RECT -47.085 35.195 -46.755 35.525 ;
        RECT -47.085 33.835 -46.755 34.165 ;
        RECT -47.085 32.475 -46.755 32.805 ;
        RECT -47.085 31.115 -46.755 31.445 ;
        RECT -47.085 29.755 -46.755 30.085 ;
        RECT -47.085 28.395 -46.755 28.725 ;
        RECT -47.085 27.035 -46.755 27.365 ;
        RECT -47.085 25.675 -46.755 26.005 ;
        RECT -47.085 24.315 -46.755 24.645 ;
        RECT -47.085 22.955 -46.755 23.285 ;
        RECT -47.085 21.595 -46.755 21.925 ;
        RECT -47.085 20.235 -46.755 20.565 ;
        RECT -47.085 18.875 -46.755 19.205 ;
        RECT -47.085 17.515 -46.755 17.845 ;
        RECT -47.085 16.155 -46.755 16.485 ;
        RECT -47.085 14.795 -46.755 15.125 ;
        RECT -47.085 13.435 -46.755 13.765 ;
        RECT -47.085 12.075 -46.755 12.405 ;
        RECT -47.085 10.715 -46.755 11.045 ;
        RECT -47.085 9.355 -46.755 9.685 ;
        RECT -47.085 7.995 -46.755 8.325 ;
        RECT -47.085 6.635 -46.755 6.965 ;
        RECT -47.085 5.275 -46.755 5.605 ;
        RECT -47.085 3.915 -46.755 4.245 ;
        RECT -47.085 2.555 -46.755 2.885 ;
        RECT -47.085 1.195 -46.755 1.525 ;
        RECT -47.085 -0.165 -46.755 0.165 ;
        RECT -47.085 -1.525 -46.755 -1.195 ;
        RECT -47.085 -2.885 -46.755 -2.555 ;
        RECT -47.085 -4.245 -46.755 -3.915 ;
        RECT -47.085 -5.605 -46.755 -5.275 ;
        RECT -47.085 -6.965 -46.755 -6.635 ;
        RECT -47.085 -8.325 -46.755 -7.995 ;
        RECT -47.085 -9.685 -46.755 -9.355 ;
        RECT -47.085 -11.045 -46.755 -10.715 ;
        RECT -47.085 -12.405 -46.755 -12.075 ;
        RECT -47.085 -13.765 -46.755 -13.435 ;
        RECT -47.085 -15.125 -46.755 -14.795 ;
        RECT -47.085 -16.485 -46.755 -16.155 ;
        RECT -47.085 -17.845 -46.755 -17.515 ;
        RECT -47.085 -19.205 -46.755 -18.875 ;
        RECT -47.085 -20.565 -46.755 -20.235 ;
        RECT -47.085 -21.925 -46.755 -21.595 ;
        RECT -47.085 -23.285 -46.755 -22.955 ;
        RECT -47.085 -24.645 -46.755 -24.315 ;
        RECT -47.085 -26.005 -46.755 -25.675 ;
        RECT -47.085 -27.365 -46.755 -27.035 ;
        RECT -47.085 -28.725 -46.755 -28.395 ;
        RECT -47.085 -30.085 -46.755 -29.755 ;
        RECT -47.085 -31.445 -46.755 -31.115 ;
        RECT -47.085 -32.805 -46.755 -32.475 ;
        RECT -47.085 -35.525 -46.755 -35.195 ;
        RECT -47.085 -36.885 -46.755 -36.555 ;
        RECT -47.085 -39.605 -46.755 -39.275 ;
        RECT -47.085 -40.965 -46.755 -40.635 ;
        RECT -47.085 -42.325 -46.755 -41.995 ;
        RECT -47.085 -43.685 -46.755 -43.355 ;
        RECT -47.085 -45.045 -46.755 -44.715 ;
    END
    PORT
      LAYER met3 ;
        RECT -57.965 129.8 -57.635 130.93 ;
        RECT -57.965 127.675 -57.635 128.005 ;
        RECT -57.965 126.315 -57.635 126.645 ;
        RECT -57.965 124.955 -57.635 125.285 ;
        RECT -57.965 123.595 -57.635 123.925 ;
        RECT -57.965 122.235 -57.635 122.565 ;
        RECT -57.965 120.875 -57.635 121.205 ;
        RECT -57.965 119.515 -57.635 119.845 ;
        RECT -57.965 118.155 -57.635 118.485 ;
        RECT -57.965 116.795 -57.635 117.125 ;
        RECT -57.965 115.435 -57.635 115.765 ;
        RECT -57.965 114.075 -57.635 114.405 ;
        RECT -57.965 112.715 -57.635 113.045 ;
        RECT -57.965 111.355 -57.635 111.685 ;
        RECT -57.965 109.995 -57.635 110.325 ;
        RECT -57.965 108.635 -57.635 108.965 ;
        RECT -57.965 107.275 -57.635 107.605 ;
        RECT -57.965 105.915 -57.635 106.245 ;
        RECT -57.965 104.555 -57.635 104.885 ;
        RECT -57.965 103.195 -57.635 103.525 ;
        RECT -57.965 101.835 -57.635 102.165 ;
        RECT -57.965 100.475 -57.635 100.805 ;
        RECT -57.965 99.115 -57.635 99.445 ;
        RECT -57.965 97.755 -57.635 98.085 ;
        RECT -57.965 96.395 -57.635 96.725 ;
        RECT -57.965 95.035 -57.635 95.365 ;
        RECT -57.965 93.675 -57.635 94.005 ;
        RECT -57.965 92.315 -57.635 92.645 ;
        RECT -57.965 90.955 -57.635 91.285 ;
        RECT -57.965 89.595 -57.635 89.925 ;
        RECT -57.965 88.235 -57.635 88.565 ;
        RECT -57.965 86.875 -57.635 87.205 ;
        RECT -57.965 85.515 -57.635 85.845 ;
        RECT -57.965 84.155 -57.635 84.485 ;
        RECT -57.965 82.795 -57.635 83.125 ;
        RECT -57.965 81.435 -57.635 81.765 ;
        RECT -57.965 80.075 -57.635 80.405 ;
        RECT -57.965 78.715 -57.635 79.045 ;
        RECT -57.965 77.355 -57.635 77.685 ;
        RECT -57.965 75.995 -57.635 76.325 ;
        RECT -57.965 74.635 -57.635 74.965 ;
        RECT -57.965 73.275 -57.635 73.605 ;
        RECT -57.965 71.915 -57.635 72.245 ;
        RECT -57.965 70.555 -57.635 70.885 ;
        RECT -57.965 69.195 -57.635 69.525 ;
        RECT -57.965 67.835 -57.635 68.165 ;
        RECT -57.965 66.475 -57.635 66.805 ;
        RECT -57.965 65.115 -57.635 65.445 ;
        RECT -57.965 63.755 -57.635 64.085 ;
        RECT -57.965 62.395 -57.635 62.725 ;
        RECT -57.965 61.035 -57.635 61.365 ;
        RECT -57.965 59.675 -57.635 60.005 ;
        RECT -57.965 58.315 -57.635 58.645 ;
        RECT -57.965 56.955 -57.635 57.285 ;
        RECT -57.965 55.595 -57.635 55.925 ;
        RECT -57.965 54.235 -57.635 54.565 ;
        RECT -57.965 52.875 -57.635 53.205 ;
        RECT -57.965 51.515 -57.635 51.845 ;
        RECT -57.965 50.155 -57.635 50.485 ;
        RECT -57.965 48.795 -57.635 49.125 ;
        RECT -57.965 47.435 -57.635 47.765 ;
        RECT -57.965 46.075 -57.635 46.405 ;
        RECT -57.965 44.715 -57.635 45.045 ;
        RECT -57.965 43.355 -57.635 43.685 ;
        RECT -57.965 41.995 -57.635 42.325 ;
        RECT -57.965 40.635 -57.635 40.965 ;
        RECT -57.965 39.275 -57.635 39.605 ;
        RECT -57.965 37.915 -57.635 38.245 ;
        RECT -57.965 36.555 -57.635 36.885 ;
        RECT -57.965 35.195 -57.635 35.525 ;
        RECT -57.965 33.835 -57.635 34.165 ;
        RECT -57.965 32.475 -57.635 32.805 ;
        RECT -57.965 31.115 -57.635 31.445 ;
        RECT -57.965 29.755 -57.635 30.085 ;
        RECT -57.965 28.395 -57.635 28.725 ;
        RECT -57.965 27.035 -57.635 27.365 ;
        RECT -57.965 25.675 -57.635 26.005 ;
        RECT -57.965 24.315 -57.635 24.645 ;
        RECT -57.965 22.955 -57.635 23.285 ;
        RECT -57.965 21.595 -57.635 21.925 ;
        RECT -57.965 20.235 -57.635 20.565 ;
        RECT -57.965 18.875 -57.635 19.205 ;
        RECT -57.965 17.515 -57.635 17.845 ;
        RECT -57.965 16.155 -57.635 16.485 ;
        RECT -57.965 14.795 -57.635 15.125 ;
        RECT -57.965 13.435 -57.635 13.765 ;
        RECT -57.965 12.075 -57.635 12.405 ;
        RECT -57.965 10.715 -57.635 11.045 ;
        RECT -57.965 9.355 -57.635 9.685 ;
        RECT -57.965 7.995 -57.635 8.325 ;
        RECT -57.965 6.635 -57.635 6.965 ;
        RECT -57.965 5.275 -57.635 5.605 ;
        RECT -57.965 3.915 -57.635 4.245 ;
        RECT -57.965 2.555 -57.635 2.885 ;
        RECT -57.965 1.195 -57.635 1.525 ;
        RECT -57.965 -0.165 -57.635 0.165 ;
        RECT -57.965 -1.525 -57.635 -1.195 ;
        RECT -57.965 -2.885 -57.635 -2.555 ;
        RECT -57.965 -4.245 -57.635 -3.915 ;
        RECT -57.965 -5.605 -57.635 -5.275 ;
        RECT -57.965 -6.965 -57.635 -6.635 ;
        RECT -57.965 -8.325 -57.635 -7.995 ;
        RECT -57.965 -9.685 -57.635 -9.355 ;
        RECT -57.965 -11.045 -57.635 -10.715 ;
        RECT -57.965 -12.405 -57.635 -12.075 ;
        RECT -57.965 -13.765 -57.635 -13.435 ;
        RECT -57.965 -15.125 -57.635 -14.795 ;
        RECT -57.965 -16.485 -57.635 -16.155 ;
        RECT -57.965 -17.845 -57.635 -17.515 ;
        RECT -57.965 -19.205 -57.635 -18.875 ;
        RECT -57.965 -20.565 -57.635 -20.235 ;
        RECT -57.965 -21.925 -57.635 -21.595 ;
        RECT -57.965 -23.285 -57.635 -22.955 ;
        RECT -57.965 -24.645 -57.635 -24.315 ;
        RECT -57.965 -26.005 -57.635 -25.675 ;
        RECT -57.965 -27.365 -57.635 -27.035 ;
        RECT -57.965 -28.725 -57.635 -28.395 ;
        RECT -57.965 -30.085 -57.635 -29.755 ;
        RECT -57.965 -31.445 -57.635 -31.115 ;
        RECT -57.965 -32.805 -57.635 -32.475 ;
        RECT -57.965 -34.165 -57.635 -33.835 ;
        RECT -57.965 -35.525 -57.635 -35.195 ;
        RECT -57.965 -36.885 -57.635 -36.555 ;
        RECT -57.965 -38.245 -57.635 -37.915 ;
        RECT -57.965 -39.605 -57.635 -39.275 ;
        RECT -57.965 -40.965 -57.635 -40.635 ;
        RECT -57.965 -42.325 -57.635 -41.995 ;
        RECT -57.965 -43.685 -57.635 -43.355 ;
        RECT -57.965 -45.045 -57.635 -44.715 ;
        RECT -57.965 -46.405 -57.635 -46.075 ;
        RECT -57.965 -47.765 -57.635 -47.435 ;
        RECT -57.965 -49.125 -57.635 -48.795 ;
        RECT -57.965 -50.485 -57.635 -50.155 ;
        RECT -57.965 -51.845 -57.635 -51.515 ;
        RECT -57.965 -53.205 -57.635 -52.875 ;
        RECT -57.965 -54.565 -57.635 -54.235 ;
        RECT -57.965 -55.925 -57.635 -55.595 ;
        RECT -57.965 -57.285 -57.635 -56.955 ;
        RECT -57.965 -58.645 -57.635 -58.315 ;
        RECT -57.965 -60.005 -57.635 -59.675 ;
        RECT -57.965 -61.365 -57.635 -61.035 ;
        RECT -57.965 -62.725 -57.635 -62.395 ;
        RECT -57.965 -64.085 -57.635 -63.755 ;
        RECT -57.965 -65.445 -57.635 -65.115 ;
        RECT -57.965 -66.805 -57.635 -66.475 ;
        RECT -57.965 -68.165 -57.635 -67.835 ;
        RECT -57.965 -69.525 -57.635 -69.195 ;
        RECT -57.965 -70.885 -57.635 -70.555 ;
        RECT -57.965 -72.245 -57.635 -71.915 ;
        RECT -57.965 -73.605 -57.635 -73.275 ;
        RECT -57.965 -74.965 -57.635 -74.635 ;
        RECT -57.965 -76.325 -57.635 -75.995 ;
        RECT -57.965 -77.685 -57.635 -77.355 ;
        RECT -57.965 -79.045 -57.635 -78.715 ;
        RECT -57.965 -80.405 -57.635 -80.075 ;
        RECT -57.965 -81.765 -57.635 -81.435 ;
        RECT -57.965 -83.125 -57.635 -82.795 ;
        RECT -57.965 -84.485 -57.635 -84.155 ;
        RECT -57.965 -85.845 -57.635 -85.515 ;
        RECT -57.965 -87.205 -57.635 -86.875 ;
        RECT -57.965 -88.565 -57.635 -88.235 ;
        RECT -57.965 -89.925 -57.635 -89.595 ;
        RECT -57.965 -91.285 -57.635 -90.955 ;
        RECT -57.965 -92.645 -57.635 -92.315 ;
        RECT -57.965 -94.005 -57.635 -93.675 ;
        RECT -57.965 -95.365 -57.635 -95.035 ;
        RECT -57.965 -96.725 -57.635 -96.395 ;
        RECT -57.965 -98.085 -57.635 -97.755 ;
        RECT -57.965 -99.445 -57.635 -99.115 ;
        RECT -57.965 -100.805 -57.635 -100.475 ;
        RECT -57.965 -102.165 -57.635 -101.835 ;
        RECT -57.965 -103.525 -57.635 -103.195 ;
        RECT -57.965 -104.885 -57.635 -104.555 ;
        RECT -57.965 -106.245 -57.635 -105.915 ;
        RECT -57.965 -107.605 -57.635 -107.275 ;
        RECT -57.965 -108.965 -57.635 -108.635 ;
        RECT -57.965 -110.325 -57.635 -109.995 ;
        RECT -57.965 -111.685 -57.635 -111.355 ;
        RECT -57.965 -113.045 -57.635 -112.715 ;
        RECT -57.965 -114.405 -57.635 -114.075 ;
        RECT -57.965 -115.765 -57.635 -115.435 ;
        RECT -57.965 -117.125 -57.635 -116.795 ;
        RECT -57.965 -118.485 -57.635 -118.155 ;
        RECT -57.965 -119.845 -57.635 -119.515 ;
        RECT -57.965 -121.205 -57.635 -120.875 ;
        RECT -57.965 -122.565 -57.635 -122.235 ;
        RECT -57.965 -123.925 -57.635 -123.595 ;
        RECT -57.965 -125.285 -57.635 -124.955 ;
        RECT -57.965 -126.645 -57.635 -126.315 ;
        RECT -57.965 -128.005 -57.635 -127.675 ;
        RECT -57.965 -129.365 -57.635 -129.035 ;
        RECT -57.965 -130.725 -57.635 -130.395 ;
        RECT -57.965 -132.085 -57.635 -131.755 ;
        RECT -57.965 -134.805 -57.635 -134.475 ;
        RECT -57.965 -136.165 -57.635 -135.835 ;
        RECT -57.965 -137.525 -57.635 -137.195 ;
        RECT -57.965 -138.885 -57.635 -138.555 ;
        RECT -57.965 -140.245 -57.635 -139.915 ;
        RECT -57.965 -141.605 -57.635 -141.275 ;
        RECT -57.965 -142.965 -57.635 -142.635 ;
        RECT -57.965 -144.325 -57.635 -143.995 ;
        RECT -57.965 -145.685 -57.635 -145.355 ;
        RECT -57.965 -147.045 -57.635 -146.715 ;
        RECT -57.965 -148.405 -57.635 -148.075 ;
        RECT -57.965 -149.765 -57.635 -149.435 ;
        RECT -57.965 -151.125 -57.635 -150.795 ;
        RECT -57.965 -152.485 -57.635 -152.155 ;
        RECT -57.965 -153.845 -57.635 -153.515 ;
        RECT -57.965 -155.205 -57.635 -154.875 ;
        RECT -57.965 -156.565 -57.635 -156.235 ;
        RECT -57.965 -157.925 -57.635 -157.595 ;
        RECT -57.965 -159.285 -57.635 -158.955 ;
        RECT -57.965 -160.645 -57.635 -160.315 ;
        RECT -57.965 -162.005 -57.635 -161.675 ;
        RECT -57.965 -163.365 -57.635 -163.035 ;
        RECT -57.965 -164.725 -57.635 -164.395 ;
        RECT -57.965 -166.085 -57.635 -165.755 ;
        RECT -57.965 -167.445 -57.635 -167.115 ;
        RECT -57.965 -168.805 -57.635 -168.475 ;
        RECT -57.965 -170.165 -57.635 -169.835 ;
        RECT -57.965 -171.525 -57.635 -171.195 ;
        RECT -57.965 -172.885 -57.635 -172.555 ;
        RECT -57.965 -174.245 -57.635 -173.915 ;
        RECT -57.965 -175.605 -57.635 -175.275 ;
        RECT -57.965 -176.965 -57.635 -176.635 ;
        RECT -57.965 -178.325 -57.635 -177.995 ;
        RECT -57.965 -179.685 -57.635 -179.355 ;
        RECT -57.965 -181.045 -57.635 -180.715 ;
        RECT -57.965 -182.405 -57.635 -182.075 ;
        RECT -57.965 -183.765 -57.635 -183.435 ;
        RECT -57.965 -185.125 -57.635 -184.795 ;
        RECT -57.965 -186.485 -57.635 -186.155 ;
        RECT -57.965 -187.845 -57.635 -187.515 ;
        RECT -57.965 -189.205 -57.635 -188.875 ;
        RECT -57.965 -190.565 -57.635 -190.235 ;
        RECT -57.965 -191.925 -57.635 -191.595 ;
        RECT -57.965 -193.285 -57.635 -192.955 ;
        RECT -57.965 -194.645 -57.635 -194.315 ;
        RECT -57.965 -196.005 -57.635 -195.675 ;
        RECT -57.965 -197.365 -57.635 -197.035 ;
        RECT -57.965 -198.725 -57.635 -198.395 ;
        RECT -57.965 -200.085 -57.635 -199.755 ;
        RECT -57.965 -201.445 -57.635 -201.115 ;
        RECT -57.965 -202.805 -57.635 -202.475 ;
        RECT -57.965 -204.165 -57.635 -203.835 ;
        RECT -57.965 -205.525 -57.635 -205.195 ;
        RECT -57.965 -208.245 -57.635 -207.915 ;
        RECT -57.965 -210.965 -57.635 -210.635 ;
        RECT -57.965 -212.325 -57.635 -211.995 ;
        RECT -57.965 -213.625 -57.635 -213.295 ;
        RECT -57.965 -215.045 -57.635 -214.715 ;
        RECT -57.965 -216.405 -57.635 -216.075 ;
        RECT -57.965 -217.765 -57.635 -217.435 ;
        RECT -57.965 -219.125 -57.635 -218.795 ;
        RECT -57.965 -221.37 -57.635 -220.24 ;
        RECT -57.96 -221.485 -57.64 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -56.605 129.8 -56.275 130.93 ;
        RECT -56.605 127.675 -56.275 128.005 ;
        RECT -56.605 126.315 -56.275 126.645 ;
        RECT -56.605 124.955 -56.275 125.285 ;
        RECT -56.605 123.595 -56.275 123.925 ;
        RECT -56.605 122.235 -56.275 122.565 ;
        RECT -56.605 120.875 -56.275 121.205 ;
        RECT -56.605 119.515 -56.275 119.845 ;
        RECT -56.605 118.155 -56.275 118.485 ;
        RECT -56.605 116.795 -56.275 117.125 ;
        RECT -56.605 115.435 -56.275 115.765 ;
        RECT -56.605 114.075 -56.275 114.405 ;
        RECT -56.605 112.715 -56.275 113.045 ;
        RECT -56.605 111.355 -56.275 111.685 ;
        RECT -56.605 109.995 -56.275 110.325 ;
        RECT -56.605 108.635 -56.275 108.965 ;
        RECT -56.605 107.275 -56.275 107.605 ;
        RECT -56.605 105.915 -56.275 106.245 ;
        RECT -56.605 104.555 -56.275 104.885 ;
        RECT -56.605 103.195 -56.275 103.525 ;
        RECT -56.605 101.835 -56.275 102.165 ;
        RECT -56.605 100.475 -56.275 100.805 ;
        RECT -56.605 99.115 -56.275 99.445 ;
        RECT -56.605 97.755 -56.275 98.085 ;
        RECT -56.605 96.395 -56.275 96.725 ;
        RECT -56.605 95.035 -56.275 95.365 ;
        RECT -56.605 93.675 -56.275 94.005 ;
        RECT -56.605 92.315 -56.275 92.645 ;
        RECT -56.605 90.955 -56.275 91.285 ;
        RECT -56.605 89.595 -56.275 89.925 ;
        RECT -56.605 88.235 -56.275 88.565 ;
        RECT -56.605 86.875 -56.275 87.205 ;
        RECT -56.605 85.515 -56.275 85.845 ;
        RECT -56.605 84.155 -56.275 84.485 ;
        RECT -56.605 82.795 -56.275 83.125 ;
        RECT -56.605 81.435 -56.275 81.765 ;
        RECT -56.605 80.075 -56.275 80.405 ;
        RECT -56.605 78.715 -56.275 79.045 ;
        RECT -56.605 77.355 -56.275 77.685 ;
        RECT -56.605 75.995 -56.275 76.325 ;
        RECT -56.605 74.635 -56.275 74.965 ;
        RECT -56.605 73.275 -56.275 73.605 ;
        RECT -56.605 72.445 -56.275 72.775 ;
        RECT -56.605 70.395 -56.275 70.725 ;
        RECT -56.605 68.035 -56.275 68.365 ;
        RECT -56.605 66.885 -56.275 67.215 ;
        RECT -56.605 64.875 -56.275 65.205 ;
        RECT -56.605 63.725 -56.275 64.055 ;
        RECT -56.605 61.715 -56.275 62.045 ;
        RECT -56.605 60.395 -56.275 60.725 ;
        RECT -56.605 58.555 -56.275 58.885 ;
        RECT -56.605 57.405 -56.275 57.735 ;
        RECT -56.605 55.395 -56.275 55.725 ;
        RECT -56.605 54.245 -56.275 54.575 ;
        RECT -56.605 51.885 -56.275 52.215 ;
        RECT -56.605 49.83 -56.275 50.16 ;
        RECT -56.605 48.795 -56.275 49.125 ;
        RECT -56.605 47.435 -56.275 47.765 ;
        RECT -56.605 46.075 -56.275 46.405 ;
        RECT -56.605 44.715 -56.275 45.045 ;
        RECT -56.605 43.355 -56.275 43.685 ;
        RECT -56.605 41.995 -56.275 42.325 ;
        RECT -56.605 40.635 -56.275 40.965 ;
        RECT -56.605 39.275 -56.275 39.605 ;
        RECT -56.605 37.915 -56.275 38.245 ;
        RECT -56.605 36.555 -56.275 36.885 ;
        RECT -56.605 35.195 -56.275 35.525 ;
        RECT -56.605 33.835 -56.275 34.165 ;
        RECT -56.605 32.475 -56.275 32.805 ;
        RECT -56.605 31.115 -56.275 31.445 ;
        RECT -56.605 29.755 -56.275 30.085 ;
        RECT -56.605 28.395 -56.275 28.725 ;
        RECT -56.605 27.035 -56.275 27.365 ;
        RECT -56.605 25.675 -56.275 26.005 ;
        RECT -56.605 24.315 -56.275 24.645 ;
        RECT -56.605 22.955 -56.275 23.285 ;
        RECT -56.605 21.595 -56.275 21.925 ;
        RECT -56.605 20.235 -56.275 20.565 ;
        RECT -56.605 18.875 -56.275 19.205 ;
        RECT -56.605 17.515 -56.275 17.845 ;
        RECT -56.605 16.155 -56.275 16.485 ;
        RECT -56.605 14.795 -56.275 15.125 ;
        RECT -56.605 13.435 -56.275 13.765 ;
        RECT -56.605 12.075 -56.275 12.405 ;
        RECT -56.605 10.715 -56.275 11.045 ;
        RECT -56.605 9.355 -56.275 9.685 ;
        RECT -56.605 7.995 -56.275 8.325 ;
        RECT -56.605 6.635 -56.275 6.965 ;
        RECT -56.605 5.275 -56.275 5.605 ;
        RECT -56.605 3.915 -56.275 4.245 ;
        RECT -56.605 2.555 -56.275 2.885 ;
        RECT -56.605 1.195 -56.275 1.525 ;
        RECT -56.605 -0.165 -56.275 0.165 ;
        RECT -56.605 -1.525 -56.275 -1.195 ;
        RECT -56.605 -2.885 -56.275 -2.555 ;
        RECT -56.605 -4.245 -56.275 -3.915 ;
        RECT -56.605 -5.605 -56.275 -5.275 ;
        RECT -56.605 -6.965 -56.275 -6.635 ;
        RECT -56.605 -8.325 -56.275 -7.995 ;
        RECT -56.605 -9.685 -56.275 -9.355 ;
        RECT -56.605 -11.045 -56.275 -10.715 ;
        RECT -56.605 -12.405 -56.275 -12.075 ;
        RECT -56.605 -13.765 -56.275 -13.435 ;
        RECT -56.605 -15.125 -56.275 -14.795 ;
        RECT -56.605 -16.485 -56.275 -16.155 ;
        RECT -56.605 -17.845 -56.275 -17.515 ;
        RECT -56.605 -19.205 -56.275 -18.875 ;
        RECT -56.605 -20.565 -56.275 -20.235 ;
        RECT -56.605 -21.925 -56.275 -21.595 ;
        RECT -56.605 -23.285 -56.275 -22.955 ;
        RECT -56.605 -24.645 -56.275 -24.315 ;
        RECT -56.605 -26.005 -56.275 -25.675 ;
        RECT -56.605 -27.365 -56.275 -27.035 ;
        RECT -56.605 -28.725 -56.275 -28.395 ;
        RECT -56.605 -30.085 -56.275 -29.755 ;
        RECT -56.605 -31.445 -56.275 -31.115 ;
        RECT -56.605 -32.805 -56.275 -32.475 ;
        RECT -56.605 -34.165 -56.275 -33.835 ;
        RECT -56.605 -35.525 -56.275 -35.195 ;
        RECT -56.605 -36.885 -56.275 -36.555 ;
        RECT -56.605 -38.245 -56.275 -37.915 ;
        RECT -56.605 -39.605 -56.275 -39.275 ;
        RECT -56.605 -40.965 -56.275 -40.635 ;
        RECT -56.605 -42.325 -56.275 -41.995 ;
        RECT -56.605 -43.685 -56.275 -43.355 ;
        RECT -56.605 -45.045 -56.275 -44.715 ;
        RECT -56.605 -46.405 -56.275 -46.075 ;
        RECT -56.605 -47.765 -56.275 -47.435 ;
        RECT -56.605 -49.125 -56.275 -48.795 ;
        RECT -56.605 -50.485 -56.275 -50.155 ;
        RECT -56.605 -51.845 -56.275 -51.515 ;
        RECT -56.605 -53.205 -56.275 -52.875 ;
        RECT -56.605 -54.565 -56.275 -54.235 ;
        RECT -56.605 -55.925 -56.275 -55.595 ;
        RECT -56.605 -57.285 -56.275 -56.955 ;
        RECT -56.605 -58.645 -56.275 -58.315 ;
        RECT -56.605 -60.005 -56.275 -59.675 ;
        RECT -56.605 -61.365 -56.275 -61.035 ;
        RECT -56.605 -62.725 -56.275 -62.395 ;
        RECT -56.605 -64.085 -56.275 -63.755 ;
        RECT -56.605 -65.445 -56.275 -65.115 ;
        RECT -56.605 -66.805 -56.275 -66.475 ;
        RECT -56.605 -68.165 -56.275 -67.835 ;
        RECT -56.605 -69.525 -56.275 -69.195 ;
        RECT -56.605 -70.885 -56.275 -70.555 ;
        RECT -56.605 -72.245 -56.275 -71.915 ;
        RECT -56.605 -73.605 -56.275 -73.275 ;
        RECT -56.605 -74.965 -56.275 -74.635 ;
        RECT -56.605 -76.325 -56.275 -75.995 ;
        RECT -56.605 -77.685 -56.275 -77.355 ;
        RECT -56.605 -79.045 -56.275 -78.715 ;
        RECT -56.605 -80.405 -56.275 -80.075 ;
        RECT -56.605 -81.765 -56.275 -81.435 ;
        RECT -56.605 -83.125 -56.275 -82.795 ;
        RECT -56.605 -84.485 -56.275 -84.155 ;
        RECT -56.605 -85.845 -56.275 -85.515 ;
        RECT -56.605 -87.205 -56.275 -86.875 ;
        RECT -56.605 -88.565 -56.275 -88.235 ;
        RECT -56.605 -89.925 -56.275 -89.595 ;
        RECT -56.605 -91.285 -56.275 -90.955 ;
        RECT -56.605 -92.645 -56.275 -92.315 ;
        RECT -56.605 -94.005 -56.275 -93.675 ;
        RECT -56.605 -95.365 -56.275 -95.035 ;
        RECT -56.605 -96.725 -56.275 -96.395 ;
        RECT -56.605 -98.085 -56.275 -97.755 ;
        RECT -56.605 -99.445 -56.275 -99.115 ;
        RECT -56.605 -100.805 -56.275 -100.475 ;
        RECT -56.605 -102.165 -56.275 -101.835 ;
        RECT -56.605 -103.525 -56.275 -103.195 ;
        RECT -56.605 -104.885 -56.275 -104.555 ;
        RECT -56.605 -106.245 -56.275 -105.915 ;
        RECT -56.605 -107.605 -56.275 -107.275 ;
        RECT -56.605 -108.965 -56.275 -108.635 ;
        RECT -56.605 -110.325 -56.275 -109.995 ;
        RECT -56.605 -113.045 -56.275 -112.715 ;
        RECT -56.605 -114.405 -56.275 -114.075 ;
        RECT -56.605 -115.765 -56.275 -115.435 ;
        RECT -56.605 -117.125 -56.275 -116.795 ;
        RECT -56.605 -118.485 -56.275 -118.155 ;
        RECT -56.605 -121.205 -56.275 -120.875 ;
        RECT -56.605 -122.565 -56.275 -122.235 ;
        RECT -56.605 -123.925 -56.275 -123.595 ;
        RECT -56.605 -126.645 -56.275 -126.315 ;
        RECT -56.605 -129.365 -56.275 -129.035 ;
        RECT -56.605 -130.725 -56.275 -130.395 ;
        RECT -56.6 -131.4 -56.28 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -56.605 -141.605 -56.275 -141.275 ;
        RECT -56.605 -142.965 -56.275 -142.635 ;
        RECT -56.605 -144.325 -56.275 -143.995 ;
        RECT -56.605 -145.685 -56.275 -145.355 ;
        RECT -56.605 -147.045 -56.275 -146.715 ;
        RECT -56.605 -148.405 -56.275 -148.075 ;
        RECT -56.605 -149.765 -56.275 -149.435 ;
        RECT -56.605 -151.125 -56.275 -150.795 ;
        RECT -56.605 -152.485 -56.275 -152.155 ;
        RECT -56.605 -153.845 -56.275 -153.515 ;
        RECT -56.605 -155.205 -56.275 -154.875 ;
        RECT -56.605 -156.565 -56.275 -156.235 ;
        RECT -56.605 -157.925 -56.275 -157.595 ;
        RECT -56.605 -159.285 -56.275 -158.955 ;
        RECT -56.605 -160.645 -56.275 -160.315 ;
        RECT -56.605 -162.005 -56.275 -161.675 ;
        RECT -56.605 -163.365 -56.275 -163.035 ;
        RECT -56.605 -164.725 -56.275 -164.395 ;
        RECT -56.605 -166.085 -56.275 -165.755 ;
        RECT -56.605 -167.445 -56.275 -167.115 ;
        RECT -56.605 -168.805 -56.275 -168.475 ;
        RECT -56.605 -170.165 -56.275 -169.835 ;
        RECT -56.605 -171.525 -56.275 -171.195 ;
        RECT -56.605 -172.885 -56.275 -172.555 ;
        RECT -56.605 -174.245 -56.275 -173.915 ;
        RECT -56.605 -175.605 -56.275 -175.275 ;
        RECT -56.605 -176.965 -56.275 -176.635 ;
        RECT -56.605 -178.325 -56.275 -177.995 ;
        RECT -56.605 -179.685 -56.275 -179.355 ;
        RECT -56.605 -181.045 -56.275 -180.715 ;
        RECT -56.605 -182.405 -56.275 -182.075 ;
        RECT -56.605 -183.765 -56.275 -183.435 ;
        RECT -56.605 -185.125 -56.275 -184.795 ;
        RECT -56.605 -186.485 -56.275 -186.155 ;
        RECT -56.605 -187.845 -56.275 -187.515 ;
        RECT -56.605 -189.205 -56.275 -188.875 ;
        RECT -56.605 -190.565 -56.275 -190.235 ;
        RECT -56.605 -191.925 -56.275 -191.595 ;
        RECT -56.605 -193.285 -56.275 -192.955 ;
        RECT -56.605 -194.645 -56.275 -194.315 ;
        RECT -56.605 -196.005 -56.275 -195.675 ;
        RECT -56.605 -197.365 -56.275 -197.035 ;
        RECT -56.605 -198.725 -56.275 -198.395 ;
        RECT -56.605 -200.085 -56.275 -199.755 ;
        RECT -56.605 -201.445 -56.275 -201.115 ;
        RECT -56.605 -202.805 -56.275 -202.475 ;
        RECT -56.605 -204.165 -56.275 -203.835 ;
        RECT -56.605 -205.525 -56.275 -205.195 ;
        RECT -56.605 -208.245 -56.275 -207.915 ;
        RECT -56.605 -210.965 -56.275 -210.635 ;
        RECT -56.605 -212.325 -56.275 -211.995 ;
        RECT -56.605 -213.625 -56.275 -213.295 ;
        RECT -56.605 -215.045 -56.275 -214.715 ;
        RECT -56.605 -216.405 -56.275 -216.075 ;
        RECT -56.605 -217.765 -56.275 -217.435 ;
        RECT -56.605 -219.125 -56.275 -218.795 ;
        RECT -56.605 -221.37 -56.275 -220.24 ;
        RECT -56.6 -221.485 -56.28 -141.275 ;
    END
    PORT
      LAYER met3 ;
        RECT -55.245 129.8 -54.915 130.93 ;
        RECT -55.245 127.675 -54.915 128.005 ;
        RECT -55.245 126.315 -54.915 126.645 ;
        RECT -55.245 124.955 -54.915 125.285 ;
        RECT -55.245 123.595 -54.915 123.925 ;
        RECT -55.245 122.235 -54.915 122.565 ;
        RECT -55.245 120.875 -54.915 121.205 ;
        RECT -55.245 119.515 -54.915 119.845 ;
        RECT -55.245 118.155 -54.915 118.485 ;
        RECT -55.245 116.795 -54.915 117.125 ;
        RECT -55.245 115.435 -54.915 115.765 ;
        RECT -55.245 114.075 -54.915 114.405 ;
        RECT -55.245 112.715 -54.915 113.045 ;
        RECT -55.245 111.355 -54.915 111.685 ;
        RECT -55.245 109.995 -54.915 110.325 ;
        RECT -55.245 108.635 -54.915 108.965 ;
        RECT -55.245 107.275 -54.915 107.605 ;
        RECT -55.245 105.915 -54.915 106.245 ;
        RECT -55.245 104.555 -54.915 104.885 ;
        RECT -55.245 103.195 -54.915 103.525 ;
        RECT -55.245 101.835 -54.915 102.165 ;
        RECT -55.245 100.475 -54.915 100.805 ;
        RECT -55.245 99.115 -54.915 99.445 ;
        RECT -55.245 97.755 -54.915 98.085 ;
        RECT -55.245 96.395 -54.915 96.725 ;
        RECT -55.245 95.035 -54.915 95.365 ;
        RECT -55.245 93.675 -54.915 94.005 ;
        RECT -55.245 92.315 -54.915 92.645 ;
        RECT -55.245 90.955 -54.915 91.285 ;
        RECT -55.245 89.595 -54.915 89.925 ;
        RECT -55.245 88.235 -54.915 88.565 ;
        RECT -55.245 86.875 -54.915 87.205 ;
        RECT -55.245 85.515 -54.915 85.845 ;
        RECT -55.245 84.155 -54.915 84.485 ;
        RECT -55.245 82.795 -54.915 83.125 ;
        RECT -55.245 81.435 -54.915 81.765 ;
        RECT -55.245 80.075 -54.915 80.405 ;
        RECT -55.245 78.715 -54.915 79.045 ;
        RECT -55.245 77.355 -54.915 77.685 ;
        RECT -55.245 75.995 -54.915 76.325 ;
        RECT -55.245 74.635 -54.915 74.965 ;
        RECT -55.245 73.275 -54.915 73.605 ;
        RECT -55.245 72.445 -54.915 72.775 ;
        RECT -55.245 70.395 -54.915 70.725 ;
        RECT -55.245 68.035 -54.915 68.365 ;
        RECT -55.245 66.885 -54.915 67.215 ;
        RECT -55.245 64.875 -54.915 65.205 ;
        RECT -55.245 63.725 -54.915 64.055 ;
        RECT -55.245 61.715 -54.915 62.045 ;
        RECT -55.245 60.395 -54.915 60.725 ;
        RECT -55.245 58.555 -54.915 58.885 ;
        RECT -55.245 57.405 -54.915 57.735 ;
        RECT -55.245 55.395 -54.915 55.725 ;
        RECT -55.245 54.245 -54.915 54.575 ;
        RECT -55.245 51.885 -54.915 52.215 ;
        RECT -55.245 49.83 -54.915 50.16 ;
        RECT -55.245 48.795 -54.915 49.125 ;
        RECT -55.245 47.435 -54.915 47.765 ;
        RECT -55.245 46.075 -54.915 46.405 ;
        RECT -55.245 44.715 -54.915 45.045 ;
        RECT -55.245 43.355 -54.915 43.685 ;
        RECT -55.245 41.995 -54.915 42.325 ;
        RECT -55.245 40.635 -54.915 40.965 ;
        RECT -55.245 39.275 -54.915 39.605 ;
        RECT -55.245 37.915 -54.915 38.245 ;
        RECT -55.245 36.555 -54.915 36.885 ;
        RECT -55.245 35.195 -54.915 35.525 ;
        RECT -55.245 33.835 -54.915 34.165 ;
        RECT -55.245 32.475 -54.915 32.805 ;
        RECT -55.245 31.115 -54.915 31.445 ;
        RECT -55.245 29.755 -54.915 30.085 ;
        RECT -55.245 28.395 -54.915 28.725 ;
        RECT -55.245 27.035 -54.915 27.365 ;
        RECT -55.245 25.675 -54.915 26.005 ;
        RECT -55.245 24.315 -54.915 24.645 ;
        RECT -55.245 22.955 -54.915 23.285 ;
        RECT -55.245 21.595 -54.915 21.925 ;
        RECT -55.245 20.235 -54.915 20.565 ;
        RECT -55.245 18.875 -54.915 19.205 ;
        RECT -55.245 17.515 -54.915 17.845 ;
        RECT -55.245 16.155 -54.915 16.485 ;
        RECT -55.245 14.795 -54.915 15.125 ;
        RECT -55.245 13.435 -54.915 13.765 ;
        RECT -55.245 12.075 -54.915 12.405 ;
        RECT -55.245 10.715 -54.915 11.045 ;
        RECT -55.245 9.355 -54.915 9.685 ;
        RECT -55.245 7.995 -54.915 8.325 ;
        RECT -55.245 6.635 -54.915 6.965 ;
        RECT -55.245 5.275 -54.915 5.605 ;
        RECT -55.245 3.915 -54.915 4.245 ;
        RECT -55.245 2.555 -54.915 2.885 ;
        RECT -55.245 1.195 -54.915 1.525 ;
        RECT -55.245 -0.165 -54.915 0.165 ;
        RECT -55.245 -1.525 -54.915 -1.195 ;
        RECT -55.245 -2.885 -54.915 -2.555 ;
        RECT -55.245 -4.245 -54.915 -3.915 ;
        RECT -55.245 -5.605 -54.915 -5.275 ;
        RECT -55.245 -6.965 -54.915 -6.635 ;
        RECT -55.245 -8.325 -54.915 -7.995 ;
        RECT -55.245 -9.685 -54.915 -9.355 ;
        RECT -55.245 -11.045 -54.915 -10.715 ;
        RECT -55.245 -12.405 -54.915 -12.075 ;
        RECT -55.245 -13.765 -54.915 -13.435 ;
        RECT -55.245 -15.125 -54.915 -14.795 ;
        RECT -55.245 -16.485 -54.915 -16.155 ;
        RECT -55.245 -17.845 -54.915 -17.515 ;
        RECT -55.245 -19.205 -54.915 -18.875 ;
        RECT -55.245 -20.565 -54.915 -20.235 ;
        RECT -55.245 -21.925 -54.915 -21.595 ;
        RECT -55.245 -23.285 -54.915 -22.955 ;
        RECT -55.245 -24.645 -54.915 -24.315 ;
        RECT -55.245 -26.005 -54.915 -25.675 ;
        RECT -55.245 -27.365 -54.915 -27.035 ;
        RECT -55.245 -28.725 -54.915 -28.395 ;
        RECT -55.245 -30.085 -54.915 -29.755 ;
        RECT -55.245 -31.445 -54.915 -31.115 ;
        RECT -55.245 -32.805 -54.915 -32.475 ;
        RECT -55.245 -34.165 -54.915 -33.835 ;
        RECT -55.245 -35.525 -54.915 -35.195 ;
        RECT -55.245 -36.885 -54.915 -36.555 ;
        RECT -55.245 -38.245 -54.915 -37.915 ;
        RECT -55.245 -39.605 -54.915 -39.275 ;
        RECT -55.245 -40.965 -54.915 -40.635 ;
        RECT -55.245 -42.325 -54.915 -41.995 ;
        RECT -55.245 -43.685 -54.915 -43.355 ;
        RECT -55.245 -45.045 -54.915 -44.715 ;
        RECT -55.245 -46.405 -54.915 -46.075 ;
        RECT -55.245 -47.765 -54.915 -47.435 ;
        RECT -55.245 -49.125 -54.915 -48.795 ;
        RECT -55.245 -50.485 -54.915 -50.155 ;
        RECT -55.245 -51.845 -54.915 -51.515 ;
        RECT -55.245 -53.205 -54.915 -52.875 ;
        RECT -55.245 -54.565 -54.915 -54.235 ;
        RECT -55.245 -55.925 -54.915 -55.595 ;
        RECT -55.245 -57.285 -54.915 -56.955 ;
        RECT -55.245 -58.645 -54.915 -58.315 ;
        RECT -55.245 -60.005 -54.915 -59.675 ;
        RECT -55.245 -61.365 -54.915 -61.035 ;
        RECT -55.245 -62.725 -54.915 -62.395 ;
        RECT -55.245 -64.085 -54.915 -63.755 ;
        RECT -55.245 -65.445 -54.915 -65.115 ;
        RECT -55.245 -66.805 -54.915 -66.475 ;
        RECT -55.245 -68.165 -54.915 -67.835 ;
        RECT -55.245 -69.525 -54.915 -69.195 ;
        RECT -55.245 -70.885 -54.915 -70.555 ;
        RECT -55.245 -72.245 -54.915 -71.915 ;
        RECT -55.245 -73.605 -54.915 -73.275 ;
        RECT -55.245 -74.965 -54.915 -74.635 ;
        RECT -55.245 -76.325 -54.915 -75.995 ;
        RECT -55.245 -77.685 -54.915 -77.355 ;
        RECT -55.245 -79.045 -54.915 -78.715 ;
        RECT -55.245 -80.405 -54.915 -80.075 ;
        RECT -55.245 -81.765 -54.915 -81.435 ;
        RECT -55.245 -83.125 -54.915 -82.795 ;
        RECT -55.245 -84.485 -54.915 -84.155 ;
        RECT -55.245 -85.845 -54.915 -85.515 ;
        RECT -55.245 -87.205 -54.915 -86.875 ;
        RECT -55.245 -88.565 -54.915 -88.235 ;
        RECT -55.245 -89.925 -54.915 -89.595 ;
        RECT -55.245 -91.285 -54.915 -90.955 ;
        RECT -55.245 -92.645 -54.915 -92.315 ;
        RECT -55.245 -94.005 -54.915 -93.675 ;
        RECT -55.245 -95.365 -54.915 -95.035 ;
        RECT -55.245 -96.725 -54.915 -96.395 ;
        RECT -55.245 -98.085 -54.915 -97.755 ;
        RECT -55.245 -99.445 -54.915 -99.115 ;
        RECT -55.245 -100.805 -54.915 -100.475 ;
        RECT -55.245 -102.165 -54.915 -101.835 ;
        RECT -55.245 -103.525 -54.915 -103.195 ;
        RECT -55.245 -104.885 -54.915 -104.555 ;
        RECT -55.245 -106.245 -54.915 -105.915 ;
        RECT -55.245 -107.605 -54.915 -107.275 ;
        RECT -55.245 -108.965 -54.915 -108.635 ;
        RECT -55.245 -110.325 -54.915 -109.995 ;
        RECT -55.245 -113.045 -54.915 -112.715 ;
        RECT -55.245 -114.405 -54.915 -114.075 ;
        RECT -55.245 -115.765 -54.915 -115.435 ;
        RECT -55.245 -117.125 -54.915 -116.795 ;
        RECT -55.245 -118.485 -54.915 -118.155 ;
        RECT -55.245 -119.79 -54.915 -119.46 ;
        RECT -55.245 -121.205 -54.915 -120.875 ;
        RECT -55.245 -122.565 -54.915 -122.235 ;
        RECT -55.245 -123.925 -54.915 -123.595 ;
        RECT -55.245 -126.645 -54.915 -126.315 ;
        RECT -55.245 -128.43 -54.915 -128.1 ;
        RECT -55.245 -129.365 -54.915 -129.035 ;
        RECT -55.245 -130.725 -54.915 -130.395 ;
        RECT -55.245 -134.805 -54.915 -134.475 ;
        RECT -55.245 -136.165 -54.915 -135.835 ;
        RECT -55.245 -137.525 -54.915 -137.195 ;
        RECT -55.245 -138.885 -54.915 -138.555 ;
        RECT -55.245 -140.245 -54.915 -139.915 ;
        RECT -55.245 -141.605 -54.915 -141.275 ;
        RECT -55.245 -142.965 -54.915 -142.635 ;
        RECT -55.245 -144.325 -54.915 -143.995 ;
        RECT -55.245 -145.685 -54.915 -145.355 ;
        RECT -55.245 -147.045 -54.915 -146.715 ;
        RECT -55.245 -148.405 -54.915 -148.075 ;
        RECT -55.245 -149.765 -54.915 -149.435 ;
        RECT -55.245 -151.125 -54.915 -150.795 ;
        RECT -55.245 -152.485 -54.915 -152.155 ;
        RECT -55.245 -153.845 -54.915 -153.515 ;
        RECT -55.245 -155.205 -54.915 -154.875 ;
        RECT -55.245 -156.565 -54.915 -156.235 ;
        RECT -55.245 -157.925 -54.915 -157.595 ;
        RECT -55.245 -159.285 -54.915 -158.955 ;
        RECT -55.245 -160.645 -54.915 -160.315 ;
        RECT -55.245 -162.005 -54.915 -161.675 ;
        RECT -55.245 -163.365 -54.915 -163.035 ;
        RECT -55.245 -164.725 -54.915 -164.395 ;
        RECT -55.245 -166.085 -54.915 -165.755 ;
        RECT -55.245 -167.445 -54.915 -167.115 ;
        RECT -55.245 -168.805 -54.915 -168.475 ;
        RECT -55.245 -170.165 -54.915 -169.835 ;
        RECT -55.245 -171.525 -54.915 -171.195 ;
        RECT -55.245 -172.885 -54.915 -172.555 ;
        RECT -55.245 -174.245 -54.915 -173.915 ;
        RECT -55.245 -175.605 -54.915 -175.275 ;
        RECT -55.245 -176.965 -54.915 -176.635 ;
        RECT -55.245 -178.325 -54.915 -177.995 ;
        RECT -55.245 -179.685 -54.915 -179.355 ;
        RECT -55.245 -181.045 -54.915 -180.715 ;
        RECT -55.245 -182.405 -54.915 -182.075 ;
        RECT -55.245 -183.765 -54.915 -183.435 ;
        RECT -55.245 -185.125 -54.915 -184.795 ;
        RECT -55.245 -186.485 -54.915 -186.155 ;
        RECT -55.245 -187.845 -54.915 -187.515 ;
        RECT -55.245 -189.205 -54.915 -188.875 ;
        RECT -55.245 -190.565 -54.915 -190.235 ;
        RECT -55.245 -191.925 -54.915 -191.595 ;
        RECT -55.245 -193.285 -54.915 -192.955 ;
        RECT -55.245 -194.645 -54.915 -194.315 ;
        RECT -55.245 -196.005 -54.915 -195.675 ;
        RECT -55.245 -197.365 -54.915 -197.035 ;
        RECT -55.245 -198.725 -54.915 -198.395 ;
        RECT -55.245 -200.085 -54.915 -199.755 ;
        RECT -55.245 -201.445 -54.915 -201.115 ;
        RECT -55.245 -202.805 -54.915 -202.475 ;
        RECT -55.245 -204.165 -54.915 -203.835 ;
        RECT -55.245 -205.525 -54.915 -205.195 ;
        RECT -55.245 -208.245 -54.915 -207.915 ;
        RECT -55.245 -210.965 -54.915 -210.635 ;
        RECT -55.245 -212.325 -54.915 -211.995 ;
        RECT -55.245 -213.625 -54.915 -213.295 ;
        RECT -55.245 -215.045 -54.915 -214.715 ;
        RECT -55.245 -216.405 -54.915 -216.075 ;
        RECT -55.245 -217.765 -54.915 -217.435 ;
        RECT -55.245 -219.125 -54.915 -218.795 ;
        RECT -55.245 -221.37 -54.915 -220.24 ;
        RECT -55.24 -221.485 -54.92 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.885 -62.725 -53.555 -62.395 ;
        RECT -53.885 -64.085 -53.555 -63.755 ;
        RECT -53.885 -65.445 -53.555 -65.115 ;
        RECT -53.885 -66.805 -53.555 -66.475 ;
        RECT -53.885 -68.165 -53.555 -67.835 ;
        RECT -53.885 -69.525 -53.555 -69.195 ;
        RECT -53.885 -70.885 -53.555 -70.555 ;
        RECT -53.885 -72.245 -53.555 -71.915 ;
        RECT -53.885 -73.605 -53.555 -73.275 ;
        RECT -53.885 -74.965 -53.555 -74.635 ;
        RECT -53.885 -76.325 -53.555 -75.995 ;
        RECT -53.885 -77.685 -53.555 -77.355 ;
        RECT -53.885 -79.045 -53.555 -78.715 ;
        RECT -53.885 -80.405 -53.555 -80.075 ;
        RECT -53.885 -81.765 -53.555 -81.435 ;
        RECT -53.885 -83.125 -53.555 -82.795 ;
        RECT -53.885 -84.485 -53.555 -84.155 ;
        RECT -53.885 -85.845 -53.555 -85.515 ;
        RECT -53.885 -87.205 -53.555 -86.875 ;
        RECT -53.885 -88.565 -53.555 -88.235 ;
        RECT -53.885 -89.925 -53.555 -89.595 ;
        RECT -53.885 -91.285 -53.555 -90.955 ;
        RECT -53.885 -92.645 -53.555 -92.315 ;
        RECT -53.885 -94.005 -53.555 -93.675 ;
        RECT -53.885 -95.365 -53.555 -95.035 ;
        RECT -53.885 -96.725 -53.555 -96.395 ;
        RECT -53.885 -98.085 -53.555 -97.755 ;
        RECT -53.885 -99.445 -53.555 -99.115 ;
        RECT -53.885 -100.805 -53.555 -100.475 ;
        RECT -53.885 -102.165 -53.555 -101.835 ;
        RECT -53.885 -103.525 -53.555 -103.195 ;
        RECT -53.885 -104.885 -53.555 -104.555 ;
        RECT -53.885 -106.245 -53.555 -105.915 ;
        RECT -53.885 -107.605 -53.555 -107.275 ;
        RECT -53.885 -108.965 -53.555 -108.635 ;
        RECT -53.885 -110.325 -53.555 -109.995 ;
        RECT -53.885 -113.045 -53.555 -112.715 ;
        RECT -53.885 -114.405 -53.555 -114.075 ;
        RECT -53.885 -115.765 -53.555 -115.435 ;
        RECT -53.885 -117.125 -53.555 -116.795 ;
        RECT -53.885 -118.485 -53.555 -118.155 ;
        RECT -53.885 -119.79 -53.555 -119.46 ;
        RECT -53.885 -121.205 -53.555 -120.875 ;
        RECT -53.885 -122.565 -53.555 -122.235 ;
        RECT -53.885 -123.925 -53.555 -123.595 ;
        RECT -53.885 -126.645 -53.555 -126.315 ;
        RECT -53.885 -128.43 -53.555 -128.1 ;
        RECT -53.885 -129.365 -53.555 -129.035 ;
        RECT -53.885 -130.725 -53.555 -130.395 ;
        RECT -53.885 -134.805 -53.555 -134.475 ;
        RECT -53.885 -136.165 -53.555 -135.835 ;
        RECT -53.885 -137.525 -53.555 -137.195 ;
        RECT -53.885 -138.885 -53.555 -138.555 ;
        RECT -53.885 -140.245 -53.555 -139.915 ;
        RECT -53.885 -141.605 -53.555 -141.275 ;
        RECT -53.885 -142.965 -53.555 -142.635 ;
        RECT -53.885 -144.325 -53.555 -143.995 ;
        RECT -53.885 -145.685 -53.555 -145.355 ;
        RECT -53.885 -147.045 -53.555 -146.715 ;
        RECT -53.885 -148.405 -53.555 -148.075 ;
        RECT -53.885 -149.765 -53.555 -149.435 ;
        RECT -53.885 -151.125 -53.555 -150.795 ;
        RECT -53.885 -152.485 -53.555 -152.155 ;
        RECT -53.885 -153.845 -53.555 -153.515 ;
        RECT -53.885 -155.205 -53.555 -154.875 ;
        RECT -53.885 -156.565 -53.555 -156.235 ;
        RECT -53.885 -157.925 -53.555 -157.595 ;
        RECT -53.885 -159.285 -53.555 -158.955 ;
        RECT -53.885 -160.645 -53.555 -160.315 ;
        RECT -53.885 -162.005 -53.555 -161.675 ;
        RECT -53.885 -163.365 -53.555 -163.035 ;
        RECT -53.885 -164.725 -53.555 -164.395 ;
        RECT -53.885 -166.085 -53.555 -165.755 ;
        RECT -53.885 -167.445 -53.555 -167.115 ;
        RECT -53.885 -168.805 -53.555 -168.475 ;
        RECT -53.885 -170.165 -53.555 -169.835 ;
        RECT -53.885 -171.525 -53.555 -171.195 ;
        RECT -53.885 -172.885 -53.555 -172.555 ;
        RECT -53.885 -174.245 -53.555 -173.915 ;
        RECT -53.885 -175.605 -53.555 -175.275 ;
        RECT -53.885 -176.965 -53.555 -176.635 ;
        RECT -53.885 -178.325 -53.555 -177.995 ;
        RECT -53.885 -179.685 -53.555 -179.355 ;
        RECT -53.885 -181.045 -53.555 -180.715 ;
        RECT -53.885 -182.405 -53.555 -182.075 ;
        RECT -53.885 -183.765 -53.555 -183.435 ;
        RECT -53.885 -185.125 -53.555 -184.795 ;
        RECT -53.885 -186.485 -53.555 -186.155 ;
        RECT -53.885 -187.845 -53.555 -187.515 ;
        RECT -53.885 -189.205 -53.555 -188.875 ;
        RECT -53.885 -190.565 -53.555 -190.235 ;
        RECT -53.885 -191.925 -53.555 -191.595 ;
        RECT -53.885 -193.285 -53.555 -192.955 ;
        RECT -53.885 -194.645 -53.555 -194.315 ;
        RECT -53.885 -196.005 -53.555 -195.675 ;
        RECT -53.885 -197.365 -53.555 -197.035 ;
        RECT -53.885 -198.725 -53.555 -198.395 ;
        RECT -53.885 -200.085 -53.555 -199.755 ;
        RECT -53.885 -201.445 -53.555 -201.115 ;
        RECT -53.885 -202.805 -53.555 -202.475 ;
        RECT -53.885 -204.165 -53.555 -203.835 ;
        RECT -53.885 -205.525 -53.555 -205.195 ;
        RECT -53.885 -208.245 -53.555 -207.915 ;
        RECT -53.885 -212.325 -53.555 -211.995 ;
        RECT -53.885 -213.625 -53.555 -213.295 ;
        RECT -53.885 -215.045 -53.555 -214.715 ;
        RECT -53.885 -216.405 -53.555 -216.075 ;
        RECT -53.885 -217.765 -53.555 -217.435 ;
        RECT -53.885 -219.125 -53.555 -218.795 ;
        RECT -53.885 -221.37 -53.555 -220.24 ;
        RECT -53.88 -221.485 -53.56 131.045 ;
        RECT -53.885 129.8 -53.555 130.93 ;
        RECT -53.885 127.675 -53.555 128.005 ;
        RECT -53.885 126.315 -53.555 126.645 ;
        RECT -53.885 124.955 -53.555 125.285 ;
        RECT -53.885 123.595 -53.555 123.925 ;
        RECT -53.885 122.235 -53.555 122.565 ;
        RECT -53.885 120.875 -53.555 121.205 ;
        RECT -53.885 119.515 -53.555 119.845 ;
        RECT -53.885 118.155 -53.555 118.485 ;
        RECT -53.885 116.795 -53.555 117.125 ;
        RECT -53.885 115.435 -53.555 115.765 ;
        RECT -53.885 114.075 -53.555 114.405 ;
        RECT -53.885 112.715 -53.555 113.045 ;
        RECT -53.885 111.355 -53.555 111.685 ;
        RECT -53.885 109.995 -53.555 110.325 ;
        RECT -53.885 108.635 -53.555 108.965 ;
        RECT -53.885 107.275 -53.555 107.605 ;
        RECT -53.885 105.915 -53.555 106.245 ;
        RECT -53.885 104.555 -53.555 104.885 ;
        RECT -53.885 103.195 -53.555 103.525 ;
        RECT -53.885 101.835 -53.555 102.165 ;
        RECT -53.885 100.475 -53.555 100.805 ;
        RECT -53.885 99.115 -53.555 99.445 ;
        RECT -53.885 97.755 -53.555 98.085 ;
        RECT -53.885 96.395 -53.555 96.725 ;
        RECT -53.885 95.035 -53.555 95.365 ;
        RECT -53.885 93.675 -53.555 94.005 ;
        RECT -53.885 92.315 -53.555 92.645 ;
        RECT -53.885 90.955 -53.555 91.285 ;
        RECT -53.885 89.595 -53.555 89.925 ;
        RECT -53.885 88.235 -53.555 88.565 ;
        RECT -53.885 86.875 -53.555 87.205 ;
        RECT -53.885 85.515 -53.555 85.845 ;
        RECT -53.885 84.155 -53.555 84.485 ;
        RECT -53.885 82.795 -53.555 83.125 ;
        RECT -53.885 81.435 -53.555 81.765 ;
        RECT -53.885 80.075 -53.555 80.405 ;
        RECT -53.885 78.715 -53.555 79.045 ;
        RECT -53.885 77.355 -53.555 77.685 ;
        RECT -53.885 75.995 -53.555 76.325 ;
        RECT -53.885 74.635 -53.555 74.965 ;
        RECT -53.885 73.275 -53.555 73.605 ;
        RECT -53.885 72.445 -53.555 72.775 ;
        RECT -53.885 70.395 -53.555 70.725 ;
        RECT -53.885 68.035 -53.555 68.365 ;
        RECT -53.885 66.885 -53.555 67.215 ;
        RECT -53.885 64.875 -53.555 65.205 ;
        RECT -53.885 63.725 -53.555 64.055 ;
        RECT -53.885 61.715 -53.555 62.045 ;
        RECT -53.885 60.395 -53.555 60.725 ;
        RECT -53.885 58.555 -53.555 58.885 ;
        RECT -53.885 57.405 -53.555 57.735 ;
        RECT -53.885 55.395 -53.555 55.725 ;
        RECT -53.885 54.245 -53.555 54.575 ;
        RECT -53.885 51.885 -53.555 52.215 ;
        RECT -53.885 49.83 -53.555 50.16 ;
        RECT -53.885 48.795 -53.555 49.125 ;
        RECT -53.885 47.435 -53.555 47.765 ;
        RECT -53.885 46.075 -53.555 46.405 ;
        RECT -53.885 44.715 -53.555 45.045 ;
        RECT -53.885 43.355 -53.555 43.685 ;
        RECT -53.885 41.995 -53.555 42.325 ;
        RECT -53.885 40.635 -53.555 40.965 ;
        RECT -53.885 39.275 -53.555 39.605 ;
        RECT -53.885 37.915 -53.555 38.245 ;
        RECT -53.885 36.555 -53.555 36.885 ;
        RECT -53.885 35.195 -53.555 35.525 ;
        RECT -53.885 33.835 -53.555 34.165 ;
        RECT -53.885 32.475 -53.555 32.805 ;
        RECT -53.885 31.115 -53.555 31.445 ;
        RECT -53.885 29.755 -53.555 30.085 ;
        RECT -53.885 28.395 -53.555 28.725 ;
        RECT -53.885 27.035 -53.555 27.365 ;
        RECT -53.885 25.675 -53.555 26.005 ;
        RECT -53.885 24.315 -53.555 24.645 ;
        RECT -53.885 22.955 -53.555 23.285 ;
        RECT -53.885 21.595 -53.555 21.925 ;
        RECT -53.885 20.235 -53.555 20.565 ;
        RECT -53.885 18.875 -53.555 19.205 ;
        RECT -53.885 17.515 -53.555 17.845 ;
        RECT -53.885 16.155 -53.555 16.485 ;
        RECT -53.885 14.795 -53.555 15.125 ;
        RECT -53.885 13.435 -53.555 13.765 ;
        RECT -53.885 12.075 -53.555 12.405 ;
        RECT -53.885 10.715 -53.555 11.045 ;
        RECT -53.885 9.355 -53.555 9.685 ;
        RECT -53.885 7.995 -53.555 8.325 ;
        RECT -53.885 6.635 -53.555 6.965 ;
        RECT -53.885 5.275 -53.555 5.605 ;
        RECT -53.885 3.915 -53.555 4.245 ;
        RECT -53.885 2.555 -53.555 2.885 ;
        RECT -53.885 1.195 -53.555 1.525 ;
        RECT -53.885 -0.165 -53.555 0.165 ;
        RECT -53.885 -1.525 -53.555 -1.195 ;
        RECT -53.885 -2.885 -53.555 -2.555 ;
        RECT -53.885 -4.245 -53.555 -3.915 ;
        RECT -53.885 -5.605 -53.555 -5.275 ;
        RECT -53.885 -6.965 -53.555 -6.635 ;
        RECT -53.885 -8.325 -53.555 -7.995 ;
        RECT -53.885 -9.685 -53.555 -9.355 ;
        RECT -53.885 -11.045 -53.555 -10.715 ;
        RECT -53.885 -12.405 -53.555 -12.075 ;
        RECT -53.885 -13.765 -53.555 -13.435 ;
        RECT -53.885 -15.125 -53.555 -14.795 ;
        RECT -53.885 -16.485 -53.555 -16.155 ;
        RECT -53.885 -17.845 -53.555 -17.515 ;
        RECT -53.885 -19.205 -53.555 -18.875 ;
        RECT -53.885 -20.565 -53.555 -20.235 ;
        RECT -53.885 -21.925 -53.555 -21.595 ;
        RECT -53.885 -23.285 -53.555 -22.955 ;
        RECT -53.885 -24.645 -53.555 -24.315 ;
        RECT -53.885 -26.005 -53.555 -25.675 ;
        RECT -53.885 -27.365 -53.555 -27.035 ;
        RECT -53.885 -28.725 -53.555 -28.395 ;
        RECT -53.885 -30.085 -53.555 -29.755 ;
        RECT -53.885 -31.445 -53.555 -31.115 ;
        RECT -53.885 -32.805 -53.555 -32.475 ;
        RECT -53.885 -34.165 -53.555 -33.835 ;
        RECT -53.885 -35.525 -53.555 -35.195 ;
        RECT -53.885 -36.885 -53.555 -36.555 ;
        RECT -53.885 -39.605 -53.555 -39.275 ;
        RECT -53.885 -40.965 -53.555 -40.635 ;
        RECT -53.885 -42.325 -53.555 -41.995 ;
        RECT -53.885 -43.685 -53.555 -43.355 ;
        RECT -53.885 -45.045 -53.555 -44.715 ;
        RECT -53.885 -46.405 -53.555 -46.075 ;
        RECT -53.885 -47.765 -53.555 -47.435 ;
        RECT -53.885 -49.125 -53.555 -48.795 ;
        RECT -53.885 -50.485 -53.555 -50.155 ;
        RECT -53.885 -51.845 -53.555 -51.515 ;
        RECT -53.885 -53.205 -53.555 -52.875 ;
        RECT -53.885 -54.565 -53.555 -54.235 ;
        RECT -53.885 -55.925 -53.555 -55.595 ;
        RECT -53.885 -57.285 -53.555 -56.955 ;
        RECT -53.885 -58.645 -53.555 -58.315 ;
        RECT -53.885 -60.005 -53.555 -59.675 ;
        RECT -53.885 -61.365 -53.555 -61.035 ;
    END
    PORT
      LAYER met3 ;
        RECT -63.405 129.8 -63.075 130.93 ;
        RECT -63.405 127.675 -63.075 128.005 ;
        RECT -63.405 126.315 -63.075 126.645 ;
        RECT -63.405 124.955 -63.075 125.285 ;
        RECT -63.405 123.595 -63.075 123.925 ;
        RECT -63.405 122.235 -63.075 122.565 ;
        RECT -63.405 120.875 -63.075 121.205 ;
        RECT -63.405 119.515 -63.075 119.845 ;
        RECT -63.405 118.155 -63.075 118.485 ;
        RECT -63.405 116.795 -63.075 117.125 ;
        RECT -63.405 115.435 -63.075 115.765 ;
        RECT -63.405 114.075 -63.075 114.405 ;
        RECT -63.405 112.715 -63.075 113.045 ;
        RECT -63.405 111.355 -63.075 111.685 ;
        RECT -63.405 109.995 -63.075 110.325 ;
        RECT -63.405 108.635 -63.075 108.965 ;
        RECT -63.405 107.275 -63.075 107.605 ;
        RECT -63.405 105.915 -63.075 106.245 ;
        RECT -63.405 104.555 -63.075 104.885 ;
        RECT -63.405 103.195 -63.075 103.525 ;
        RECT -63.405 101.835 -63.075 102.165 ;
        RECT -63.405 100.475 -63.075 100.805 ;
        RECT -63.405 99.115 -63.075 99.445 ;
        RECT -63.405 97.755 -63.075 98.085 ;
        RECT -63.405 96.395 -63.075 96.725 ;
        RECT -63.405 95.035 -63.075 95.365 ;
        RECT -63.405 93.675 -63.075 94.005 ;
        RECT -63.405 92.315 -63.075 92.645 ;
        RECT -63.405 90.955 -63.075 91.285 ;
        RECT -63.405 89.595 -63.075 89.925 ;
        RECT -63.405 88.235 -63.075 88.565 ;
        RECT -63.405 86.875 -63.075 87.205 ;
        RECT -63.405 85.515 -63.075 85.845 ;
        RECT -63.405 84.155 -63.075 84.485 ;
        RECT -63.405 82.795 -63.075 83.125 ;
        RECT -63.405 81.435 -63.075 81.765 ;
        RECT -63.405 80.075 -63.075 80.405 ;
        RECT -63.405 78.715 -63.075 79.045 ;
        RECT -63.405 77.355 -63.075 77.685 ;
        RECT -63.405 75.995 -63.075 76.325 ;
        RECT -63.405 74.635 -63.075 74.965 ;
        RECT -63.405 73.275 -63.075 73.605 ;
        RECT -63.405 71.915 -63.075 72.245 ;
        RECT -63.405 70.555 -63.075 70.885 ;
        RECT -63.405 69.195 -63.075 69.525 ;
        RECT -63.405 67.835 -63.075 68.165 ;
        RECT -63.405 66.475 -63.075 66.805 ;
        RECT -63.405 65.115 -63.075 65.445 ;
        RECT -63.405 63.755 -63.075 64.085 ;
        RECT -63.405 62.395 -63.075 62.725 ;
        RECT -63.405 61.035 -63.075 61.365 ;
        RECT -63.405 59.675 -63.075 60.005 ;
        RECT -63.405 58.315 -63.075 58.645 ;
        RECT -63.405 56.955 -63.075 57.285 ;
        RECT -63.405 55.595 -63.075 55.925 ;
        RECT -63.405 54.235 -63.075 54.565 ;
        RECT -63.405 52.875 -63.075 53.205 ;
        RECT -63.405 51.515 -63.075 51.845 ;
        RECT -63.405 50.155 -63.075 50.485 ;
        RECT -63.405 48.795 -63.075 49.125 ;
        RECT -63.405 47.435 -63.075 47.765 ;
        RECT -63.405 46.075 -63.075 46.405 ;
        RECT -63.405 44.715 -63.075 45.045 ;
        RECT -63.405 43.355 -63.075 43.685 ;
        RECT -63.405 41.995 -63.075 42.325 ;
        RECT -63.405 40.635 -63.075 40.965 ;
        RECT -63.405 39.275 -63.075 39.605 ;
        RECT -63.405 37.915 -63.075 38.245 ;
        RECT -63.405 36.555 -63.075 36.885 ;
        RECT -63.405 35.195 -63.075 35.525 ;
        RECT -63.405 33.835 -63.075 34.165 ;
        RECT -63.405 32.475 -63.075 32.805 ;
        RECT -63.405 31.115 -63.075 31.445 ;
        RECT -63.405 29.755 -63.075 30.085 ;
        RECT -63.405 28.395 -63.075 28.725 ;
        RECT -63.405 27.035 -63.075 27.365 ;
        RECT -63.405 25.675 -63.075 26.005 ;
        RECT -63.405 24.315 -63.075 24.645 ;
        RECT -63.405 22.955 -63.075 23.285 ;
        RECT -63.405 21.595 -63.075 21.925 ;
        RECT -63.405 20.235 -63.075 20.565 ;
        RECT -63.405 18.875 -63.075 19.205 ;
        RECT -63.405 17.515 -63.075 17.845 ;
        RECT -63.405 16.155 -63.075 16.485 ;
        RECT -63.405 14.795 -63.075 15.125 ;
        RECT -63.405 13.435 -63.075 13.765 ;
        RECT -63.405 12.075 -63.075 12.405 ;
        RECT -63.405 10.715 -63.075 11.045 ;
        RECT -63.405 9.355 -63.075 9.685 ;
        RECT -63.405 7.995 -63.075 8.325 ;
        RECT -63.405 6.635 -63.075 6.965 ;
        RECT -63.405 5.275 -63.075 5.605 ;
        RECT -63.405 3.915 -63.075 4.245 ;
        RECT -63.405 2.555 -63.075 2.885 ;
        RECT -63.405 1.195 -63.075 1.525 ;
        RECT -63.405 -0.165 -63.075 0.165 ;
        RECT -63.405 -1.525 -63.075 -1.195 ;
        RECT -63.405 -2.885 -63.075 -2.555 ;
        RECT -63.405 -4.245 -63.075 -3.915 ;
        RECT -63.405 -5.605 -63.075 -5.275 ;
        RECT -63.405 -6.965 -63.075 -6.635 ;
        RECT -63.405 -8.325 -63.075 -7.995 ;
        RECT -63.405 -9.685 -63.075 -9.355 ;
        RECT -63.405 -11.045 -63.075 -10.715 ;
        RECT -63.405 -12.405 -63.075 -12.075 ;
        RECT -63.405 -13.765 -63.075 -13.435 ;
        RECT -63.405 -15.125 -63.075 -14.795 ;
        RECT -63.405 -16.485 -63.075 -16.155 ;
        RECT -63.405 -17.845 -63.075 -17.515 ;
        RECT -63.405 -19.205 -63.075 -18.875 ;
        RECT -63.405 -20.565 -63.075 -20.235 ;
        RECT -63.405 -21.925 -63.075 -21.595 ;
        RECT -63.405 -23.285 -63.075 -22.955 ;
        RECT -63.405 -24.645 -63.075 -24.315 ;
        RECT -63.405 -26.005 -63.075 -25.675 ;
        RECT -63.405 -27.365 -63.075 -27.035 ;
        RECT -63.405 -28.725 -63.075 -28.395 ;
        RECT -63.405 -30.085 -63.075 -29.755 ;
        RECT -63.405 -31.445 -63.075 -31.115 ;
        RECT -63.405 -32.805 -63.075 -32.475 ;
        RECT -63.405 -34.165 -63.075 -33.835 ;
        RECT -63.405 -35.525 -63.075 -35.195 ;
        RECT -63.405 -36.885 -63.075 -36.555 ;
        RECT -63.405 -38.245 -63.075 -37.915 ;
        RECT -63.405 -39.605 -63.075 -39.275 ;
        RECT -63.405 -40.965 -63.075 -40.635 ;
        RECT -63.405 -42.325 -63.075 -41.995 ;
        RECT -63.405 -43.685 -63.075 -43.355 ;
        RECT -63.405 -45.045 -63.075 -44.715 ;
        RECT -63.405 -46.405 -63.075 -46.075 ;
        RECT -63.405 -47.765 -63.075 -47.435 ;
        RECT -63.405 -49.125 -63.075 -48.795 ;
        RECT -63.405 -50.485 -63.075 -50.155 ;
        RECT -63.405 -51.845 -63.075 -51.515 ;
        RECT -63.405 -53.205 -63.075 -52.875 ;
        RECT -63.405 -54.565 -63.075 -54.235 ;
        RECT -63.405 -55.925 -63.075 -55.595 ;
        RECT -63.405 -57.285 -63.075 -56.955 ;
        RECT -63.405 -58.645 -63.075 -58.315 ;
        RECT -63.405 -60.005 -63.075 -59.675 ;
        RECT -63.405 -61.365 -63.075 -61.035 ;
        RECT -63.405 -62.725 -63.075 -62.395 ;
        RECT -63.405 -64.085 -63.075 -63.755 ;
        RECT -63.405 -65.445 -63.075 -65.115 ;
        RECT -63.405 -66.805 -63.075 -66.475 ;
        RECT -63.405 -68.165 -63.075 -67.835 ;
        RECT -63.405 -69.525 -63.075 -69.195 ;
        RECT -63.405 -70.885 -63.075 -70.555 ;
        RECT -63.405 -72.245 -63.075 -71.915 ;
        RECT -63.405 -73.605 -63.075 -73.275 ;
        RECT -63.405 -74.965 -63.075 -74.635 ;
        RECT -63.405 -76.325 -63.075 -75.995 ;
        RECT -63.405 -77.685 -63.075 -77.355 ;
        RECT -63.405 -79.045 -63.075 -78.715 ;
        RECT -63.405 -80.405 -63.075 -80.075 ;
        RECT -63.405 -81.765 -63.075 -81.435 ;
        RECT -63.405 -83.125 -63.075 -82.795 ;
        RECT -63.405 -84.485 -63.075 -84.155 ;
        RECT -63.405 -85.845 -63.075 -85.515 ;
        RECT -63.405 -87.205 -63.075 -86.875 ;
        RECT -63.405 -88.565 -63.075 -88.235 ;
        RECT -63.405 -89.925 -63.075 -89.595 ;
        RECT -63.405 -91.285 -63.075 -90.955 ;
        RECT -63.405 -92.645 -63.075 -92.315 ;
        RECT -63.405 -94.005 -63.075 -93.675 ;
        RECT -63.405 -95.365 -63.075 -95.035 ;
        RECT -63.405 -96.725 -63.075 -96.395 ;
        RECT -63.405 -98.085 -63.075 -97.755 ;
        RECT -63.405 -99.445 -63.075 -99.115 ;
        RECT -63.405 -100.805 -63.075 -100.475 ;
        RECT -63.405 -102.165 -63.075 -101.835 ;
        RECT -63.405 -103.525 -63.075 -103.195 ;
        RECT -63.405 -104.885 -63.075 -104.555 ;
        RECT -63.405 -106.245 -63.075 -105.915 ;
        RECT -63.405 -107.605 -63.075 -107.275 ;
        RECT -63.405 -108.965 -63.075 -108.635 ;
        RECT -63.405 -110.325 -63.075 -109.995 ;
        RECT -63.405 -111.685 -63.075 -111.355 ;
        RECT -63.405 -113.045 -63.075 -112.715 ;
        RECT -63.405 -114.405 -63.075 -114.075 ;
        RECT -63.405 -115.765 -63.075 -115.435 ;
        RECT -63.405 -117.125 -63.075 -116.795 ;
        RECT -63.405 -118.485 -63.075 -118.155 ;
        RECT -63.405 -119.845 -63.075 -119.515 ;
        RECT -63.405 -121.205 -63.075 -120.875 ;
        RECT -63.405 -122.565 -63.075 -122.235 ;
        RECT -63.405 -123.925 -63.075 -123.595 ;
        RECT -63.405 -125.285 -63.075 -124.955 ;
        RECT -63.405 -126.645 -63.075 -126.315 ;
        RECT -63.405 -128.005 -63.075 -127.675 ;
        RECT -63.405 -129.365 -63.075 -129.035 ;
        RECT -63.405 -130.725 -63.075 -130.395 ;
        RECT -63.405 -132.085 -63.075 -131.755 ;
        RECT -63.405 -133.445 -63.075 -133.115 ;
        RECT -63.405 -134.805 -63.075 -134.475 ;
        RECT -63.405 -136.165 -63.075 -135.835 ;
        RECT -63.405 -137.525 -63.075 -137.195 ;
        RECT -63.405 -138.885 -63.075 -138.555 ;
        RECT -63.405 -140.245 -63.075 -139.915 ;
        RECT -63.405 -141.605 -63.075 -141.275 ;
        RECT -63.405 -142.965 -63.075 -142.635 ;
        RECT -63.405 -144.325 -63.075 -143.995 ;
        RECT -63.405 -145.685 -63.075 -145.355 ;
        RECT -63.405 -147.045 -63.075 -146.715 ;
        RECT -63.405 -148.405 -63.075 -148.075 ;
        RECT -63.405 -149.765 -63.075 -149.435 ;
        RECT -63.405 -151.125 -63.075 -150.795 ;
        RECT -63.405 -152.485 -63.075 -152.155 ;
        RECT -63.405 -153.845 -63.075 -153.515 ;
        RECT -63.405 -155.205 -63.075 -154.875 ;
        RECT -63.405 -156.565 -63.075 -156.235 ;
        RECT -63.405 -157.925 -63.075 -157.595 ;
        RECT -63.405 -159.285 -63.075 -158.955 ;
        RECT -63.405 -160.645 -63.075 -160.315 ;
        RECT -63.405 -162.005 -63.075 -161.675 ;
        RECT -63.405 -163.365 -63.075 -163.035 ;
        RECT -63.405 -164.725 -63.075 -164.395 ;
        RECT -63.405 -166.085 -63.075 -165.755 ;
        RECT -63.405 -167.445 -63.075 -167.115 ;
        RECT -63.405 -168.805 -63.075 -168.475 ;
        RECT -63.405 -170.165 -63.075 -169.835 ;
        RECT -63.405 -171.525 -63.075 -171.195 ;
        RECT -63.405 -172.885 -63.075 -172.555 ;
        RECT -63.405 -174.245 -63.075 -173.915 ;
        RECT -63.405 -175.605 -63.075 -175.275 ;
        RECT -63.405 -176.965 -63.075 -176.635 ;
        RECT -63.405 -178.325 -63.075 -177.995 ;
        RECT -63.405 -179.685 -63.075 -179.355 ;
        RECT -63.405 -181.045 -63.075 -180.715 ;
        RECT -63.405 -182.405 -63.075 -182.075 ;
        RECT -63.405 -183.765 -63.075 -183.435 ;
        RECT -63.405 -185.125 -63.075 -184.795 ;
        RECT -63.405 -186.485 -63.075 -186.155 ;
        RECT -63.405 -187.845 -63.075 -187.515 ;
        RECT -63.405 -189.205 -63.075 -188.875 ;
        RECT -63.405 -190.565 -63.075 -190.235 ;
        RECT -63.405 -191.925 -63.075 -191.595 ;
        RECT -63.405 -193.285 -63.075 -192.955 ;
        RECT -63.405 -194.645 -63.075 -194.315 ;
        RECT -63.405 -196.005 -63.075 -195.675 ;
        RECT -63.405 -197.365 -63.075 -197.035 ;
        RECT -63.405 -198.725 -63.075 -198.395 ;
        RECT -63.405 -200.085 -63.075 -199.755 ;
        RECT -63.405 -201.445 -63.075 -201.115 ;
        RECT -63.405 -202.805 -63.075 -202.475 ;
        RECT -63.405 -204.165 -63.075 -203.835 ;
        RECT -63.405 -205.525 -63.075 -205.195 ;
        RECT -63.405 -208.245 -63.075 -207.915 ;
        RECT -63.405 -210.965 -63.075 -210.635 ;
        RECT -63.405 -212.325 -63.075 -211.995 ;
        RECT -63.405 -213.625 -63.075 -213.295 ;
        RECT -63.405 -215.045 -63.075 -214.715 ;
        RECT -63.405 -216.405 -63.075 -216.075 ;
        RECT -63.405 -217.765 -63.075 -217.435 ;
        RECT -63.405 -219.125 -63.075 -218.795 ;
        RECT -63.405 -221.37 -63.075 -220.24 ;
        RECT -63.4 -221.485 -63.08 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -62.045 129.8 -61.715 130.93 ;
        RECT -62.045 127.675 -61.715 128.005 ;
        RECT -62.045 126.315 -61.715 126.645 ;
        RECT -62.045 124.955 -61.715 125.285 ;
        RECT -62.045 123.595 -61.715 123.925 ;
        RECT -62.045 122.235 -61.715 122.565 ;
        RECT -62.045 120.875 -61.715 121.205 ;
        RECT -62.045 119.515 -61.715 119.845 ;
        RECT -62.045 118.155 -61.715 118.485 ;
        RECT -62.045 116.795 -61.715 117.125 ;
        RECT -62.045 115.435 -61.715 115.765 ;
        RECT -62.045 114.075 -61.715 114.405 ;
        RECT -62.045 112.715 -61.715 113.045 ;
        RECT -62.045 111.355 -61.715 111.685 ;
        RECT -62.045 109.995 -61.715 110.325 ;
        RECT -62.045 108.635 -61.715 108.965 ;
        RECT -62.045 107.275 -61.715 107.605 ;
        RECT -62.045 105.915 -61.715 106.245 ;
        RECT -62.045 104.555 -61.715 104.885 ;
        RECT -62.045 103.195 -61.715 103.525 ;
        RECT -62.045 101.835 -61.715 102.165 ;
        RECT -62.045 100.475 -61.715 100.805 ;
        RECT -62.045 99.115 -61.715 99.445 ;
        RECT -62.045 97.755 -61.715 98.085 ;
        RECT -62.045 96.395 -61.715 96.725 ;
        RECT -62.045 95.035 -61.715 95.365 ;
        RECT -62.045 93.675 -61.715 94.005 ;
        RECT -62.045 92.315 -61.715 92.645 ;
        RECT -62.045 90.955 -61.715 91.285 ;
        RECT -62.045 89.595 -61.715 89.925 ;
        RECT -62.045 88.235 -61.715 88.565 ;
        RECT -62.045 86.875 -61.715 87.205 ;
        RECT -62.045 85.515 -61.715 85.845 ;
        RECT -62.045 84.155 -61.715 84.485 ;
        RECT -62.045 82.795 -61.715 83.125 ;
        RECT -62.045 81.435 -61.715 81.765 ;
        RECT -62.045 80.075 -61.715 80.405 ;
        RECT -62.045 78.715 -61.715 79.045 ;
        RECT -62.045 77.355 -61.715 77.685 ;
        RECT -62.045 75.995 -61.715 76.325 ;
        RECT -62.045 74.635 -61.715 74.965 ;
        RECT -62.045 73.275 -61.715 73.605 ;
        RECT -62.045 71.915 -61.715 72.245 ;
        RECT -62.045 70.555 -61.715 70.885 ;
        RECT -62.045 69.195 -61.715 69.525 ;
        RECT -62.045 67.835 -61.715 68.165 ;
        RECT -62.045 66.475 -61.715 66.805 ;
        RECT -62.045 65.115 -61.715 65.445 ;
        RECT -62.045 63.755 -61.715 64.085 ;
        RECT -62.045 62.395 -61.715 62.725 ;
        RECT -62.045 61.035 -61.715 61.365 ;
        RECT -62.045 59.675 -61.715 60.005 ;
        RECT -62.045 58.315 -61.715 58.645 ;
        RECT -62.045 56.955 -61.715 57.285 ;
        RECT -62.045 55.595 -61.715 55.925 ;
        RECT -62.045 54.235 -61.715 54.565 ;
        RECT -62.045 52.875 -61.715 53.205 ;
        RECT -62.045 51.515 -61.715 51.845 ;
        RECT -62.045 50.155 -61.715 50.485 ;
        RECT -62.045 48.795 -61.715 49.125 ;
        RECT -62.045 47.435 -61.715 47.765 ;
        RECT -62.045 46.075 -61.715 46.405 ;
        RECT -62.045 44.715 -61.715 45.045 ;
        RECT -62.045 43.355 -61.715 43.685 ;
        RECT -62.045 41.995 -61.715 42.325 ;
        RECT -62.045 40.635 -61.715 40.965 ;
        RECT -62.045 39.275 -61.715 39.605 ;
        RECT -62.045 37.915 -61.715 38.245 ;
        RECT -62.045 36.555 -61.715 36.885 ;
        RECT -62.045 35.195 -61.715 35.525 ;
        RECT -62.045 33.835 -61.715 34.165 ;
        RECT -62.045 32.475 -61.715 32.805 ;
        RECT -62.045 31.115 -61.715 31.445 ;
        RECT -62.045 29.755 -61.715 30.085 ;
        RECT -62.045 28.395 -61.715 28.725 ;
        RECT -62.045 27.035 -61.715 27.365 ;
        RECT -62.045 25.675 -61.715 26.005 ;
        RECT -62.045 24.315 -61.715 24.645 ;
        RECT -62.045 22.955 -61.715 23.285 ;
        RECT -62.045 21.595 -61.715 21.925 ;
        RECT -62.045 20.235 -61.715 20.565 ;
        RECT -62.045 18.875 -61.715 19.205 ;
        RECT -62.045 17.515 -61.715 17.845 ;
        RECT -62.045 16.155 -61.715 16.485 ;
        RECT -62.045 14.795 -61.715 15.125 ;
        RECT -62.045 13.435 -61.715 13.765 ;
        RECT -62.045 12.075 -61.715 12.405 ;
        RECT -62.045 10.715 -61.715 11.045 ;
        RECT -62.045 9.355 -61.715 9.685 ;
        RECT -62.045 7.995 -61.715 8.325 ;
        RECT -62.045 6.635 -61.715 6.965 ;
        RECT -62.045 5.275 -61.715 5.605 ;
        RECT -62.045 3.915 -61.715 4.245 ;
        RECT -62.045 2.555 -61.715 2.885 ;
        RECT -62.045 1.195 -61.715 1.525 ;
        RECT -62.045 -0.165 -61.715 0.165 ;
        RECT -62.045 -1.525 -61.715 -1.195 ;
        RECT -62.045 -2.885 -61.715 -2.555 ;
        RECT -62.045 -4.245 -61.715 -3.915 ;
        RECT -62.045 -5.605 -61.715 -5.275 ;
        RECT -62.045 -6.965 -61.715 -6.635 ;
        RECT -62.045 -8.325 -61.715 -7.995 ;
        RECT -62.045 -9.685 -61.715 -9.355 ;
        RECT -62.045 -11.045 -61.715 -10.715 ;
        RECT -62.045 -12.405 -61.715 -12.075 ;
        RECT -62.045 -13.765 -61.715 -13.435 ;
        RECT -62.045 -15.125 -61.715 -14.795 ;
        RECT -62.045 -16.485 -61.715 -16.155 ;
        RECT -62.045 -17.845 -61.715 -17.515 ;
        RECT -62.045 -19.205 -61.715 -18.875 ;
        RECT -62.045 -20.565 -61.715 -20.235 ;
        RECT -62.045 -21.925 -61.715 -21.595 ;
        RECT -62.045 -23.285 -61.715 -22.955 ;
        RECT -62.045 -24.645 -61.715 -24.315 ;
        RECT -62.045 -26.005 -61.715 -25.675 ;
        RECT -62.045 -27.365 -61.715 -27.035 ;
        RECT -62.045 -28.725 -61.715 -28.395 ;
        RECT -62.045 -30.085 -61.715 -29.755 ;
        RECT -62.045 -31.445 -61.715 -31.115 ;
        RECT -62.045 -32.805 -61.715 -32.475 ;
        RECT -62.045 -34.165 -61.715 -33.835 ;
        RECT -62.045 -35.525 -61.715 -35.195 ;
        RECT -62.045 -36.885 -61.715 -36.555 ;
        RECT -62.045 -38.245 -61.715 -37.915 ;
        RECT -62.045 -39.605 -61.715 -39.275 ;
        RECT -62.045 -40.965 -61.715 -40.635 ;
        RECT -62.045 -42.325 -61.715 -41.995 ;
        RECT -62.045 -43.685 -61.715 -43.355 ;
        RECT -62.045 -45.045 -61.715 -44.715 ;
        RECT -62.045 -46.405 -61.715 -46.075 ;
        RECT -62.045 -47.765 -61.715 -47.435 ;
        RECT -62.045 -49.125 -61.715 -48.795 ;
        RECT -62.045 -50.485 -61.715 -50.155 ;
        RECT -62.045 -51.845 -61.715 -51.515 ;
        RECT -62.045 -53.205 -61.715 -52.875 ;
        RECT -62.045 -54.565 -61.715 -54.235 ;
        RECT -62.045 -55.925 -61.715 -55.595 ;
        RECT -62.045 -57.285 -61.715 -56.955 ;
        RECT -62.045 -58.645 -61.715 -58.315 ;
        RECT -62.045 -60.005 -61.715 -59.675 ;
        RECT -62.045 -61.365 -61.715 -61.035 ;
        RECT -62.045 -62.725 -61.715 -62.395 ;
        RECT -62.045 -64.085 -61.715 -63.755 ;
        RECT -62.045 -65.445 -61.715 -65.115 ;
        RECT -62.045 -66.805 -61.715 -66.475 ;
        RECT -62.045 -68.165 -61.715 -67.835 ;
        RECT -62.045 -69.525 -61.715 -69.195 ;
        RECT -62.045 -70.885 -61.715 -70.555 ;
        RECT -62.045 -72.245 -61.715 -71.915 ;
        RECT -62.045 -73.605 -61.715 -73.275 ;
        RECT -62.045 -74.965 -61.715 -74.635 ;
        RECT -62.045 -76.325 -61.715 -75.995 ;
        RECT -62.045 -77.685 -61.715 -77.355 ;
        RECT -62.045 -79.045 -61.715 -78.715 ;
        RECT -62.045 -80.405 -61.715 -80.075 ;
        RECT -62.045 -81.765 -61.715 -81.435 ;
        RECT -62.045 -83.125 -61.715 -82.795 ;
        RECT -62.045 -84.485 -61.715 -84.155 ;
        RECT -62.045 -85.845 -61.715 -85.515 ;
        RECT -62.045 -87.205 -61.715 -86.875 ;
        RECT -62.045 -88.565 -61.715 -88.235 ;
        RECT -62.045 -89.925 -61.715 -89.595 ;
        RECT -62.045 -91.285 -61.715 -90.955 ;
        RECT -62.045 -92.645 -61.715 -92.315 ;
        RECT -62.045 -94.005 -61.715 -93.675 ;
        RECT -62.045 -95.365 -61.715 -95.035 ;
        RECT -62.045 -96.725 -61.715 -96.395 ;
        RECT -62.045 -98.085 -61.715 -97.755 ;
        RECT -62.045 -99.445 -61.715 -99.115 ;
        RECT -62.045 -100.805 -61.715 -100.475 ;
        RECT -62.045 -102.165 -61.715 -101.835 ;
        RECT -62.045 -103.525 -61.715 -103.195 ;
        RECT -62.045 -104.885 -61.715 -104.555 ;
        RECT -62.045 -106.245 -61.715 -105.915 ;
        RECT -62.045 -107.605 -61.715 -107.275 ;
        RECT -62.045 -108.965 -61.715 -108.635 ;
        RECT -62.045 -110.325 -61.715 -109.995 ;
        RECT -62.045 -111.685 -61.715 -111.355 ;
        RECT -62.045 -113.045 -61.715 -112.715 ;
        RECT -62.045 -114.405 -61.715 -114.075 ;
        RECT -62.045 -115.765 -61.715 -115.435 ;
        RECT -62.045 -117.125 -61.715 -116.795 ;
        RECT -62.045 -118.485 -61.715 -118.155 ;
        RECT -62.045 -119.845 -61.715 -119.515 ;
        RECT -62.045 -121.205 -61.715 -120.875 ;
        RECT -62.045 -122.565 -61.715 -122.235 ;
        RECT -62.045 -123.925 -61.715 -123.595 ;
        RECT -62.045 -125.285 -61.715 -124.955 ;
        RECT -62.045 -126.645 -61.715 -126.315 ;
        RECT -62.045 -128.005 -61.715 -127.675 ;
        RECT -62.045 -129.365 -61.715 -129.035 ;
        RECT -62.045 -130.725 -61.715 -130.395 ;
        RECT -62.045 -132.085 -61.715 -131.755 ;
        RECT -62.045 -133.445 -61.715 -133.115 ;
        RECT -62.045 -134.805 -61.715 -134.475 ;
        RECT -62.045 -136.165 -61.715 -135.835 ;
        RECT -62.045 -137.525 -61.715 -137.195 ;
        RECT -62.045 -138.885 -61.715 -138.555 ;
        RECT -62.045 -140.245 -61.715 -139.915 ;
        RECT -62.045 -141.605 -61.715 -141.275 ;
        RECT -62.045 -142.965 -61.715 -142.635 ;
        RECT -62.045 -144.325 -61.715 -143.995 ;
        RECT -62.045 -145.685 -61.715 -145.355 ;
        RECT -62.045 -147.045 -61.715 -146.715 ;
        RECT -62.045 -148.405 -61.715 -148.075 ;
        RECT -62.045 -149.765 -61.715 -149.435 ;
        RECT -62.045 -151.125 -61.715 -150.795 ;
        RECT -62.045 -152.485 -61.715 -152.155 ;
        RECT -62.045 -153.845 -61.715 -153.515 ;
        RECT -62.045 -155.205 -61.715 -154.875 ;
        RECT -62.045 -156.565 -61.715 -156.235 ;
        RECT -62.045 -157.925 -61.715 -157.595 ;
        RECT -62.045 -159.285 -61.715 -158.955 ;
        RECT -62.045 -160.645 -61.715 -160.315 ;
        RECT -62.045 -162.005 -61.715 -161.675 ;
        RECT -62.045 -163.365 -61.715 -163.035 ;
        RECT -62.045 -164.725 -61.715 -164.395 ;
        RECT -62.045 -166.085 -61.715 -165.755 ;
        RECT -62.045 -167.445 -61.715 -167.115 ;
        RECT -62.045 -168.805 -61.715 -168.475 ;
        RECT -62.045 -170.165 -61.715 -169.835 ;
        RECT -62.045 -171.525 -61.715 -171.195 ;
        RECT -62.045 -172.885 -61.715 -172.555 ;
        RECT -62.045 -174.245 -61.715 -173.915 ;
        RECT -62.045 -175.605 -61.715 -175.275 ;
        RECT -62.045 -176.965 -61.715 -176.635 ;
        RECT -62.045 -178.325 -61.715 -177.995 ;
        RECT -62.045 -179.685 -61.715 -179.355 ;
        RECT -62.045 -181.045 -61.715 -180.715 ;
        RECT -62.045 -182.405 -61.715 -182.075 ;
        RECT -62.045 -183.765 -61.715 -183.435 ;
        RECT -62.045 -185.125 -61.715 -184.795 ;
        RECT -62.045 -186.485 -61.715 -186.155 ;
        RECT -62.045 -187.845 -61.715 -187.515 ;
        RECT -62.045 -189.205 -61.715 -188.875 ;
        RECT -62.045 -190.565 -61.715 -190.235 ;
        RECT -62.045 -191.925 -61.715 -191.595 ;
        RECT -62.045 -193.285 -61.715 -192.955 ;
        RECT -62.045 -194.645 -61.715 -194.315 ;
        RECT -62.045 -196.005 -61.715 -195.675 ;
        RECT -62.045 -197.365 -61.715 -197.035 ;
        RECT -62.045 -198.725 -61.715 -198.395 ;
        RECT -62.045 -200.085 -61.715 -199.755 ;
        RECT -62.045 -201.445 -61.715 -201.115 ;
        RECT -62.045 -202.805 -61.715 -202.475 ;
        RECT -62.045 -204.165 -61.715 -203.835 ;
        RECT -62.045 -205.525 -61.715 -205.195 ;
        RECT -62.045 -208.245 -61.715 -207.915 ;
        RECT -62.045 -210.965 -61.715 -210.635 ;
        RECT -62.045 -212.325 -61.715 -211.995 ;
        RECT -62.045 -213.625 -61.715 -213.295 ;
        RECT -62.045 -215.045 -61.715 -214.715 ;
        RECT -62.045 -216.405 -61.715 -216.075 ;
        RECT -62.045 -217.765 -61.715 -217.435 ;
        RECT -62.045 -219.125 -61.715 -218.795 ;
        RECT -62.045 -221.37 -61.715 -220.24 ;
        RECT -62.04 -221.485 -61.72 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -60.685 129.8 -60.355 130.93 ;
        RECT -60.685 127.675 -60.355 128.005 ;
        RECT -60.685 126.315 -60.355 126.645 ;
        RECT -60.685 124.955 -60.355 125.285 ;
        RECT -60.685 123.595 -60.355 123.925 ;
        RECT -60.685 122.235 -60.355 122.565 ;
        RECT -60.685 120.875 -60.355 121.205 ;
        RECT -60.685 119.515 -60.355 119.845 ;
        RECT -60.685 118.155 -60.355 118.485 ;
        RECT -60.685 116.795 -60.355 117.125 ;
        RECT -60.685 115.435 -60.355 115.765 ;
        RECT -60.685 114.075 -60.355 114.405 ;
        RECT -60.685 112.715 -60.355 113.045 ;
        RECT -60.685 111.355 -60.355 111.685 ;
        RECT -60.685 109.995 -60.355 110.325 ;
        RECT -60.685 108.635 -60.355 108.965 ;
        RECT -60.685 107.275 -60.355 107.605 ;
        RECT -60.685 105.915 -60.355 106.245 ;
        RECT -60.685 104.555 -60.355 104.885 ;
        RECT -60.685 103.195 -60.355 103.525 ;
        RECT -60.685 101.835 -60.355 102.165 ;
        RECT -60.685 100.475 -60.355 100.805 ;
        RECT -60.685 99.115 -60.355 99.445 ;
        RECT -60.685 97.755 -60.355 98.085 ;
        RECT -60.685 96.395 -60.355 96.725 ;
        RECT -60.685 95.035 -60.355 95.365 ;
        RECT -60.685 93.675 -60.355 94.005 ;
        RECT -60.685 92.315 -60.355 92.645 ;
        RECT -60.685 90.955 -60.355 91.285 ;
        RECT -60.685 89.595 -60.355 89.925 ;
        RECT -60.685 88.235 -60.355 88.565 ;
        RECT -60.685 86.875 -60.355 87.205 ;
        RECT -60.685 85.515 -60.355 85.845 ;
        RECT -60.685 84.155 -60.355 84.485 ;
        RECT -60.685 82.795 -60.355 83.125 ;
        RECT -60.685 81.435 -60.355 81.765 ;
        RECT -60.685 80.075 -60.355 80.405 ;
        RECT -60.685 78.715 -60.355 79.045 ;
        RECT -60.685 77.355 -60.355 77.685 ;
        RECT -60.685 75.995 -60.355 76.325 ;
        RECT -60.685 74.635 -60.355 74.965 ;
        RECT -60.685 73.275 -60.355 73.605 ;
        RECT -60.685 71.915 -60.355 72.245 ;
        RECT -60.685 70.555 -60.355 70.885 ;
        RECT -60.685 69.195 -60.355 69.525 ;
        RECT -60.685 67.835 -60.355 68.165 ;
        RECT -60.685 66.475 -60.355 66.805 ;
        RECT -60.685 65.115 -60.355 65.445 ;
        RECT -60.685 63.755 -60.355 64.085 ;
        RECT -60.685 62.395 -60.355 62.725 ;
        RECT -60.685 61.035 -60.355 61.365 ;
        RECT -60.685 59.675 -60.355 60.005 ;
        RECT -60.685 58.315 -60.355 58.645 ;
        RECT -60.685 56.955 -60.355 57.285 ;
        RECT -60.685 55.595 -60.355 55.925 ;
        RECT -60.685 54.235 -60.355 54.565 ;
        RECT -60.685 52.875 -60.355 53.205 ;
        RECT -60.685 51.515 -60.355 51.845 ;
        RECT -60.685 50.155 -60.355 50.485 ;
        RECT -60.685 48.795 -60.355 49.125 ;
        RECT -60.685 47.435 -60.355 47.765 ;
        RECT -60.685 46.075 -60.355 46.405 ;
        RECT -60.685 44.715 -60.355 45.045 ;
        RECT -60.685 43.355 -60.355 43.685 ;
        RECT -60.685 41.995 -60.355 42.325 ;
        RECT -60.685 40.635 -60.355 40.965 ;
        RECT -60.685 39.275 -60.355 39.605 ;
        RECT -60.685 37.915 -60.355 38.245 ;
        RECT -60.685 36.555 -60.355 36.885 ;
        RECT -60.685 35.195 -60.355 35.525 ;
        RECT -60.685 33.835 -60.355 34.165 ;
        RECT -60.685 32.475 -60.355 32.805 ;
        RECT -60.685 31.115 -60.355 31.445 ;
        RECT -60.685 29.755 -60.355 30.085 ;
        RECT -60.685 28.395 -60.355 28.725 ;
        RECT -60.685 27.035 -60.355 27.365 ;
        RECT -60.685 25.675 -60.355 26.005 ;
        RECT -60.685 24.315 -60.355 24.645 ;
        RECT -60.685 22.955 -60.355 23.285 ;
        RECT -60.685 21.595 -60.355 21.925 ;
        RECT -60.685 20.235 -60.355 20.565 ;
        RECT -60.685 18.875 -60.355 19.205 ;
        RECT -60.685 17.515 -60.355 17.845 ;
        RECT -60.685 16.155 -60.355 16.485 ;
        RECT -60.685 14.795 -60.355 15.125 ;
        RECT -60.685 13.435 -60.355 13.765 ;
        RECT -60.685 12.075 -60.355 12.405 ;
        RECT -60.685 10.715 -60.355 11.045 ;
        RECT -60.685 9.355 -60.355 9.685 ;
        RECT -60.685 7.995 -60.355 8.325 ;
        RECT -60.685 6.635 -60.355 6.965 ;
        RECT -60.685 5.275 -60.355 5.605 ;
        RECT -60.685 3.915 -60.355 4.245 ;
        RECT -60.685 2.555 -60.355 2.885 ;
        RECT -60.685 1.195 -60.355 1.525 ;
        RECT -60.685 -0.165 -60.355 0.165 ;
        RECT -60.685 -1.525 -60.355 -1.195 ;
        RECT -60.685 -2.885 -60.355 -2.555 ;
        RECT -60.685 -4.245 -60.355 -3.915 ;
        RECT -60.685 -5.605 -60.355 -5.275 ;
        RECT -60.685 -6.965 -60.355 -6.635 ;
        RECT -60.685 -8.325 -60.355 -7.995 ;
        RECT -60.685 -9.685 -60.355 -9.355 ;
        RECT -60.685 -11.045 -60.355 -10.715 ;
        RECT -60.685 -12.405 -60.355 -12.075 ;
        RECT -60.685 -13.765 -60.355 -13.435 ;
        RECT -60.685 -15.125 -60.355 -14.795 ;
        RECT -60.685 -16.485 -60.355 -16.155 ;
        RECT -60.685 -17.845 -60.355 -17.515 ;
        RECT -60.685 -19.205 -60.355 -18.875 ;
        RECT -60.685 -20.565 -60.355 -20.235 ;
        RECT -60.685 -21.925 -60.355 -21.595 ;
        RECT -60.685 -23.285 -60.355 -22.955 ;
        RECT -60.685 -24.645 -60.355 -24.315 ;
        RECT -60.685 -26.005 -60.355 -25.675 ;
        RECT -60.685 -27.365 -60.355 -27.035 ;
        RECT -60.685 -28.725 -60.355 -28.395 ;
        RECT -60.685 -30.085 -60.355 -29.755 ;
        RECT -60.685 -31.445 -60.355 -31.115 ;
        RECT -60.685 -32.805 -60.355 -32.475 ;
        RECT -60.685 -34.165 -60.355 -33.835 ;
        RECT -60.685 -35.525 -60.355 -35.195 ;
        RECT -60.685 -36.885 -60.355 -36.555 ;
        RECT -60.685 -38.245 -60.355 -37.915 ;
        RECT -60.685 -39.605 -60.355 -39.275 ;
        RECT -60.685 -40.965 -60.355 -40.635 ;
        RECT -60.685 -42.325 -60.355 -41.995 ;
        RECT -60.685 -43.685 -60.355 -43.355 ;
        RECT -60.685 -45.045 -60.355 -44.715 ;
        RECT -60.685 -46.405 -60.355 -46.075 ;
        RECT -60.685 -47.765 -60.355 -47.435 ;
        RECT -60.685 -49.125 -60.355 -48.795 ;
        RECT -60.685 -50.485 -60.355 -50.155 ;
        RECT -60.685 -51.845 -60.355 -51.515 ;
        RECT -60.685 -53.205 -60.355 -52.875 ;
        RECT -60.685 -54.565 -60.355 -54.235 ;
        RECT -60.685 -55.925 -60.355 -55.595 ;
        RECT -60.685 -57.285 -60.355 -56.955 ;
        RECT -60.685 -58.645 -60.355 -58.315 ;
        RECT -60.685 -60.005 -60.355 -59.675 ;
        RECT -60.685 -61.365 -60.355 -61.035 ;
        RECT -60.685 -62.725 -60.355 -62.395 ;
        RECT -60.685 -64.085 -60.355 -63.755 ;
        RECT -60.685 -65.445 -60.355 -65.115 ;
        RECT -60.685 -66.805 -60.355 -66.475 ;
        RECT -60.685 -68.165 -60.355 -67.835 ;
        RECT -60.685 -69.525 -60.355 -69.195 ;
        RECT -60.685 -70.885 -60.355 -70.555 ;
        RECT -60.685 -72.245 -60.355 -71.915 ;
        RECT -60.685 -73.605 -60.355 -73.275 ;
        RECT -60.685 -74.965 -60.355 -74.635 ;
        RECT -60.685 -76.325 -60.355 -75.995 ;
        RECT -60.685 -77.685 -60.355 -77.355 ;
        RECT -60.685 -79.045 -60.355 -78.715 ;
        RECT -60.685 -80.405 -60.355 -80.075 ;
        RECT -60.685 -81.765 -60.355 -81.435 ;
        RECT -60.685 -83.125 -60.355 -82.795 ;
        RECT -60.685 -84.485 -60.355 -84.155 ;
        RECT -60.685 -85.845 -60.355 -85.515 ;
        RECT -60.685 -87.205 -60.355 -86.875 ;
        RECT -60.685 -88.565 -60.355 -88.235 ;
        RECT -60.685 -89.925 -60.355 -89.595 ;
        RECT -60.685 -91.285 -60.355 -90.955 ;
        RECT -60.685 -92.645 -60.355 -92.315 ;
        RECT -60.685 -94.005 -60.355 -93.675 ;
        RECT -60.685 -95.365 -60.355 -95.035 ;
        RECT -60.685 -96.725 -60.355 -96.395 ;
        RECT -60.685 -98.085 -60.355 -97.755 ;
        RECT -60.685 -99.445 -60.355 -99.115 ;
        RECT -60.685 -100.805 -60.355 -100.475 ;
        RECT -60.685 -102.165 -60.355 -101.835 ;
        RECT -60.685 -103.525 -60.355 -103.195 ;
        RECT -60.685 -104.885 -60.355 -104.555 ;
        RECT -60.685 -106.245 -60.355 -105.915 ;
        RECT -60.685 -107.605 -60.355 -107.275 ;
        RECT -60.685 -108.965 -60.355 -108.635 ;
        RECT -60.685 -110.325 -60.355 -109.995 ;
        RECT -60.685 -111.685 -60.355 -111.355 ;
        RECT -60.685 -113.045 -60.355 -112.715 ;
        RECT -60.685 -114.405 -60.355 -114.075 ;
        RECT -60.685 -115.765 -60.355 -115.435 ;
        RECT -60.685 -117.125 -60.355 -116.795 ;
        RECT -60.685 -118.485 -60.355 -118.155 ;
        RECT -60.685 -119.845 -60.355 -119.515 ;
        RECT -60.685 -121.205 -60.355 -120.875 ;
        RECT -60.685 -122.565 -60.355 -122.235 ;
        RECT -60.685 -123.925 -60.355 -123.595 ;
        RECT -60.685 -125.285 -60.355 -124.955 ;
        RECT -60.685 -126.645 -60.355 -126.315 ;
        RECT -60.685 -128.005 -60.355 -127.675 ;
        RECT -60.685 -129.365 -60.355 -129.035 ;
        RECT -60.685 -130.725 -60.355 -130.395 ;
        RECT -60.685 -132.085 -60.355 -131.755 ;
        RECT -60.68 -132.76 -60.36 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -60.685 -212.325 -60.355 -211.995 ;
        RECT -60.685 -213.625 -60.355 -213.295 ;
        RECT -60.685 -215.045 -60.355 -214.715 ;
        RECT -60.685 -216.405 -60.355 -216.075 ;
        RECT -60.685 -217.765 -60.355 -217.435 ;
        RECT -60.685 -219.125 -60.355 -218.795 ;
        RECT -60.685 -221.37 -60.355 -220.24 ;
        RECT -60.68 -221.485 -60.36 -211.995 ;
    END
    PORT
      LAYER met3 ;
        RECT -59.325 -60.005 -58.995 -59.675 ;
        RECT -59.325 -61.365 -58.995 -61.035 ;
        RECT -59.325 -62.725 -58.995 -62.395 ;
        RECT -59.325 -64.085 -58.995 -63.755 ;
        RECT -59.325 -65.445 -58.995 -65.115 ;
        RECT -59.325 -66.805 -58.995 -66.475 ;
        RECT -59.325 -68.165 -58.995 -67.835 ;
        RECT -59.325 -69.525 -58.995 -69.195 ;
        RECT -59.325 -70.885 -58.995 -70.555 ;
        RECT -59.325 -72.245 -58.995 -71.915 ;
        RECT -59.325 -73.605 -58.995 -73.275 ;
        RECT -59.325 -74.965 -58.995 -74.635 ;
        RECT -59.325 -76.325 -58.995 -75.995 ;
        RECT -59.325 -77.685 -58.995 -77.355 ;
        RECT -59.325 -79.045 -58.995 -78.715 ;
        RECT -59.325 -80.405 -58.995 -80.075 ;
        RECT -59.325 -81.765 -58.995 -81.435 ;
        RECT -59.325 -83.125 -58.995 -82.795 ;
        RECT -59.325 -84.485 -58.995 -84.155 ;
        RECT -59.325 -85.845 -58.995 -85.515 ;
        RECT -59.325 -87.205 -58.995 -86.875 ;
        RECT -59.325 -88.565 -58.995 -88.235 ;
        RECT -59.325 -89.925 -58.995 -89.595 ;
        RECT -59.325 -91.285 -58.995 -90.955 ;
        RECT -59.325 -92.645 -58.995 -92.315 ;
        RECT -59.325 -94.005 -58.995 -93.675 ;
        RECT -59.325 -95.365 -58.995 -95.035 ;
        RECT -59.325 -96.725 -58.995 -96.395 ;
        RECT -59.325 -98.085 -58.995 -97.755 ;
        RECT -59.325 -99.445 -58.995 -99.115 ;
        RECT -59.325 -100.805 -58.995 -100.475 ;
        RECT -59.325 -102.165 -58.995 -101.835 ;
        RECT -59.325 -103.525 -58.995 -103.195 ;
        RECT -59.325 -104.885 -58.995 -104.555 ;
        RECT -59.325 -106.245 -58.995 -105.915 ;
        RECT -59.325 -107.605 -58.995 -107.275 ;
        RECT -59.325 -108.965 -58.995 -108.635 ;
        RECT -59.325 -110.325 -58.995 -109.995 ;
        RECT -59.325 -111.685 -58.995 -111.355 ;
        RECT -59.325 -113.045 -58.995 -112.715 ;
        RECT -59.325 -114.405 -58.995 -114.075 ;
        RECT -59.325 -115.765 -58.995 -115.435 ;
        RECT -59.325 -117.125 -58.995 -116.795 ;
        RECT -59.325 -118.485 -58.995 -118.155 ;
        RECT -59.325 -119.845 -58.995 -119.515 ;
        RECT -59.325 -121.205 -58.995 -120.875 ;
        RECT -59.325 -122.565 -58.995 -122.235 ;
        RECT -59.325 -123.925 -58.995 -123.595 ;
        RECT -59.325 -125.285 -58.995 -124.955 ;
        RECT -59.325 -126.645 -58.995 -126.315 ;
        RECT -59.325 -128.005 -58.995 -127.675 ;
        RECT -59.325 -129.365 -58.995 -129.035 ;
        RECT -59.325 -130.725 -58.995 -130.395 ;
        RECT -59.325 -132.085 -58.995 -131.755 ;
        RECT -59.325 -134.805 -58.995 -134.475 ;
        RECT -59.325 -136.165 -58.995 -135.835 ;
        RECT -59.325 -137.525 -58.995 -137.195 ;
        RECT -59.325 -138.885 -58.995 -138.555 ;
        RECT -59.325 -140.245 -58.995 -139.915 ;
        RECT -59.325 -141.605 -58.995 -141.275 ;
        RECT -59.325 -142.965 -58.995 -142.635 ;
        RECT -59.325 -144.325 -58.995 -143.995 ;
        RECT -59.325 -145.685 -58.995 -145.355 ;
        RECT -59.325 -147.045 -58.995 -146.715 ;
        RECT -59.325 -148.405 -58.995 -148.075 ;
        RECT -59.325 -149.765 -58.995 -149.435 ;
        RECT -59.325 -151.125 -58.995 -150.795 ;
        RECT -59.325 -152.485 -58.995 -152.155 ;
        RECT -59.325 -153.845 -58.995 -153.515 ;
        RECT -59.325 -155.205 -58.995 -154.875 ;
        RECT -59.325 -156.565 -58.995 -156.235 ;
        RECT -59.325 -157.925 -58.995 -157.595 ;
        RECT -59.325 -159.285 -58.995 -158.955 ;
        RECT -59.325 -160.645 -58.995 -160.315 ;
        RECT -59.325 -162.005 -58.995 -161.675 ;
        RECT -59.325 -163.365 -58.995 -163.035 ;
        RECT -59.325 -164.725 -58.995 -164.395 ;
        RECT -59.325 -166.085 -58.995 -165.755 ;
        RECT -59.325 -167.445 -58.995 -167.115 ;
        RECT -59.325 -168.805 -58.995 -168.475 ;
        RECT -59.325 -170.165 -58.995 -169.835 ;
        RECT -59.325 -171.525 -58.995 -171.195 ;
        RECT -59.325 -172.885 -58.995 -172.555 ;
        RECT -59.325 -174.245 -58.995 -173.915 ;
        RECT -59.325 -175.605 -58.995 -175.275 ;
        RECT -59.325 -176.965 -58.995 -176.635 ;
        RECT -59.325 -178.325 -58.995 -177.995 ;
        RECT -59.325 -179.685 -58.995 -179.355 ;
        RECT -59.325 -181.045 -58.995 -180.715 ;
        RECT -59.325 -182.405 -58.995 -182.075 ;
        RECT -59.325 -183.765 -58.995 -183.435 ;
        RECT -59.325 -185.125 -58.995 -184.795 ;
        RECT -59.325 -186.485 -58.995 -186.155 ;
        RECT -59.325 -187.845 -58.995 -187.515 ;
        RECT -59.325 -189.205 -58.995 -188.875 ;
        RECT -59.325 -190.565 -58.995 -190.235 ;
        RECT -59.325 -191.925 -58.995 -191.595 ;
        RECT -59.325 -193.285 -58.995 -192.955 ;
        RECT -59.325 -194.645 -58.995 -194.315 ;
        RECT -59.325 -196.005 -58.995 -195.675 ;
        RECT -59.325 -197.365 -58.995 -197.035 ;
        RECT -59.325 -198.725 -58.995 -198.395 ;
        RECT -59.325 -200.085 -58.995 -199.755 ;
        RECT -59.325 -201.445 -58.995 -201.115 ;
        RECT -59.325 -202.805 -58.995 -202.475 ;
        RECT -59.325 -204.165 -58.995 -203.835 ;
        RECT -59.325 -205.525 -58.995 -205.195 ;
        RECT -59.325 -208.245 -58.995 -207.915 ;
        RECT -59.325 -212.325 -58.995 -211.995 ;
        RECT -59.325 -213.625 -58.995 -213.295 ;
        RECT -59.325 -215.045 -58.995 -214.715 ;
        RECT -59.325 -216.405 -58.995 -216.075 ;
        RECT -59.325 -217.765 -58.995 -217.435 ;
        RECT -59.325 -219.125 -58.995 -218.795 ;
        RECT -59.325 -221.37 -58.995 -220.24 ;
        RECT -59.32 -221.485 -59 131.045 ;
        RECT -59.325 129.8 -58.995 130.93 ;
        RECT -59.325 127.675 -58.995 128.005 ;
        RECT -59.325 126.315 -58.995 126.645 ;
        RECT -59.325 124.955 -58.995 125.285 ;
        RECT -59.325 123.595 -58.995 123.925 ;
        RECT -59.325 122.235 -58.995 122.565 ;
        RECT -59.325 120.875 -58.995 121.205 ;
        RECT -59.325 119.515 -58.995 119.845 ;
        RECT -59.325 118.155 -58.995 118.485 ;
        RECT -59.325 116.795 -58.995 117.125 ;
        RECT -59.325 115.435 -58.995 115.765 ;
        RECT -59.325 114.075 -58.995 114.405 ;
        RECT -59.325 112.715 -58.995 113.045 ;
        RECT -59.325 111.355 -58.995 111.685 ;
        RECT -59.325 109.995 -58.995 110.325 ;
        RECT -59.325 108.635 -58.995 108.965 ;
        RECT -59.325 107.275 -58.995 107.605 ;
        RECT -59.325 105.915 -58.995 106.245 ;
        RECT -59.325 104.555 -58.995 104.885 ;
        RECT -59.325 103.195 -58.995 103.525 ;
        RECT -59.325 101.835 -58.995 102.165 ;
        RECT -59.325 100.475 -58.995 100.805 ;
        RECT -59.325 99.115 -58.995 99.445 ;
        RECT -59.325 97.755 -58.995 98.085 ;
        RECT -59.325 96.395 -58.995 96.725 ;
        RECT -59.325 95.035 -58.995 95.365 ;
        RECT -59.325 93.675 -58.995 94.005 ;
        RECT -59.325 92.315 -58.995 92.645 ;
        RECT -59.325 90.955 -58.995 91.285 ;
        RECT -59.325 89.595 -58.995 89.925 ;
        RECT -59.325 88.235 -58.995 88.565 ;
        RECT -59.325 86.875 -58.995 87.205 ;
        RECT -59.325 85.515 -58.995 85.845 ;
        RECT -59.325 84.155 -58.995 84.485 ;
        RECT -59.325 82.795 -58.995 83.125 ;
        RECT -59.325 81.435 -58.995 81.765 ;
        RECT -59.325 80.075 -58.995 80.405 ;
        RECT -59.325 78.715 -58.995 79.045 ;
        RECT -59.325 77.355 -58.995 77.685 ;
        RECT -59.325 75.995 -58.995 76.325 ;
        RECT -59.325 74.635 -58.995 74.965 ;
        RECT -59.325 73.275 -58.995 73.605 ;
        RECT -59.325 71.915 -58.995 72.245 ;
        RECT -59.325 70.555 -58.995 70.885 ;
        RECT -59.325 69.195 -58.995 69.525 ;
        RECT -59.325 67.835 -58.995 68.165 ;
        RECT -59.325 66.475 -58.995 66.805 ;
        RECT -59.325 65.115 -58.995 65.445 ;
        RECT -59.325 63.755 -58.995 64.085 ;
        RECT -59.325 62.395 -58.995 62.725 ;
        RECT -59.325 61.035 -58.995 61.365 ;
        RECT -59.325 59.675 -58.995 60.005 ;
        RECT -59.325 58.315 -58.995 58.645 ;
        RECT -59.325 56.955 -58.995 57.285 ;
        RECT -59.325 55.595 -58.995 55.925 ;
        RECT -59.325 54.235 -58.995 54.565 ;
        RECT -59.325 52.875 -58.995 53.205 ;
        RECT -59.325 51.515 -58.995 51.845 ;
        RECT -59.325 50.155 -58.995 50.485 ;
        RECT -59.325 48.795 -58.995 49.125 ;
        RECT -59.325 47.435 -58.995 47.765 ;
        RECT -59.325 46.075 -58.995 46.405 ;
        RECT -59.325 44.715 -58.995 45.045 ;
        RECT -59.325 43.355 -58.995 43.685 ;
        RECT -59.325 41.995 -58.995 42.325 ;
        RECT -59.325 40.635 -58.995 40.965 ;
        RECT -59.325 39.275 -58.995 39.605 ;
        RECT -59.325 37.915 -58.995 38.245 ;
        RECT -59.325 36.555 -58.995 36.885 ;
        RECT -59.325 35.195 -58.995 35.525 ;
        RECT -59.325 33.835 -58.995 34.165 ;
        RECT -59.325 32.475 -58.995 32.805 ;
        RECT -59.325 31.115 -58.995 31.445 ;
        RECT -59.325 29.755 -58.995 30.085 ;
        RECT -59.325 28.395 -58.995 28.725 ;
        RECT -59.325 27.035 -58.995 27.365 ;
        RECT -59.325 25.675 -58.995 26.005 ;
        RECT -59.325 24.315 -58.995 24.645 ;
        RECT -59.325 22.955 -58.995 23.285 ;
        RECT -59.325 21.595 -58.995 21.925 ;
        RECT -59.325 20.235 -58.995 20.565 ;
        RECT -59.325 18.875 -58.995 19.205 ;
        RECT -59.325 17.515 -58.995 17.845 ;
        RECT -59.325 16.155 -58.995 16.485 ;
        RECT -59.325 14.795 -58.995 15.125 ;
        RECT -59.325 13.435 -58.995 13.765 ;
        RECT -59.325 12.075 -58.995 12.405 ;
        RECT -59.325 10.715 -58.995 11.045 ;
        RECT -59.325 9.355 -58.995 9.685 ;
        RECT -59.325 7.995 -58.995 8.325 ;
        RECT -59.325 6.635 -58.995 6.965 ;
        RECT -59.325 5.275 -58.995 5.605 ;
        RECT -59.325 3.915 -58.995 4.245 ;
        RECT -59.325 2.555 -58.995 2.885 ;
        RECT -59.325 1.195 -58.995 1.525 ;
        RECT -59.325 -0.165 -58.995 0.165 ;
        RECT -59.325 -1.525 -58.995 -1.195 ;
        RECT -59.325 -2.885 -58.995 -2.555 ;
        RECT -59.325 -4.245 -58.995 -3.915 ;
        RECT -59.325 -5.605 -58.995 -5.275 ;
        RECT -59.325 -6.965 -58.995 -6.635 ;
        RECT -59.325 -8.325 -58.995 -7.995 ;
        RECT -59.325 -9.685 -58.995 -9.355 ;
        RECT -59.325 -11.045 -58.995 -10.715 ;
        RECT -59.325 -12.405 -58.995 -12.075 ;
        RECT -59.325 -13.765 -58.995 -13.435 ;
        RECT -59.325 -15.125 -58.995 -14.795 ;
        RECT -59.325 -16.485 -58.995 -16.155 ;
        RECT -59.325 -17.845 -58.995 -17.515 ;
        RECT -59.325 -19.205 -58.995 -18.875 ;
        RECT -59.325 -20.565 -58.995 -20.235 ;
        RECT -59.325 -21.925 -58.995 -21.595 ;
        RECT -59.325 -23.285 -58.995 -22.955 ;
        RECT -59.325 -24.645 -58.995 -24.315 ;
        RECT -59.325 -26.005 -58.995 -25.675 ;
        RECT -59.325 -27.365 -58.995 -27.035 ;
        RECT -59.325 -28.725 -58.995 -28.395 ;
        RECT -59.325 -30.085 -58.995 -29.755 ;
        RECT -59.325 -31.445 -58.995 -31.115 ;
        RECT -59.325 -32.805 -58.995 -32.475 ;
        RECT -59.325 -34.165 -58.995 -33.835 ;
        RECT -59.325 -35.525 -58.995 -35.195 ;
        RECT -59.325 -36.885 -58.995 -36.555 ;
        RECT -59.325 -38.245 -58.995 -37.915 ;
        RECT -59.325 -39.605 -58.995 -39.275 ;
        RECT -59.325 -40.965 -58.995 -40.635 ;
        RECT -59.325 -42.325 -58.995 -41.995 ;
        RECT -59.325 -43.685 -58.995 -43.355 ;
        RECT -59.325 -45.045 -58.995 -44.715 ;
        RECT -59.325 -46.405 -58.995 -46.075 ;
        RECT -59.325 -47.765 -58.995 -47.435 ;
        RECT -59.325 -49.125 -58.995 -48.795 ;
        RECT -59.325 -50.485 -58.995 -50.155 ;
        RECT -59.325 -51.845 -58.995 -51.515 ;
        RECT -59.325 -53.205 -58.995 -52.875 ;
        RECT -59.325 -54.565 -58.995 -54.235 ;
        RECT -59.325 -55.925 -58.995 -55.595 ;
        RECT -59.325 -57.285 -58.995 -56.955 ;
        RECT -59.325 -58.645 -58.995 -58.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -68.845 129.8 -68.515 130.93 ;
        RECT -68.845 127.675 -68.515 128.005 ;
        RECT -68.845 126.315 -68.515 126.645 ;
        RECT -68.845 124.955 -68.515 125.285 ;
        RECT -68.845 123.595 -68.515 123.925 ;
        RECT -68.845 122.235 -68.515 122.565 ;
        RECT -68.845 120.875 -68.515 121.205 ;
        RECT -68.845 119.515 -68.515 119.845 ;
        RECT -68.845 118.155 -68.515 118.485 ;
        RECT -68.845 116.795 -68.515 117.125 ;
        RECT -68.845 115.435 -68.515 115.765 ;
        RECT -68.845 114.075 -68.515 114.405 ;
        RECT -68.845 112.715 -68.515 113.045 ;
        RECT -68.845 111.355 -68.515 111.685 ;
        RECT -68.845 109.995 -68.515 110.325 ;
        RECT -68.845 108.635 -68.515 108.965 ;
        RECT -68.845 107.275 -68.515 107.605 ;
        RECT -68.845 105.915 -68.515 106.245 ;
        RECT -68.845 104.555 -68.515 104.885 ;
        RECT -68.845 103.195 -68.515 103.525 ;
        RECT -68.845 101.835 -68.515 102.165 ;
        RECT -68.845 100.475 -68.515 100.805 ;
        RECT -68.845 99.115 -68.515 99.445 ;
        RECT -68.845 97.755 -68.515 98.085 ;
        RECT -68.845 96.395 -68.515 96.725 ;
        RECT -68.845 95.035 -68.515 95.365 ;
        RECT -68.845 93.675 -68.515 94.005 ;
        RECT -68.845 92.315 -68.515 92.645 ;
        RECT -68.845 90.955 -68.515 91.285 ;
        RECT -68.845 89.595 -68.515 89.925 ;
        RECT -68.845 88.235 -68.515 88.565 ;
        RECT -68.845 86.875 -68.515 87.205 ;
        RECT -68.845 85.515 -68.515 85.845 ;
        RECT -68.845 84.155 -68.515 84.485 ;
        RECT -68.845 82.795 -68.515 83.125 ;
        RECT -68.845 81.435 -68.515 81.765 ;
        RECT -68.845 80.075 -68.515 80.405 ;
        RECT -68.845 78.715 -68.515 79.045 ;
        RECT -68.845 77.355 -68.515 77.685 ;
        RECT -68.845 75.995 -68.515 76.325 ;
        RECT -68.845 74.635 -68.515 74.965 ;
        RECT -68.845 73.275 -68.515 73.605 ;
        RECT -68.845 71.915 -68.515 72.245 ;
        RECT -68.845 70.555 -68.515 70.885 ;
        RECT -68.845 69.195 -68.515 69.525 ;
        RECT -68.845 67.835 -68.515 68.165 ;
        RECT -68.845 66.475 -68.515 66.805 ;
        RECT -68.845 65.115 -68.515 65.445 ;
        RECT -68.845 63.755 -68.515 64.085 ;
        RECT -68.845 62.395 -68.515 62.725 ;
        RECT -68.845 61.035 -68.515 61.365 ;
        RECT -68.845 59.675 -68.515 60.005 ;
        RECT -68.845 58.315 -68.515 58.645 ;
        RECT -68.845 56.955 -68.515 57.285 ;
        RECT -68.845 55.595 -68.515 55.925 ;
        RECT -68.845 54.235 -68.515 54.565 ;
        RECT -68.845 52.875 -68.515 53.205 ;
        RECT -68.845 51.515 -68.515 51.845 ;
        RECT -68.845 50.155 -68.515 50.485 ;
        RECT -68.845 48.795 -68.515 49.125 ;
        RECT -68.845 47.435 -68.515 47.765 ;
        RECT -68.845 46.075 -68.515 46.405 ;
        RECT -68.845 44.715 -68.515 45.045 ;
        RECT -68.845 43.355 -68.515 43.685 ;
        RECT -68.845 41.995 -68.515 42.325 ;
        RECT -68.845 40.635 -68.515 40.965 ;
        RECT -68.845 39.275 -68.515 39.605 ;
        RECT -68.845 37.915 -68.515 38.245 ;
        RECT -68.845 36.555 -68.515 36.885 ;
        RECT -68.845 35.195 -68.515 35.525 ;
        RECT -68.845 33.835 -68.515 34.165 ;
        RECT -68.845 32.475 -68.515 32.805 ;
        RECT -68.845 31.115 -68.515 31.445 ;
        RECT -68.845 29.755 -68.515 30.085 ;
        RECT -68.845 28.395 -68.515 28.725 ;
        RECT -68.845 27.035 -68.515 27.365 ;
        RECT -68.845 25.675 -68.515 26.005 ;
        RECT -68.845 24.315 -68.515 24.645 ;
        RECT -68.845 22.955 -68.515 23.285 ;
        RECT -68.845 21.595 -68.515 21.925 ;
        RECT -68.845 20.235 -68.515 20.565 ;
        RECT -68.845 18.875 -68.515 19.205 ;
        RECT -68.845 17.515 -68.515 17.845 ;
        RECT -68.845 16.155 -68.515 16.485 ;
        RECT -68.845 14.795 -68.515 15.125 ;
        RECT -68.845 13.435 -68.515 13.765 ;
        RECT -68.845 12.075 -68.515 12.405 ;
        RECT -68.845 10.715 -68.515 11.045 ;
        RECT -68.845 9.355 -68.515 9.685 ;
        RECT -68.845 7.995 -68.515 8.325 ;
        RECT -68.845 6.635 -68.515 6.965 ;
        RECT -68.845 5.275 -68.515 5.605 ;
        RECT -68.845 3.915 -68.515 4.245 ;
        RECT -68.845 2.555 -68.515 2.885 ;
        RECT -68.845 1.195 -68.515 1.525 ;
        RECT -68.845 -0.165 -68.515 0.165 ;
        RECT -68.845 -1.525 -68.515 -1.195 ;
        RECT -68.845 -2.885 -68.515 -2.555 ;
        RECT -68.845 -4.245 -68.515 -3.915 ;
        RECT -68.845 -5.605 -68.515 -5.275 ;
        RECT -68.845 -6.965 -68.515 -6.635 ;
        RECT -68.845 -8.325 -68.515 -7.995 ;
        RECT -68.845 -9.685 -68.515 -9.355 ;
        RECT -68.845 -11.045 -68.515 -10.715 ;
        RECT -68.845 -12.405 -68.515 -12.075 ;
        RECT -68.845 -13.765 -68.515 -13.435 ;
        RECT -68.845 -15.125 -68.515 -14.795 ;
        RECT -68.845 -16.485 -68.515 -16.155 ;
        RECT -68.845 -17.845 -68.515 -17.515 ;
        RECT -68.845 -19.205 -68.515 -18.875 ;
        RECT -68.845 -20.565 -68.515 -20.235 ;
        RECT -68.845 -21.925 -68.515 -21.595 ;
        RECT -68.845 -23.285 -68.515 -22.955 ;
        RECT -68.845 -24.645 -68.515 -24.315 ;
        RECT -68.845 -26.005 -68.515 -25.675 ;
        RECT -68.845 -27.365 -68.515 -27.035 ;
        RECT -68.845 -28.725 -68.515 -28.395 ;
        RECT -68.845 -30.085 -68.515 -29.755 ;
        RECT -68.845 -31.445 -68.515 -31.115 ;
        RECT -68.845 -32.805 -68.515 -32.475 ;
        RECT -68.845 -34.165 -68.515 -33.835 ;
        RECT -68.845 -35.525 -68.515 -35.195 ;
        RECT -68.845 -36.885 -68.515 -36.555 ;
        RECT -68.845 -38.245 -68.515 -37.915 ;
        RECT -68.845 -39.605 -68.515 -39.275 ;
        RECT -68.845 -40.965 -68.515 -40.635 ;
        RECT -68.845 -42.325 -68.515 -41.995 ;
        RECT -68.845 -43.685 -68.515 -43.355 ;
        RECT -68.845 -45.045 -68.515 -44.715 ;
        RECT -68.845 -46.405 -68.515 -46.075 ;
        RECT -68.845 -47.765 -68.515 -47.435 ;
        RECT -68.845 -49.125 -68.515 -48.795 ;
        RECT -68.845 -50.485 -68.515 -50.155 ;
        RECT -68.845 -51.845 -68.515 -51.515 ;
        RECT -68.845 -53.205 -68.515 -52.875 ;
        RECT -68.845 -54.565 -68.515 -54.235 ;
        RECT -68.845 -55.925 -68.515 -55.595 ;
        RECT -68.845 -57.285 -68.515 -56.955 ;
        RECT -68.845 -58.645 -68.515 -58.315 ;
        RECT -68.845 -60.005 -68.515 -59.675 ;
        RECT -68.845 -61.365 -68.515 -61.035 ;
        RECT -68.845 -62.725 -68.515 -62.395 ;
        RECT -68.845 -64.085 -68.515 -63.755 ;
        RECT -68.845 -65.445 -68.515 -65.115 ;
        RECT -68.845 -66.805 -68.515 -66.475 ;
        RECT -68.845 -68.165 -68.515 -67.835 ;
        RECT -68.845 -69.525 -68.515 -69.195 ;
        RECT -68.845 -70.885 -68.515 -70.555 ;
        RECT -68.845 -72.245 -68.515 -71.915 ;
        RECT -68.845 -73.605 -68.515 -73.275 ;
        RECT -68.845 -74.965 -68.515 -74.635 ;
        RECT -68.845 -76.325 -68.515 -75.995 ;
        RECT -68.845 -77.685 -68.515 -77.355 ;
        RECT -68.845 -79.045 -68.515 -78.715 ;
        RECT -68.845 -80.405 -68.515 -80.075 ;
        RECT -68.845 -81.765 -68.515 -81.435 ;
        RECT -68.845 -83.125 -68.515 -82.795 ;
        RECT -68.845 -84.485 -68.515 -84.155 ;
        RECT -68.845 -85.845 -68.515 -85.515 ;
        RECT -68.845 -87.205 -68.515 -86.875 ;
        RECT -68.845 -88.565 -68.515 -88.235 ;
        RECT -68.845 -89.925 -68.515 -89.595 ;
        RECT -68.845 -91.285 -68.515 -90.955 ;
        RECT -68.845 -92.645 -68.515 -92.315 ;
        RECT -68.845 -94.005 -68.515 -93.675 ;
        RECT -68.845 -95.365 -68.515 -95.035 ;
        RECT -68.845 -96.725 -68.515 -96.395 ;
        RECT -68.845 -98.085 -68.515 -97.755 ;
        RECT -68.845 -99.445 -68.515 -99.115 ;
        RECT -68.845 -100.805 -68.515 -100.475 ;
        RECT -68.845 -102.165 -68.515 -101.835 ;
        RECT -68.845 -103.525 -68.515 -103.195 ;
        RECT -68.845 -104.885 -68.515 -104.555 ;
        RECT -68.845 -106.245 -68.515 -105.915 ;
        RECT -68.845 -107.605 -68.515 -107.275 ;
        RECT -68.845 -108.965 -68.515 -108.635 ;
        RECT -68.845 -110.325 -68.515 -109.995 ;
        RECT -68.845 -111.685 -68.515 -111.355 ;
        RECT -68.845 -113.045 -68.515 -112.715 ;
        RECT -68.845 -114.405 -68.515 -114.075 ;
        RECT -68.845 -115.765 -68.515 -115.435 ;
        RECT -68.845 -117.125 -68.515 -116.795 ;
        RECT -68.845 -118.485 -68.515 -118.155 ;
        RECT -68.845 -119.845 -68.515 -119.515 ;
        RECT -68.845 -121.205 -68.515 -120.875 ;
        RECT -68.845 -122.565 -68.515 -122.235 ;
        RECT -68.845 -123.925 -68.515 -123.595 ;
        RECT -68.845 -125.285 -68.515 -124.955 ;
        RECT -68.845 -126.645 -68.515 -126.315 ;
        RECT -68.845 -128.005 -68.515 -127.675 ;
        RECT -68.845 -129.365 -68.515 -129.035 ;
        RECT -68.845 -130.725 -68.515 -130.395 ;
        RECT -68.845 -132.085 -68.515 -131.755 ;
        RECT -68.845 -133.445 -68.515 -133.115 ;
        RECT -68.845 -134.805 -68.515 -134.475 ;
        RECT -68.845 -136.165 -68.515 -135.835 ;
        RECT -68.845 -137.525 -68.515 -137.195 ;
        RECT -68.845 -138.885 -68.515 -138.555 ;
        RECT -68.845 -140.245 -68.515 -139.915 ;
        RECT -68.845 -141.605 -68.515 -141.275 ;
        RECT -68.845 -142.965 -68.515 -142.635 ;
        RECT -68.845 -144.325 -68.515 -143.995 ;
        RECT -68.845 -145.685 -68.515 -145.355 ;
        RECT -68.845 -147.045 -68.515 -146.715 ;
        RECT -68.845 -148.405 -68.515 -148.075 ;
        RECT -68.845 -149.765 -68.515 -149.435 ;
        RECT -68.845 -151.125 -68.515 -150.795 ;
        RECT -68.845 -152.485 -68.515 -152.155 ;
        RECT -68.845 -153.845 -68.515 -153.515 ;
        RECT -68.845 -155.205 -68.515 -154.875 ;
        RECT -68.845 -156.565 -68.515 -156.235 ;
        RECT -68.845 -157.925 -68.515 -157.595 ;
        RECT -68.845 -159.285 -68.515 -158.955 ;
        RECT -68.845 -160.645 -68.515 -160.315 ;
        RECT -68.845 -162.005 -68.515 -161.675 ;
        RECT -68.845 -163.365 -68.515 -163.035 ;
        RECT -68.845 -164.725 -68.515 -164.395 ;
        RECT -68.845 -166.085 -68.515 -165.755 ;
        RECT -68.845 -167.445 -68.515 -167.115 ;
        RECT -68.845 -168.805 -68.515 -168.475 ;
        RECT -68.845 -170.165 -68.515 -169.835 ;
        RECT -68.845 -171.525 -68.515 -171.195 ;
        RECT -68.845 -172.885 -68.515 -172.555 ;
        RECT -68.845 -174.245 -68.515 -173.915 ;
        RECT -68.845 -175.605 -68.515 -175.275 ;
        RECT -68.845 -176.965 -68.515 -176.635 ;
        RECT -68.845 -178.325 -68.515 -177.995 ;
        RECT -68.845 -179.685 -68.515 -179.355 ;
        RECT -68.845 -181.045 -68.515 -180.715 ;
        RECT -68.845 -182.405 -68.515 -182.075 ;
        RECT -68.845 -183.765 -68.515 -183.435 ;
        RECT -68.845 -185.125 -68.515 -184.795 ;
        RECT -68.845 -186.485 -68.515 -186.155 ;
        RECT -68.845 -187.845 -68.515 -187.515 ;
        RECT -68.845 -189.205 -68.515 -188.875 ;
        RECT -68.845 -190.565 -68.515 -190.235 ;
        RECT -68.845 -191.925 -68.515 -191.595 ;
        RECT -68.845 -193.285 -68.515 -192.955 ;
        RECT -68.845 -194.645 -68.515 -194.315 ;
        RECT -68.845 -196.005 -68.515 -195.675 ;
        RECT -68.845 -197.365 -68.515 -197.035 ;
        RECT -68.845 -198.725 -68.515 -198.395 ;
        RECT -68.845 -200.085 -68.515 -199.755 ;
        RECT -68.845 -201.445 -68.515 -201.115 ;
        RECT -68.845 -202.805 -68.515 -202.475 ;
        RECT -68.845 -204.165 -68.515 -203.835 ;
        RECT -68.845 -205.525 -68.515 -205.195 ;
        RECT -68.845 -206.885 -68.515 -206.555 ;
        RECT -68.845 -208.245 -68.515 -207.915 ;
        RECT -68.845 -209.605 -68.515 -209.275 ;
        RECT -68.845 -210.965 -68.515 -210.635 ;
        RECT -68.845 -212.325 -68.515 -211.995 ;
        RECT -68.845 -213.685 -68.515 -213.355 ;
        RECT -68.845 -215.045 -68.515 -214.715 ;
        RECT -68.845 -216.405 -68.515 -216.075 ;
        RECT -68.845 -217.765 -68.515 -217.435 ;
        RECT -68.845 -219.125 -68.515 -218.795 ;
        RECT -68.845 -221.37 -68.515 -220.24 ;
        RECT -68.84 -221.485 -68.52 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -67.485 129.8 -67.155 130.93 ;
        RECT -67.485 127.675 -67.155 128.005 ;
        RECT -67.485 126.315 -67.155 126.645 ;
        RECT -67.485 124.955 -67.155 125.285 ;
        RECT -67.485 123.595 -67.155 123.925 ;
        RECT -67.485 122.235 -67.155 122.565 ;
        RECT -67.485 120.875 -67.155 121.205 ;
        RECT -67.485 119.515 -67.155 119.845 ;
        RECT -67.485 118.155 -67.155 118.485 ;
        RECT -67.485 116.795 -67.155 117.125 ;
        RECT -67.485 115.435 -67.155 115.765 ;
        RECT -67.485 114.075 -67.155 114.405 ;
        RECT -67.485 112.715 -67.155 113.045 ;
        RECT -67.485 111.355 -67.155 111.685 ;
        RECT -67.485 109.995 -67.155 110.325 ;
        RECT -67.485 108.635 -67.155 108.965 ;
        RECT -67.485 107.275 -67.155 107.605 ;
        RECT -67.485 105.915 -67.155 106.245 ;
        RECT -67.485 104.555 -67.155 104.885 ;
        RECT -67.485 103.195 -67.155 103.525 ;
        RECT -67.485 101.835 -67.155 102.165 ;
        RECT -67.485 100.475 -67.155 100.805 ;
        RECT -67.485 99.115 -67.155 99.445 ;
        RECT -67.485 97.755 -67.155 98.085 ;
        RECT -67.485 96.395 -67.155 96.725 ;
        RECT -67.485 95.035 -67.155 95.365 ;
        RECT -67.485 93.675 -67.155 94.005 ;
        RECT -67.485 92.315 -67.155 92.645 ;
        RECT -67.485 90.955 -67.155 91.285 ;
        RECT -67.485 89.595 -67.155 89.925 ;
        RECT -67.485 88.235 -67.155 88.565 ;
        RECT -67.485 86.875 -67.155 87.205 ;
        RECT -67.485 85.515 -67.155 85.845 ;
        RECT -67.485 84.155 -67.155 84.485 ;
        RECT -67.485 82.795 -67.155 83.125 ;
        RECT -67.485 81.435 -67.155 81.765 ;
        RECT -67.485 80.075 -67.155 80.405 ;
        RECT -67.485 78.715 -67.155 79.045 ;
        RECT -67.485 77.355 -67.155 77.685 ;
        RECT -67.485 75.995 -67.155 76.325 ;
        RECT -67.485 74.635 -67.155 74.965 ;
        RECT -67.485 73.275 -67.155 73.605 ;
        RECT -67.485 71.915 -67.155 72.245 ;
        RECT -67.485 70.555 -67.155 70.885 ;
        RECT -67.485 69.195 -67.155 69.525 ;
        RECT -67.485 67.835 -67.155 68.165 ;
        RECT -67.485 66.475 -67.155 66.805 ;
        RECT -67.485 65.115 -67.155 65.445 ;
        RECT -67.485 63.755 -67.155 64.085 ;
        RECT -67.485 62.395 -67.155 62.725 ;
        RECT -67.485 61.035 -67.155 61.365 ;
        RECT -67.485 59.675 -67.155 60.005 ;
        RECT -67.485 58.315 -67.155 58.645 ;
        RECT -67.485 56.955 -67.155 57.285 ;
        RECT -67.485 55.595 -67.155 55.925 ;
        RECT -67.485 54.235 -67.155 54.565 ;
        RECT -67.485 52.875 -67.155 53.205 ;
        RECT -67.485 51.515 -67.155 51.845 ;
        RECT -67.485 50.155 -67.155 50.485 ;
        RECT -67.485 48.795 -67.155 49.125 ;
        RECT -67.485 47.435 -67.155 47.765 ;
        RECT -67.485 46.075 -67.155 46.405 ;
        RECT -67.485 44.715 -67.155 45.045 ;
        RECT -67.485 43.355 -67.155 43.685 ;
        RECT -67.485 41.995 -67.155 42.325 ;
        RECT -67.485 40.635 -67.155 40.965 ;
        RECT -67.485 39.275 -67.155 39.605 ;
        RECT -67.485 37.915 -67.155 38.245 ;
        RECT -67.485 36.555 -67.155 36.885 ;
        RECT -67.485 35.195 -67.155 35.525 ;
        RECT -67.485 33.835 -67.155 34.165 ;
        RECT -67.485 32.475 -67.155 32.805 ;
        RECT -67.485 31.115 -67.155 31.445 ;
        RECT -67.485 29.755 -67.155 30.085 ;
        RECT -67.485 28.395 -67.155 28.725 ;
        RECT -67.485 27.035 -67.155 27.365 ;
        RECT -67.485 25.675 -67.155 26.005 ;
        RECT -67.485 24.315 -67.155 24.645 ;
        RECT -67.485 22.955 -67.155 23.285 ;
        RECT -67.485 21.595 -67.155 21.925 ;
        RECT -67.485 20.235 -67.155 20.565 ;
        RECT -67.485 18.875 -67.155 19.205 ;
        RECT -67.485 17.515 -67.155 17.845 ;
        RECT -67.485 16.155 -67.155 16.485 ;
        RECT -67.485 14.795 -67.155 15.125 ;
        RECT -67.485 13.435 -67.155 13.765 ;
        RECT -67.485 12.075 -67.155 12.405 ;
        RECT -67.485 10.715 -67.155 11.045 ;
        RECT -67.485 9.355 -67.155 9.685 ;
        RECT -67.485 7.995 -67.155 8.325 ;
        RECT -67.485 6.635 -67.155 6.965 ;
        RECT -67.485 5.275 -67.155 5.605 ;
        RECT -67.485 3.915 -67.155 4.245 ;
        RECT -67.485 2.555 -67.155 2.885 ;
        RECT -67.485 1.195 -67.155 1.525 ;
        RECT -67.485 -0.165 -67.155 0.165 ;
        RECT -67.485 -1.525 -67.155 -1.195 ;
        RECT -67.485 -2.885 -67.155 -2.555 ;
        RECT -67.485 -4.245 -67.155 -3.915 ;
        RECT -67.485 -5.605 -67.155 -5.275 ;
        RECT -67.485 -6.965 -67.155 -6.635 ;
        RECT -67.485 -8.325 -67.155 -7.995 ;
        RECT -67.485 -9.685 -67.155 -9.355 ;
        RECT -67.485 -11.045 -67.155 -10.715 ;
        RECT -67.485 -12.405 -67.155 -12.075 ;
        RECT -67.485 -13.765 -67.155 -13.435 ;
        RECT -67.485 -15.125 -67.155 -14.795 ;
        RECT -67.485 -16.485 -67.155 -16.155 ;
        RECT -67.485 -17.845 -67.155 -17.515 ;
        RECT -67.485 -19.205 -67.155 -18.875 ;
        RECT -67.485 -20.565 -67.155 -20.235 ;
        RECT -67.485 -21.925 -67.155 -21.595 ;
        RECT -67.485 -23.285 -67.155 -22.955 ;
        RECT -67.485 -24.645 -67.155 -24.315 ;
        RECT -67.485 -26.005 -67.155 -25.675 ;
        RECT -67.485 -27.365 -67.155 -27.035 ;
        RECT -67.485 -28.725 -67.155 -28.395 ;
        RECT -67.485 -30.085 -67.155 -29.755 ;
        RECT -67.485 -31.445 -67.155 -31.115 ;
        RECT -67.485 -32.805 -67.155 -32.475 ;
        RECT -67.485 -34.165 -67.155 -33.835 ;
        RECT -67.485 -35.525 -67.155 -35.195 ;
        RECT -67.485 -36.885 -67.155 -36.555 ;
        RECT -67.485 -38.245 -67.155 -37.915 ;
        RECT -67.485 -39.605 -67.155 -39.275 ;
        RECT -67.485 -40.965 -67.155 -40.635 ;
        RECT -67.485 -42.325 -67.155 -41.995 ;
        RECT -67.485 -43.685 -67.155 -43.355 ;
        RECT -67.485 -45.045 -67.155 -44.715 ;
        RECT -67.485 -46.405 -67.155 -46.075 ;
        RECT -67.485 -47.765 -67.155 -47.435 ;
        RECT -67.485 -49.125 -67.155 -48.795 ;
        RECT -67.485 -50.485 -67.155 -50.155 ;
        RECT -67.485 -51.845 -67.155 -51.515 ;
        RECT -67.485 -53.205 -67.155 -52.875 ;
        RECT -67.485 -54.565 -67.155 -54.235 ;
        RECT -67.485 -55.925 -67.155 -55.595 ;
        RECT -67.485 -57.285 -67.155 -56.955 ;
        RECT -67.485 -58.645 -67.155 -58.315 ;
        RECT -67.485 -60.005 -67.155 -59.675 ;
        RECT -67.485 -61.365 -67.155 -61.035 ;
        RECT -67.485 -62.725 -67.155 -62.395 ;
        RECT -67.485 -64.085 -67.155 -63.755 ;
        RECT -67.485 -65.445 -67.155 -65.115 ;
        RECT -67.485 -66.805 -67.155 -66.475 ;
        RECT -67.485 -68.165 -67.155 -67.835 ;
        RECT -67.485 -69.525 -67.155 -69.195 ;
        RECT -67.485 -70.885 -67.155 -70.555 ;
        RECT -67.485 -72.245 -67.155 -71.915 ;
        RECT -67.485 -73.605 -67.155 -73.275 ;
        RECT -67.485 -74.965 -67.155 -74.635 ;
        RECT -67.485 -76.325 -67.155 -75.995 ;
        RECT -67.485 -77.685 -67.155 -77.355 ;
        RECT -67.485 -79.045 -67.155 -78.715 ;
        RECT -67.485 -80.405 -67.155 -80.075 ;
        RECT -67.485 -81.765 -67.155 -81.435 ;
        RECT -67.485 -83.125 -67.155 -82.795 ;
        RECT -67.485 -84.485 -67.155 -84.155 ;
        RECT -67.485 -85.845 -67.155 -85.515 ;
        RECT -67.485 -87.205 -67.155 -86.875 ;
        RECT -67.485 -88.565 -67.155 -88.235 ;
        RECT -67.485 -89.925 -67.155 -89.595 ;
        RECT -67.485 -91.285 -67.155 -90.955 ;
        RECT -67.485 -92.645 -67.155 -92.315 ;
        RECT -67.485 -94.005 -67.155 -93.675 ;
        RECT -67.485 -95.365 -67.155 -95.035 ;
        RECT -67.485 -96.725 -67.155 -96.395 ;
        RECT -67.485 -98.085 -67.155 -97.755 ;
        RECT -67.485 -99.445 -67.155 -99.115 ;
        RECT -67.485 -100.805 -67.155 -100.475 ;
        RECT -67.485 -102.165 -67.155 -101.835 ;
        RECT -67.485 -103.525 -67.155 -103.195 ;
        RECT -67.485 -104.885 -67.155 -104.555 ;
        RECT -67.485 -106.245 -67.155 -105.915 ;
        RECT -67.485 -107.605 -67.155 -107.275 ;
        RECT -67.485 -108.965 -67.155 -108.635 ;
        RECT -67.485 -110.325 -67.155 -109.995 ;
        RECT -67.485 -111.685 -67.155 -111.355 ;
        RECT -67.485 -113.045 -67.155 -112.715 ;
        RECT -67.485 -114.405 -67.155 -114.075 ;
        RECT -67.485 -115.765 -67.155 -115.435 ;
        RECT -67.485 -117.125 -67.155 -116.795 ;
        RECT -67.485 -118.485 -67.155 -118.155 ;
        RECT -67.485 -119.845 -67.155 -119.515 ;
        RECT -67.485 -121.205 -67.155 -120.875 ;
        RECT -67.485 -122.565 -67.155 -122.235 ;
        RECT -67.485 -123.925 -67.155 -123.595 ;
        RECT -67.485 -125.285 -67.155 -124.955 ;
        RECT -67.485 -126.645 -67.155 -126.315 ;
        RECT -67.485 -128.005 -67.155 -127.675 ;
        RECT -67.485 -129.365 -67.155 -129.035 ;
        RECT -67.485 -130.725 -67.155 -130.395 ;
        RECT -67.485 -132.085 -67.155 -131.755 ;
        RECT -67.485 -133.445 -67.155 -133.115 ;
        RECT -67.485 -134.805 -67.155 -134.475 ;
        RECT -67.485 -136.165 -67.155 -135.835 ;
        RECT -67.485 -137.525 -67.155 -137.195 ;
        RECT -67.485 -138.885 -67.155 -138.555 ;
        RECT -67.485 -140.245 -67.155 -139.915 ;
        RECT -67.485 -141.605 -67.155 -141.275 ;
        RECT -67.485 -142.965 -67.155 -142.635 ;
        RECT -67.485 -144.325 -67.155 -143.995 ;
        RECT -67.485 -145.685 -67.155 -145.355 ;
        RECT -67.485 -147.045 -67.155 -146.715 ;
        RECT -67.485 -148.405 -67.155 -148.075 ;
        RECT -67.485 -149.765 -67.155 -149.435 ;
        RECT -67.485 -151.125 -67.155 -150.795 ;
        RECT -67.485 -152.485 -67.155 -152.155 ;
        RECT -67.485 -153.845 -67.155 -153.515 ;
        RECT -67.485 -155.205 -67.155 -154.875 ;
        RECT -67.485 -156.565 -67.155 -156.235 ;
        RECT -67.485 -157.925 -67.155 -157.595 ;
        RECT -67.485 -159.285 -67.155 -158.955 ;
        RECT -67.485 -160.645 -67.155 -160.315 ;
        RECT -67.485 -162.005 -67.155 -161.675 ;
        RECT -67.485 -163.365 -67.155 -163.035 ;
        RECT -67.485 -164.725 -67.155 -164.395 ;
        RECT -67.485 -166.085 -67.155 -165.755 ;
        RECT -67.485 -167.445 -67.155 -167.115 ;
        RECT -67.485 -168.805 -67.155 -168.475 ;
        RECT -67.485 -170.165 -67.155 -169.835 ;
        RECT -67.485 -171.525 -67.155 -171.195 ;
        RECT -67.485 -172.885 -67.155 -172.555 ;
        RECT -67.485 -174.245 -67.155 -173.915 ;
        RECT -67.485 -175.605 -67.155 -175.275 ;
        RECT -67.485 -176.965 -67.155 -176.635 ;
        RECT -67.485 -178.325 -67.155 -177.995 ;
        RECT -67.485 -179.685 -67.155 -179.355 ;
        RECT -67.485 -181.045 -67.155 -180.715 ;
        RECT -67.485 -182.405 -67.155 -182.075 ;
        RECT -67.485 -183.765 -67.155 -183.435 ;
        RECT -67.485 -185.125 -67.155 -184.795 ;
        RECT -67.485 -186.485 -67.155 -186.155 ;
        RECT -67.485 -187.845 -67.155 -187.515 ;
        RECT -67.485 -189.205 -67.155 -188.875 ;
        RECT -67.485 -190.565 -67.155 -190.235 ;
        RECT -67.485 -191.925 -67.155 -191.595 ;
        RECT -67.485 -193.285 -67.155 -192.955 ;
        RECT -67.485 -194.645 -67.155 -194.315 ;
        RECT -67.485 -196.005 -67.155 -195.675 ;
        RECT -67.485 -197.365 -67.155 -197.035 ;
        RECT -67.485 -198.725 -67.155 -198.395 ;
        RECT -67.485 -200.085 -67.155 -199.755 ;
        RECT -67.485 -201.445 -67.155 -201.115 ;
        RECT -67.485 -202.805 -67.155 -202.475 ;
        RECT -67.485 -204.165 -67.155 -203.835 ;
        RECT -67.485 -205.525 -67.155 -205.195 ;
        RECT -67.485 -206.885 -67.155 -206.555 ;
        RECT -67.485 -208.245 -67.155 -207.915 ;
        RECT -67.485 -209.605 -67.155 -209.275 ;
        RECT -67.485 -210.965 -67.155 -210.635 ;
        RECT -67.485 -212.325 -67.155 -211.995 ;
        RECT -67.485 -213.685 -67.155 -213.355 ;
        RECT -67.485 -215.045 -67.155 -214.715 ;
        RECT -67.485 -216.405 -67.155 -216.075 ;
        RECT -67.485 -217.765 -67.155 -217.435 ;
        RECT -67.485 -219.125 -67.155 -218.795 ;
        RECT -67.485 -221.37 -67.155 -220.24 ;
        RECT -67.48 -221.485 -67.16 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -66.125 129.8 -65.795 130.93 ;
        RECT -66.125 127.675 -65.795 128.005 ;
        RECT -66.125 126.315 -65.795 126.645 ;
        RECT -66.125 124.955 -65.795 125.285 ;
        RECT -66.125 123.595 -65.795 123.925 ;
        RECT -66.125 122.235 -65.795 122.565 ;
        RECT -66.125 120.875 -65.795 121.205 ;
        RECT -66.125 119.515 -65.795 119.845 ;
        RECT -66.125 118.155 -65.795 118.485 ;
        RECT -66.125 116.795 -65.795 117.125 ;
        RECT -66.125 115.435 -65.795 115.765 ;
        RECT -66.125 114.075 -65.795 114.405 ;
        RECT -66.125 112.715 -65.795 113.045 ;
        RECT -66.125 111.355 -65.795 111.685 ;
        RECT -66.125 109.995 -65.795 110.325 ;
        RECT -66.125 108.635 -65.795 108.965 ;
        RECT -66.125 107.275 -65.795 107.605 ;
        RECT -66.125 105.915 -65.795 106.245 ;
        RECT -66.125 104.555 -65.795 104.885 ;
        RECT -66.125 103.195 -65.795 103.525 ;
        RECT -66.125 101.835 -65.795 102.165 ;
        RECT -66.125 100.475 -65.795 100.805 ;
        RECT -66.125 99.115 -65.795 99.445 ;
        RECT -66.125 97.755 -65.795 98.085 ;
        RECT -66.125 96.395 -65.795 96.725 ;
        RECT -66.125 95.035 -65.795 95.365 ;
        RECT -66.125 93.675 -65.795 94.005 ;
        RECT -66.125 92.315 -65.795 92.645 ;
        RECT -66.125 90.955 -65.795 91.285 ;
        RECT -66.125 89.595 -65.795 89.925 ;
        RECT -66.125 88.235 -65.795 88.565 ;
        RECT -66.125 86.875 -65.795 87.205 ;
        RECT -66.125 85.515 -65.795 85.845 ;
        RECT -66.125 84.155 -65.795 84.485 ;
        RECT -66.125 82.795 -65.795 83.125 ;
        RECT -66.125 81.435 -65.795 81.765 ;
        RECT -66.125 80.075 -65.795 80.405 ;
        RECT -66.125 78.715 -65.795 79.045 ;
        RECT -66.125 77.355 -65.795 77.685 ;
        RECT -66.125 75.995 -65.795 76.325 ;
        RECT -66.125 74.635 -65.795 74.965 ;
        RECT -66.125 73.275 -65.795 73.605 ;
        RECT -66.125 71.915 -65.795 72.245 ;
        RECT -66.125 70.555 -65.795 70.885 ;
        RECT -66.125 69.195 -65.795 69.525 ;
        RECT -66.125 67.835 -65.795 68.165 ;
        RECT -66.125 66.475 -65.795 66.805 ;
        RECT -66.125 65.115 -65.795 65.445 ;
        RECT -66.125 63.755 -65.795 64.085 ;
        RECT -66.125 62.395 -65.795 62.725 ;
        RECT -66.125 61.035 -65.795 61.365 ;
        RECT -66.125 59.675 -65.795 60.005 ;
        RECT -66.125 58.315 -65.795 58.645 ;
        RECT -66.125 56.955 -65.795 57.285 ;
        RECT -66.125 55.595 -65.795 55.925 ;
        RECT -66.125 54.235 -65.795 54.565 ;
        RECT -66.125 52.875 -65.795 53.205 ;
        RECT -66.125 51.515 -65.795 51.845 ;
        RECT -66.125 50.155 -65.795 50.485 ;
        RECT -66.125 48.795 -65.795 49.125 ;
        RECT -66.125 47.435 -65.795 47.765 ;
        RECT -66.125 46.075 -65.795 46.405 ;
        RECT -66.125 44.715 -65.795 45.045 ;
        RECT -66.125 43.355 -65.795 43.685 ;
        RECT -66.125 41.995 -65.795 42.325 ;
        RECT -66.125 40.635 -65.795 40.965 ;
        RECT -66.125 39.275 -65.795 39.605 ;
        RECT -66.125 37.915 -65.795 38.245 ;
        RECT -66.125 36.555 -65.795 36.885 ;
        RECT -66.125 35.195 -65.795 35.525 ;
        RECT -66.125 33.835 -65.795 34.165 ;
        RECT -66.125 32.475 -65.795 32.805 ;
        RECT -66.125 31.115 -65.795 31.445 ;
        RECT -66.125 29.755 -65.795 30.085 ;
        RECT -66.125 28.395 -65.795 28.725 ;
        RECT -66.125 27.035 -65.795 27.365 ;
        RECT -66.125 25.675 -65.795 26.005 ;
        RECT -66.125 24.315 -65.795 24.645 ;
        RECT -66.125 22.955 -65.795 23.285 ;
        RECT -66.125 21.595 -65.795 21.925 ;
        RECT -66.125 20.235 -65.795 20.565 ;
        RECT -66.125 18.875 -65.795 19.205 ;
        RECT -66.125 17.515 -65.795 17.845 ;
        RECT -66.125 16.155 -65.795 16.485 ;
        RECT -66.125 14.795 -65.795 15.125 ;
        RECT -66.125 13.435 -65.795 13.765 ;
        RECT -66.125 12.075 -65.795 12.405 ;
        RECT -66.125 10.715 -65.795 11.045 ;
        RECT -66.125 9.355 -65.795 9.685 ;
        RECT -66.125 7.995 -65.795 8.325 ;
        RECT -66.125 6.635 -65.795 6.965 ;
        RECT -66.125 5.275 -65.795 5.605 ;
        RECT -66.125 3.915 -65.795 4.245 ;
        RECT -66.125 2.555 -65.795 2.885 ;
        RECT -66.125 1.195 -65.795 1.525 ;
        RECT -66.125 -0.165 -65.795 0.165 ;
        RECT -66.125 -1.525 -65.795 -1.195 ;
        RECT -66.125 -2.885 -65.795 -2.555 ;
        RECT -66.125 -4.245 -65.795 -3.915 ;
        RECT -66.125 -5.605 -65.795 -5.275 ;
        RECT -66.125 -6.965 -65.795 -6.635 ;
        RECT -66.125 -8.325 -65.795 -7.995 ;
        RECT -66.125 -9.685 -65.795 -9.355 ;
        RECT -66.125 -11.045 -65.795 -10.715 ;
        RECT -66.125 -12.405 -65.795 -12.075 ;
        RECT -66.125 -13.765 -65.795 -13.435 ;
        RECT -66.125 -15.125 -65.795 -14.795 ;
        RECT -66.125 -16.485 -65.795 -16.155 ;
        RECT -66.125 -17.845 -65.795 -17.515 ;
        RECT -66.125 -19.205 -65.795 -18.875 ;
        RECT -66.125 -20.565 -65.795 -20.235 ;
        RECT -66.125 -21.925 -65.795 -21.595 ;
        RECT -66.125 -23.285 -65.795 -22.955 ;
        RECT -66.125 -24.645 -65.795 -24.315 ;
        RECT -66.125 -26.005 -65.795 -25.675 ;
        RECT -66.125 -27.365 -65.795 -27.035 ;
        RECT -66.125 -28.725 -65.795 -28.395 ;
        RECT -66.125 -30.085 -65.795 -29.755 ;
        RECT -66.125 -31.445 -65.795 -31.115 ;
        RECT -66.125 -32.805 -65.795 -32.475 ;
        RECT -66.125 -34.165 -65.795 -33.835 ;
        RECT -66.125 -35.525 -65.795 -35.195 ;
        RECT -66.125 -36.885 -65.795 -36.555 ;
        RECT -66.125 -38.245 -65.795 -37.915 ;
        RECT -66.125 -39.605 -65.795 -39.275 ;
        RECT -66.125 -40.965 -65.795 -40.635 ;
        RECT -66.125 -42.325 -65.795 -41.995 ;
        RECT -66.125 -43.685 -65.795 -43.355 ;
        RECT -66.125 -45.045 -65.795 -44.715 ;
        RECT -66.125 -46.405 -65.795 -46.075 ;
        RECT -66.125 -47.765 -65.795 -47.435 ;
        RECT -66.125 -49.125 -65.795 -48.795 ;
        RECT -66.125 -50.485 -65.795 -50.155 ;
        RECT -66.125 -51.845 -65.795 -51.515 ;
        RECT -66.125 -53.205 -65.795 -52.875 ;
        RECT -66.125 -54.565 -65.795 -54.235 ;
        RECT -66.125 -55.925 -65.795 -55.595 ;
        RECT -66.125 -57.285 -65.795 -56.955 ;
        RECT -66.125 -58.645 -65.795 -58.315 ;
        RECT -66.125 -60.005 -65.795 -59.675 ;
        RECT -66.125 -61.365 -65.795 -61.035 ;
        RECT -66.125 -62.725 -65.795 -62.395 ;
        RECT -66.125 -64.085 -65.795 -63.755 ;
        RECT -66.125 -65.445 -65.795 -65.115 ;
        RECT -66.125 -66.805 -65.795 -66.475 ;
        RECT -66.125 -68.165 -65.795 -67.835 ;
        RECT -66.125 -69.525 -65.795 -69.195 ;
        RECT -66.125 -70.885 -65.795 -70.555 ;
        RECT -66.125 -72.245 -65.795 -71.915 ;
        RECT -66.125 -73.605 -65.795 -73.275 ;
        RECT -66.125 -74.965 -65.795 -74.635 ;
        RECT -66.125 -76.325 -65.795 -75.995 ;
        RECT -66.125 -77.685 -65.795 -77.355 ;
        RECT -66.125 -79.045 -65.795 -78.715 ;
        RECT -66.125 -80.405 -65.795 -80.075 ;
        RECT -66.125 -81.765 -65.795 -81.435 ;
        RECT -66.125 -83.125 -65.795 -82.795 ;
        RECT -66.125 -84.485 -65.795 -84.155 ;
        RECT -66.125 -85.845 -65.795 -85.515 ;
        RECT -66.125 -87.205 -65.795 -86.875 ;
        RECT -66.125 -88.565 -65.795 -88.235 ;
        RECT -66.125 -89.925 -65.795 -89.595 ;
        RECT -66.125 -91.285 -65.795 -90.955 ;
        RECT -66.125 -92.645 -65.795 -92.315 ;
        RECT -66.125 -94.005 -65.795 -93.675 ;
        RECT -66.125 -95.365 -65.795 -95.035 ;
        RECT -66.125 -96.725 -65.795 -96.395 ;
        RECT -66.125 -98.085 -65.795 -97.755 ;
        RECT -66.125 -99.445 -65.795 -99.115 ;
        RECT -66.125 -100.805 -65.795 -100.475 ;
        RECT -66.125 -102.165 -65.795 -101.835 ;
        RECT -66.125 -103.525 -65.795 -103.195 ;
        RECT -66.125 -104.885 -65.795 -104.555 ;
        RECT -66.125 -106.245 -65.795 -105.915 ;
        RECT -66.125 -107.605 -65.795 -107.275 ;
        RECT -66.125 -108.965 -65.795 -108.635 ;
        RECT -66.125 -110.325 -65.795 -109.995 ;
        RECT -66.125 -111.685 -65.795 -111.355 ;
        RECT -66.125 -113.045 -65.795 -112.715 ;
        RECT -66.125 -114.405 -65.795 -114.075 ;
        RECT -66.125 -115.765 -65.795 -115.435 ;
        RECT -66.125 -117.125 -65.795 -116.795 ;
        RECT -66.125 -118.485 -65.795 -118.155 ;
        RECT -66.125 -119.845 -65.795 -119.515 ;
        RECT -66.125 -121.205 -65.795 -120.875 ;
        RECT -66.125 -122.565 -65.795 -122.235 ;
        RECT -66.125 -123.925 -65.795 -123.595 ;
        RECT -66.125 -125.285 -65.795 -124.955 ;
        RECT -66.125 -126.645 -65.795 -126.315 ;
        RECT -66.125 -128.005 -65.795 -127.675 ;
        RECT -66.125 -129.365 -65.795 -129.035 ;
        RECT -66.125 -130.725 -65.795 -130.395 ;
        RECT -66.125 -132.085 -65.795 -131.755 ;
        RECT -66.125 -133.445 -65.795 -133.115 ;
        RECT -66.125 -134.805 -65.795 -134.475 ;
        RECT -66.125 -136.165 -65.795 -135.835 ;
        RECT -66.125 -137.525 -65.795 -137.195 ;
        RECT -66.125 -138.885 -65.795 -138.555 ;
        RECT -66.125 -140.245 -65.795 -139.915 ;
        RECT -66.125 -141.605 -65.795 -141.275 ;
        RECT -66.125 -142.965 -65.795 -142.635 ;
        RECT -66.125 -144.325 -65.795 -143.995 ;
        RECT -66.125 -145.685 -65.795 -145.355 ;
        RECT -66.125 -147.045 -65.795 -146.715 ;
        RECT -66.125 -148.405 -65.795 -148.075 ;
        RECT -66.125 -149.765 -65.795 -149.435 ;
        RECT -66.125 -151.125 -65.795 -150.795 ;
        RECT -66.125 -152.485 -65.795 -152.155 ;
        RECT -66.125 -153.845 -65.795 -153.515 ;
        RECT -66.125 -155.205 -65.795 -154.875 ;
        RECT -66.125 -156.565 -65.795 -156.235 ;
        RECT -66.125 -157.925 -65.795 -157.595 ;
        RECT -66.125 -159.285 -65.795 -158.955 ;
        RECT -66.125 -160.645 -65.795 -160.315 ;
        RECT -66.125 -162.005 -65.795 -161.675 ;
        RECT -66.125 -163.365 -65.795 -163.035 ;
        RECT -66.125 -164.725 -65.795 -164.395 ;
        RECT -66.125 -166.085 -65.795 -165.755 ;
        RECT -66.125 -167.445 -65.795 -167.115 ;
        RECT -66.125 -168.805 -65.795 -168.475 ;
        RECT -66.125 -170.165 -65.795 -169.835 ;
        RECT -66.125 -171.525 -65.795 -171.195 ;
        RECT -66.125 -172.885 -65.795 -172.555 ;
        RECT -66.125 -174.245 -65.795 -173.915 ;
        RECT -66.125 -175.605 -65.795 -175.275 ;
        RECT -66.125 -176.965 -65.795 -176.635 ;
        RECT -66.125 -178.325 -65.795 -177.995 ;
        RECT -66.125 -179.685 -65.795 -179.355 ;
        RECT -66.125 -181.045 -65.795 -180.715 ;
        RECT -66.125 -182.405 -65.795 -182.075 ;
        RECT -66.125 -183.765 -65.795 -183.435 ;
        RECT -66.125 -185.125 -65.795 -184.795 ;
        RECT -66.125 -186.485 -65.795 -186.155 ;
        RECT -66.125 -187.845 -65.795 -187.515 ;
        RECT -66.125 -189.205 -65.795 -188.875 ;
        RECT -66.125 -190.565 -65.795 -190.235 ;
        RECT -66.125 -191.925 -65.795 -191.595 ;
        RECT -66.125 -193.285 -65.795 -192.955 ;
        RECT -66.125 -194.645 -65.795 -194.315 ;
        RECT -66.125 -196.005 -65.795 -195.675 ;
        RECT -66.125 -197.365 -65.795 -197.035 ;
        RECT -66.125 -198.725 -65.795 -198.395 ;
        RECT -66.125 -200.085 -65.795 -199.755 ;
        RECT -66.125 -201.445 -65.795 -201.115 ;
        RECT -66.125 -202.805 -65.795 -202.475 ;
        RECT -66.125 -204.165 -65.795 -203.835 ;
        RECT -66.125 -205.525 -65.795 -205.195 ;
        RECT -66.125 -208.245 -65.795 -207.915 ;
        RECT -66.125 -209.605 -65.795 -209.275 ;
        RECT -66.125 -210.965 -65.795 -210.635 ;
        RECT -66.125 -212.325 -65.795 -211.995 ;
        RECT -66.125 -215.045 -65.795 -214.715 ;
        RECT -66.125 -216.405 -65.795 -216.075 ;
        RECT -66.125 -217.765 -65.795 -217.435 ;
        RECT -66.125 -219.125 -65.795 -218.795 ;
        RECT -66.125 -221.37 -65.795 -220.24 ;
        RECT -66.12 -221.485 -65.8 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -64.765 -99.445 -64.435 -99.115 ;
        RECT -64.765 -100.805 -64.435 -100.475 ;
        RECT -64.765 -102.165 -64.435 -101.835 ;
        RECT -64.765 -103.525 -64.435 -103.195 ;
        RECT -64.765 -104.885 -64.435 -104.555 ;
        RECT -64.765 -106.245 -64.435 -105.915 ;
        RECT -64.765 -107.605 -64.435 -107.275 ;
        RECT -64.765 -108.965 -64.435 -108.635 ;
        RECT -64.765 -110.325 -64.435 -109.995 ;
        RECT -64.765 -111.685 -64.435 -111.355 ;
        RECT -64.765 -113.045 -64.435 -112.715 ;
        RECT -64.765 -114.405 -64.435 -114.075 ;
        RECT -64.765 -115.765 -64.435 -115.435 ;
        RECT -64.765 -117.125 -64.435 -116.795 ;
        RECT -64.765 -118.485 -64.435 -118.155 ;
        RECT -64.765 -119.845 -64.435 -119.515 ;
        RECT -64.765 -121.205 -64.435 -120.875 ;
        RECT -64.765 -122.565 -64.435 -122.235 ;
        RECT -64.765 -123.925 -64.435 -123.595 ;
        RECT -64.765 -125.285 -64.435 -124.955 ;
        RECT -64.765 -126.645 -64.435 -126.315 ;
        RECT -64.765 -128.005 -64.435 -127.675 ;
        RECT -64.765 -129.365 -64.435 -129.035 ;
        RECT -64.765 -130.725 -64.435 -130.395 ;
        RECT -64.765 -132.085 -64.435 -131.755 ;
        RECT -64.765 -133.445 -64.435 -133.115 ;
        RECT -64.765 -134.805 -64.435 -134.475 ;
        RECT -64.765 -136.165 -64.435 -135.835 ;
        RECT -64.765 -137.525 -64.435 -137.195 ;
        RECT -64.765 -138.885 -64.435 -138.555 ;
        RECT -64.765 -140.245 -64.435 -139.915 ;
        RECT -64.765 -141.605 -64.435 -141.275 ;
        RECT -64.765 -142.965 -64.435 -142.635 ;
        RECT -64.765 -144.325 -64.435 -143.995 ;
        RECT -64.765 -145.685 -64.435 -145.355 ;
        RECT -64.765 -147.045 -64.435 -146.715 ;
        RECT -64.765 -148.405 -64.435 -148.075 ;
        RECT -64.765 -149.765 -64.435 -149.435 ;
        RECT -64.765 -151.125 -64.435 -150.795 ;
        RECT -64.765 -152.485 -64.435 -152.155 ;
        RECT -64.765 -153.845 -64.435 -153.515 ;
        RECT -64.765 -155.205 -64.435 -154.875 ;
        RECT -64.765 -156.565 -64.435 -156.235 ;
        RECT -64.765 -157.925 -64.435 -157.595 ;
        RECT -64.765 -159.285 -64.435 -158.955 ;
        RECT -64.765 -160.645 -64.435 -160.315 ;
        RECT -64.765 -162.005 -64.435 -161.675 ;
        RECT -64.765 -163.365 -64.435 -163.035 ;
        RECT -64.765 -164.725 -64.435 -164.395 ;
        RECT -64.765 -166.085 -64.435 -165.755 ;
        RECT -64.765 -167.445 -64.435 -167.115 ;
        RECT -64.765 -168.805 -64.435 -168.475 ;
        RECT -64.765 -170.165 -64.435 -169.835 ;
        RECT -64.765 -171.525 -64.435 -171.195 ;
        RECT -64.765 -172.885 -64.435 -172.555 ;
        RECT -64.765 -174.245 -64.435 -173.915 ;
        RECT -64.765 -175.605 -64.435 -175.275 ;
        RECT -64.765 -176.965 -64.435 -176.635 ;
        RECT -64.765 -178.325 -64.435 -177.995 ;
        RECT -64.765 -179.685 -64.435 -179.355 ;
        RECT -64.765 -181.045 -64.435 -180.715 ;
        RECT -64.765 -182.405 -64.435 -182.075 ;
        RECT -64.765 -183.765 -64.435 -183.435 ;
        RECT -64.765 -185.125 -64.435 -184.795 ;
        RECT -64.765 -186.485 -64.435 -186.155 ;
        RECT -64.765 -187.845 -64.435 -187.515 ;
        RECT -64.765 -189.205 -64.435 -188.875 ;
        RECT -64.765 -190.565 -64.435 -190.235 ;
        RECT -64.765 -191.925 -64.435 -191.595 ;
        RECT -64.765 -193.285 -64.435 -192.955 ;
        RECT -64.765 -194.645 -64.435 -194.315 ;
        RECT -64.765 -196.005 -64.435 -195.675 ;
        RECT -64.765 -197.365 -64.435 -197.035 ;
        RECT -64.765 -198.725 -64.435 -198.395 ;
        RECT -64.765 -200.085 -64.435 -199.755 ;
        RECT -64.765 -201.445 -64.435 -201.115 ;
        RECT -64.765 -202.805 -64.435 -202.475 ;
        RECT -64.765 -204.165 -64.435 -203.835 ;
        RECT -64.765 -205.525 -64.435 -205.195 ;
        RECT -64.765 -208.245 -64.435 -207.915 ;
        RECT -64.765 -209.605 -64.435 -209.275 ;
        RECT -64.76 -209.605 -64.44 131.045 ;
        RECT -64.765 129.8 -64.435 130.93 ;
        RECT -64.765 127.675 -64.435 128.005 ;
        RECT -64.765 126.315 -64.435 126.645 ;
        RECT -64.765 124.955 -64.435 125.285 ;
        RECT -64.765 123.595 -64.435 123.925 ;
        RECT -64.765 122.235 -64.435 122.565 ;
        RECT -64.765 120.875 -64.435 121.205 ;
        RECT -64.765 119.515 -64.435 119.845 ;
        RECT -64.765 118.155 -64.435 118.485 ;
        RECT -64.765 116.795 -64.435 117.125 ;
        RECT -64.765 115.435 -64.435 115.765 ;
        RECT -64.765 114.075 -64.435 114.405 ;
        RECT -64.765 112.715 -64.435 113.045 ;
        RECT -64.765 111.355 -64.435 111.685 ;
        RECT -64.765 109.995 -64.435 110.325 ;
        RECT -64.765 108.635 -64.435 108.965 ;
        RECT -64.765 107.275 -64.435 107.605 ;
        RECT -64.765 105.915 -64.435 106.245 ;
        RECT -64.765 104.555 -64.435 104.885 ;
        RECT -64.765 103.195 -64.435 103.525 ;
        RECT -64.765 101.835 -64.435 102.165 ;
        RECT -64.765 100.475 -64.435 100.805 ;
        RECT -64.765 99.115 -64.435 99.445 ;
        RECT -64.765 97.755 -64.435 98.085 ;
        RECT -64.765 96.395 -64.435 96.725 ;
        RECT -64.765 95.035 -64.435 95.365 ;
        RECT -64.765 93.675 -64.435 94.005 ;
        RECT -64.765 92.315 -64.435 92.645 ;
        RECT -64.765 90.955 -64.435 91.285 ;
        RECT -64.765 89.595 -64.435 89.925 ;
        RECT -64.765 88.235 -64.435 88.565 ;
        RECT -64.765 86.875 -64.435 87.205 ;
        RECT -64.765 85.515 -64.435 85.845 ;
        RECT -64.765 84.155 -64.435 84.485 ;
        RECT -64.765 82.795 -64.435 83.125 ;
        RECT -64.765 81.435 -64.435 81.765 ;
        RECT -64.765 80.075 -64.435 80.405 ;
        RECT -64.765 78.715 -64.435 79.045 ;
        RECT -64.765 77.355 -64.435 77.685 ;
        RECT -64.765 75.995 -64.435 76.325 ;
        RECT -64.765 74.635 -64.435 74.965 ;
        RECT -64.765 73.275 -64.435 73.605 ;
        RECT -64.765 71.915 -64.435 72.245 ;
        RECT -64.765 70.555 -64.435 70.885 ;
        RECT -64.765 69.195 -64.435 69.525 ;
        RECT -64.765 67.835 -64.435 68.165 ;
        RECT -64.765 66.475 -64.435 66.805 ;
        RECT -64.765 65.115 -64.435 65.445 ;
        RECT -64.765 63.755 -64.435 64.085 ;
        RECT -64.765 62.395 -64.435 62.725 ;
        RECT -64.765 61.035 -64.435 61.365 ;
        RECT -64.765 59.675 -64.435 60.005 ;
        RECT -64.765 58.315 -64.435 58.645 ;
        RECT -64.765 56.955 -64.435 57.285 ;
        RECT -64.765 55.595 -64.435 55.925 ;
        RECT -64.765 54.235 -64.435 54.565 ;
        RECT -64.765 52.875 -64.435 53.205 ;
        RECT -64.765 51.515 -64.435 51.845 ;
        RECT -64.765 50.155 -64.435 50.485 ;
        RECT -64.765 48.795 -64.435 49.125 ;
        RECT -64.765 47.435 -64.435 47.765 ;
        RECT -64.765 46.075 -64.435 46.405 ;
        RECT -64.765 44.715 -64.435 45.045 ;
        RECT -64.765 43.355 -64.435 43.685 ;
        RECT -64.765 41.995 -64.435 42.325 ;
        RECT -64.765 40.635 -64.435 40.965 ;
        RECT -64.765 39.275 -64.435 39.605 ;
        RECT -64.765 37.915 -64.435 38.245 ;
        RECT -64.765 36.555 -64.435 36.885 ;
        RECT -64.765 35.195 -64.435 35.525 ;
        RECT -64.765 33.835 -64.435 34.165 ;
        RECT -64.765 32.475 -64.435 32.805 ;
        RECT -64.765 31.115 -64.435 31.445 ;
        RECT -64.765 29.755 -64.435 30.085 ;
        RECT -64.765 28.395 -64.435 28.725 ;
        RECT -64.765 27.035 -64.435 27.365 ;
        RECT -64.765 25.675 -64.435 26.005 ;
        RECT -64.765 24.315 -64.435 24.645 ;
        RECT -64.765 22.955 -64.435 23.285 ;
        RECT -64.765 21.595 -64.435 21.925 ;
        RECT -64.765 20.235 -64.435 20.565 ;
        RECT -64.765 18.875 -64.435 19.205 ;
        RECT -64.765 17.515 -64.435 17.845 ;
        RECT -64.765 16.155 -64.435 16.485 ;
        RECT -64.765 14.795 -64.435 15.125 ;
        RECT -64.765 13.435 -64.435 13.765 ;
        RECT -64.765 12.075 -64.435 12.405 ;
        RECT -64.765 10.715 -64.435 11.045 ;
        RECT -64.765 9.355 -64.435 9.685 ;
        RECT -64.765 7.995 -64.435 8.325 ;
        RECT -64.765 6.635 -64.435 6.965 ;
        RECT -64.765 5.275 -64.435 5.605 ;
        RECT -64.765 3.915 -64.435 4.245 ;
        RECT -64.765 2.555 -64.435 2.885 ;
        RECT -64.765 1.195 -64.435 1.525 ;
        RECT -64.765 -0.165 -64.435 0.165 ;
        RECT -64.765 -1.525 -64.435 -1.195 ;
        RECT -64.765 -2.885 -64.435 -2.555 ;
        RECT -64.765 -4.245 -64.435 -3.915 ;
        RECT -64.765 -5.605 -64.435 -5.275 ;
        RECT -64.765 -6.965 -64.435 -6.635 ;
        RECT -64.765 -8.325 -64.435 -7.995 ;
        RECT -64.765 -9.685 -64.435 -9.355 ;
        RECT -64.765 -11.045 -64.435 -10.715 ;
        RECT -64.765 -12.405 -64.435 -12.075 ;
        RECT -64.765 -13.765 -64.435 -13.435 ;
        RECT -64.765 -15.125 -64.435 -14.795 ;
        RECT -64.765 -16.485 -64.435 -16.155 ;
        RECT -64.765 -17.845 -64.435 -17.515 ;
        RECT -64.765 -19.205 -64.435 -18.875 ;
        RECT -64.765 -20.565 -64.435 -20.235 ;
        RECT -64.765 -21.925 -64.435 -21.595 ;
        RECT -64.765 -23.285 -64.435 -22.955 ;
        RECT -64.765 -24.645 -64.435 -24.315 ;
        RECT -64.765 -26.005 -64.435 -25.675 ;
        RECT -64.765 -27.365 -64.435 -27.035 ;
        RECT -64.765 -28.725 -64.435 -28.395 ;
        RECT -64.765 -30.085 -64.435 -29.755 ;
        RECT -64.765 -31.445 -64.435 -31.115 ;
        RECT -64.765 -32.805 -64.435 -32.475 ;
        RECT -64.765 -34.165 -64.435 -33.835 ;
        RECT -64.765 -35.525 -64.435 -35.195 ;
        RECT -64.765 -36.885 -64.435 -36.555 ;
        RECT -64.765 -38.245 -64.435 -37.915 ;
        RECT -64.765 -39.605 -64.435 -39.275 ;
        RECT -64.765 -40.965 -64.435 -40.635 ;
        RECT -64.765 -42.325 -64.435 -41.995 ;
        RECT -64.765 -43.685 -64.435 -43.355 ;
        RECT -64.765 -45.045 -64.435 -44.715 ;
        RECT -64.765 -46.405 -64.435 -46.075 ;
        RECT -64.765 -47.765 -64.435 -47.435 ;
        RECT -64.765 -49.125 -64.435 -48.795 ;
        RECT -64.765 -50.485 -64.435 -50.155 ;
        RECT -64.765 -51.845 -64.435 -51.515 ;
        RECT -64.765 -53.205 -64.435 -52.875 ;
        RECT -64.765 -54.565 -64.435 -54.235 ;
        RECT -64.765 -55.925 -64.435 -55.595 ;
        RECT -64.765 -57.285 -64.435 -56.955 ;
        RECT -64.765 -58.645 -64.435 -58.315 ;
        RECT -64.765 -60.005 -64.435 -59.675 ;
        RECT -64.765 -61.365 -64.435 -61.035 ;
        RECT -64.765 -62.725 -64.435 -62.395 ;
        RECT -64.765 -64.085 -64.435 -63.755 ;
        RECT -64.765 -65.445 -64.435 -65.115 ;
        RECT -64.765 -66.805 -64.435 -66.475 ;
        RECT -64.765 -68.165 -64.435 -67.835 ;
        RECT -64.765 -69.525 -64.435 -69.195 ;
        RECT -64.765 -70.885 -64.435 -70.555 ;
        RECT -64.765 -72.245 -64.435 -71.915 ;
        RECT -64.765 -73.605 -64.435 -73.275 ;
        RECT -64.765 -74.965 -64.435 -74.635 ;
        RECT -64.765 -76.325 -64.435 -75.995 ;
        RECT -64.765 -77.685 -64.435 -77.355 ;
        RECT -64.765 -79.045 -64.435 -78.715 ;
        RECT -64.765 -80.405 -64.435 -80.075 ;
        RECT -64.765 -81.765 -64.435 -81.435 ;
        RECT -64.765 -83.125 -64.435 -82.795 ;
        RECT -64.765 -84.485 -64.435 -84.155 ;
        RECT -64.765 -85.845 -64.435 -85.515 ;
        RECT -64.765 -87.205 -64.435 -86.875 ;
        RECT -64.765 -88.565 -64.435 -88.235 ;
        RECT -64.765 -89.925 -64.435 -89.595 ;
        RECT -64.765 -91.285 -64.435 -90.955 ;
        RECT -64.765 -92.645 -64.435 -92.315 ;
        RECT -64.765 -94.005 -64.435 -93.675 ;
        RECT -64.765 -95.365 -64.435 -95.035 ;
        RECT -64.765 -96.725 -64.435 -96.395 ;
        RECT -64.765 -98.085 -64.435 -97.755 ;
    END
    PORT
      LAYER met3 ;
        RECT -71.565 129.8 -71.235 130.93 ;
        RECT -71.565 127.675 -71.235 128.005 ;
        RECT -71.565 126.315 -71.235 126.645 ;
        RECT -71.565 124.955 -71.235 125.285 ;
        RECT -71.565 123.595 -71.235 123.925 ;
        RECT -71.565 122.235 -71.235 122.565 ;
        RECT -71.565 120.875 -71.235 121.205 ;
        RECT -71.565 119.515 -71.235 119.845 ;
        RECT -71.565 118.155 -71.235 118.485 ;
        RECT -71.565 116.795 -71.235 117.125 ;
        RECT -71.565 115.435 -71.235 115.765 ;
        RECT -71.565 114.075 -71.235 114.405 ;
        RECT -71.565 112.715 -71.235 113.045 ;
        RECT -71.565 111.355 -71.235 111.685 ;
        RECT -71.565 109.995 -71.235 110.325 ;
        RECT -71.565 108.635 -71.235 108.965 ;
        RECT -71.565 107.275 -71.235 107.605 ;
        RECT -71.565 105.915 -71.235 106.245 ;
        RECT -71.565 104.555 -71.235 104.885 ;
        RECT -71.565 103.195 -71.235 103.525 ;
        RECT -71.565 101.835 -71.235 102.165 ;
        RECT -71.565 100.475 -71.235 100.805 ;
        RECT -71.565 99.115 -71.235 99.445 ;
        RECT -71.565 97.755 -71.235 98.085 ;
        RECT -71.565 96.395 -71.235 96.725 ;
        RECT -71.565 95.035 -71.235 95.365 ;
        RECT -71.565 93.675 -71.235 94.005 ;
        RECT -71.565 92.315 -71.235 92.645 ;
        RECT -71.565 90.955 -71.235 91.285 ;
        RECT -71.565 89.595 -71.235 89.925 ;
        RECT -71.565 88.235 -71.235 88.565 ;
        RECT -71.565 86.875 -71.235 87.205 ;
        RECT -71.565 85.515 -71.235 85.845 ;
        RECT -71.565 84.155 -71.235 84.485 ;
        RECT -71.565 82.795 -71.235 83.125 ;
        RECT -71.565 81.435 -71.235 81.765 ;
        RECT -71.565 80.075 -71.235 80.405 ;
        RECT -71.565 78.715 -71.235 79.045 ;
        RECT -71.565 77.355 -71.235 77.685 ;
        RECT -71.565 75.995 -71.235 76.325 ;
        RECT -71.565 74.635 -71.235 74.965 ;
        RECT -71.565 73.275 -71.235 73.605 ;
        RECT -71.565 71.915 -71.235 72.245 ;
        RECT -71.565 70.555 -71.235 70.885 ;
        RECT -71.565 69.195 -71.235 69.525 ;
        RECT -71.565 67.835 -71.235 68.165 ;
        RECT -71.565 66.475 -71.235 66.805 ;
        RECT -71.565 65.115 -71.235 65.445 ;
        RECT -71.565 63.755 -71.235 64.085 ;
        RECT -71.565 62.395 -71.235 62.725 ;
        RECT -71.565 61.035 -71.235 61.365 ;
        RECT -71.565 59.675 -71.235 60.005 ;
        RECT -71.565 58.315 -71.235 58.645 ;
        RECT -71.565 56.955 -71.235 57.285 ;
        RECT -71.565 55.595 -71.235 55.925 ;
        RECT -71.565 54.235 -71.235 54.565 ;
        RECT -71.565 52.875 -71.235 53.205 ;
        RECT -71.565 51.515 -71.235 51.845 ;
        RECT -71.565 50.155 -71.235 50.485 ;
        RECT -71.565 48.795 -71.235 49.125 ;
        RECT -71.565 47.435 -71.235 47.765 ;
        RECT -71.565 46.075 -71.235 46.405 ;
        RECT -71.565 44.715 -71.235 45.045 ;
        RECT -71.565 43.355 -71.235 43.685 ;
        RECT -71.565 41.995 -71.235 42.325 ;
        RECT -71.565 40.635 -71.235 40.965 ;
        RECT -71.565 39.275 -71.235 39.605 ;
        RECT -71.565 37.915 -71.235 38.245 ;
        RECT -71.565 36.555 -71.235 36.885 ;
        RECT -71.565 35.195 -71.235 35.525 ;
        RECT -71.565 33.835 -71.235 34.165 ;
        RECT -71.565 32.475 -71.235 32.805 ;
        RECT -71.565 31.115 -71.235 31.445 ;
        RECT -71.565 29.755 -71.235 30.085 ;
        RECT -71.565 28.395 -71.235 28.725 ;
        RECT -71.565 27.035 -71.235 27.365 ;
        RECT -71.565 25.675 -71.235 26.005 ;
        RECT -71.565 24.315 -71.235 24.645 ;
        RECT -71.565 22.955 -71.235 23.285 ;
        RECT -71.565 21.595 -71.235 21.925 ;
        RECT -71.565 20.235 -71.235 20.565 ;
        RECT -71.565 18.875 -71.235 19.205 ;
        RECT -71.565 17.515 -71.235 17.845 ;
        RECT -71.565 16.155 -71.235 16.485 ;
        RECT -71.565 14.795 -71.235 15.125 ;
        RECT -71.565 13.435 -71.235 13.765 ;
        RECT -71.565 12.075 -71.235 12.405 ;
        RECT -71.565 10.715 -71.235 11.045 ;
        RECT -71.565 9.355 -71.235 9.685 ;
        RECT -71.565 7.995 -71.235 8.325 ;
        RECT -71.565 6.635 -71.235 6.965 ;
        RECT -71.565 5.275 -71.235 5.605 ;
        RECT -71.565 3.915 -71.235 4.245 ;
        RECT -71.565 2.555 -71.235 2.885 ;
        RECT -71.565 1.195 -71.235 1.525 ;
        RECT -71.565 -0.165 -71.235 0.165 ;
        RECT -71.565 -1.525 -71.235 -1.195 ;
        RECT -71.565 -2.885 -71.235 -2.555 ;
        RECT -71.565 -4.245 -71.235 -3.915 ;
        RECT -71.565 -5.605 -71.235 -5.275 ;
        RECT -71.565 -6.965 -71.235 -6.635 ;
        RECT -71.565 -8.325 -71.235 -7.995 ;
        RECT -71.565 -9.685 -71.235 -9.355 ;
        RECT -71.565 -11.045 -71.235 -10.715 ;
        RECT -71.565 -12.405 -71.235 -12.075 ;
        RECT -71.565 -13.765 -71.235 -13.435 ;
        RECT -71.565 -15.125 -71.235 -14.795 ;
        RECT -71.565 -16.485 -71.235 -16.155 ;
        RECT -71.565 -17.845 -71.235 -17.515 ;
        RECT -71.565 -19.205 -71.235 -18.875 ;
        RECT -71.565 -20.565 -71.235 -20.235 ;
        RECT -71.565 -21.925 -71.235 -21.595 ;
        RECT -71.565 -23.285 -71.235 -22.955 ;
        RECT -71.565 -24.645 -71.235 -24.315 ;
        RECT -71.565 -26.005 -71.235 -25.675 ;
        RECT -71.565 -27.365 -71.235 -27.035 ;
        RECT -71.565 -28.725 -71.235 -28.395 ;
        RECT -71.565 -30.085 -71.235 -29.755 ;
        RECT -71.565 -31.445 -71.235 -31.115 ;
        RECT -71.565 -32.805 -71.235 -32.475 ;
        RECT -71.565 -34.165 -71.235 -33.835 ;
        RECT -71.565 -35.525 -71.235 -35.195 ;
        RECT -71.565 -36.885 -71.235 -36.555 ;
        RECT -71.565 -38.245 -71.235 -37.915 ;
        RECT -71.565 -39.605 -71.235 -39.275 ;
        RECT -71.565 -40.965 -71.235 -40.635 ;
        RECT -71.565 -42.325 -71.235 -41.995 ;
        RECT -71.565 -43.685 -71.235 -43.355 ;
        RECT -71.565 -45.045 -71.235 -44.715 ;
        RECT -71.565 -46.405 -71.235 -46.075 ;
        RECT -71.565 -47.765 -71.235 -47.435 ;
        RECT -71.565 -49.125 -71.235 -48.795 ;
        RECT -71.565 -50.485 -71.235 -50.155 ;
        RECT -71.565 -51.845 -71.235 -51.515 ;
        RECT -71.565 -53.205 -71.235 -52.875 ;
        RECT -71.565 -54.565 -71.235 -54.235 ;
        RECT -71.565 -55.925 -71.235 -55.595 ;
        RECT -71.565 -57.285 -71.235 -56.955 ;
        RECT -71.565 -58.645 -71.235 -58.315 ;
        RECT -71.565 -60.005 -71.235 -59.675 ;
        RECT -71.565 -61.365 -71.235 -61.035 ;
        RECT -71.565 -62.725 -71.235 -62.395 ;
        RECT -71.565 -64.085 -71.235 -63.755 ;
        RECT -71.565 -65.445 -71.235 -65.115 ;
        RECT -71.565 -66.805 -71.235 -66.475 ;
        RECT -71.565 -68.165 -71.235 -67.835 ;
        RECT -71.565 -69.525 -71.235 -69.195 ;
        RECT -71.565 -70.885 -71.235 -70.555 ;
        RECT -71.565 -72.245 -71.235 -71.915 ;
        RECT -71.565 -73.605 -71.235 -73.275 ;
        RECT -71.565 -74.965 -71.235 -74.635 ;
        RECT -71.565 -76.325 -71.235 -75.995 ;
        RECT -71.565 -77.685 -71.235 -77.355 ;
        RECT -71.565 -79.045 -71.235 -78.715 ;
        RECT -71.565 -80.405 -71.235 -80.075 ;
        RECT -71.565 -81.765 -71.235 -81.435 ;
        RECT -71.565 -83.125 -71.235 -82.795 ;
        RECT -71.565 -84.485 -71.235 -84.155 ;
        RECT -71.565 -85.845 -71.235 -85.515 ;
        RECT -71.565 -87.205 -71.235 -86.875 ;
        RECT -71.565 -88.565 -71.235 -88.235 ;
        RECT -71.565 -89.925 -71.235 -89.595 ;
        RECT -71.565 -91.285 -71.235 -90.955 ;
        RECT -71.565 -92.645 -71.235 -92.315 ;
        RECT -71.565 -94.005 -71.235 -93.675 ;
        RECT -71.565 -95.365 -71.235 -95.035 ;
        RECT -71.565 -96.725 -71.235 -96.395 ;
        RECT -71.565 -98.085 -71.235 -97.755 ;
        RECT -71.565 -99.445 -71.235 -99.115 ;
        RECT -71.565 -100.805 -71.235 -100.475 ;
        RECT -71.565 -102.165 -71.235 -101.835 ;
        RECT -71.565 -103.525 -71.235 -103.195 ;
        RECT -71.565 -104.885 -71.235 -104.555 ;
        RECT -71.565 -106.245 -71.235 -105.915 ;
        RECT -71.565 -107.605 -71.235 -107.275 ;
        RECT -71.565 -108.965 -71.235 -108.635 ;
        RECT -71.565 -110.325 -71.235 -109.995 ;
        RECT -71.565 -111.685 -71.235 -111.355 ;
        RECT -71.565 -113.045 -71.235 -112.715 ;
        RECT -71.565 -114.405 -71.235 -114.075 ;
        RECT -71.565 -115.765 -71.235 -115.435 ;
        RECT -71.565 -117.125 -71.235 -116.795 ;
        RECT -71.565 -118.485 -71.235 -118.155 ;
        RECT -71.565 -119.845 -71.235 -119.515 ;
        RECT -71.565 -121.205 -71.235 -120.875 ;
        RECT -71.565 -122.565 -71.235 -122.235 ;
        RECT -71.565 -123.925 -71.235 -123.595 ;
        RECT -71.565 -125.285 -71.235 -124.955 ;
        RECT -71.565 -126.645 -71.235 -126.315 ;
        RECT -71.565 -128.005 -71.235 -127.675 ;
        RECT -71.565 -129.365 -71.235 -129.035 ;
        RECT -71.565 -130.725 -71.235 -130.395 ;
        RECT -71.565 -132.085 -71.235 -131.755 ;
        RECT -71.565 -133.445 -71.235 -133.115 ;
        RECT -71.565 -134.805 -71.235 -134.475 ;
        RECT -71.565 -136.165 -71.235 -135.835 ;
        RECT -71.565 -137.525 -71.235 -137.195 ;
        RECT -71.565 -138.885 -71.235 -138.555 ;
        RECT -71.565 -140.245 -71.235 -139.915 ;
        RECT -71.565 -141.605 -71.235 -141.275 ;
        RECT -71.565 -142.965 -71.235 -142.635 ;
        RECT -71.565 -144.325 -71.235 -143.995 ;
        RECT -71.565 -145.685 -71.235 -145.355 ;
        RECT -71.565 -147.045 -71.235 -146.715 ;
        RECT -71.565 -148.405 -71.235 -148.075 ;
        RECT -71.565 -149.765 -71.235 -149.435 ;
        RECT -71.565 -151.125 -71.235 -150.795 ;
        RECT -71.565 -152.485 -71.235 -152.155 ;
        RECT -71.565 -153.845 -71.235 -153.515 ;
        RECT -71.565 -155.205 -71.235 -154.875 ;
        RECT -71.565 -156.565 -71.235 -156.235 ;
        RECT -71.565 -157.925 -71.235 -157.595 ;
        RECT -71.565 -159.285 -71.235 -158.955 ;
        RECT -71.565 -160.645 -71.235 -160.315 ;
        RECT -71.565 -162.005 -71.235 -161.675 ;
        RECT -71.565 -163.365 -71.235 -163.035 ;
        RECT -71.565 -164.725 -71.235 -164.395 ;
        RECT -71.565 -166.085 -71.235 -165.755 ;
        RECT -71.565 -167.445 -71.235 -167.115 ;
        RECT -71.565 -168.805 -71.235 -168.475 ;
        RECT -71.565 -170.165 -71.235 -169.835 ;
        RECT -71.565 -171.525 -71.235 -171.195 ;
        RECT -71.565 -172.885 -71.235 -172.555 ;
        RECT -71.565 -174.245 -71.235 -173.915 ;
        RECT -71.565 -175.605 -71.235 -175.275 ;
        RECT -71.565 -176.965 -71.235 -176.635 ;
        RECT -71.565 -178.325 -71.235 -177.995 ;
        RECT -71.565 -179.685 -71.235 -179.355 ;
        RECT -71.565 -181.045 -71.235 -180.715 ;
        RECT -71.565 -182.405 -71.235 -182.075 ;
        RECT -71.565 -183.765 -71.235 -183.435 ;
        RECT -71.565 -185.125 -71.235 -184.795 ;
        RECT -71.565 -186.485 -71.235 -186.155 ;
        RECT -71.565 -187.845 -71.235 -187.515 ;
        RECT -71.565 -189.205 -71.235 -188.875 ;
        RECT -71.565 -190.565 -71.235 -190.235 ;
        RECT -71.565 -191.925 -71.235 -191.595 ;
        RECT -71.565 -193.285 -71.235 -192.955 ;
        RECT -71.565 -194.645 -71.235 -194.315 ;
        RECT -71.565 -196.005 -71.235 -195.675 ;
        RECT -71.565 -197.365 -71.235 -197.035 ;
        RECT -71.565 -198.725 -71.235 -198.395 ;
        RECT -71.565 -200.085 -71.235 -199.755 ;
        RECT -71.565 -201.445 -71.235 -201.115 ;
        RECT -71.565 -202.805 -71.235 -202.475 ;
        RECT -71.565 -204.165 -71.235 -203.835 ;
        RECT -71.565 -205.525 -71.235 -205.195 ;
        RECT -71.565 -206.885 -71.235 -206.555 ;
        RECT -71.565 -208.245 -71.235 -207.915 ;
        RECT -71.565 -209.605 -71.235 -209.275 ;
        RECT -71.565 -210.965 -71.235 -210.635 ;
        RECT -71.565 -212.325 -71.235 -211.995 ;
        RECT -71.565 -213.685 -71.235 -213.355 ;
        RECT -71.565 -215.045 -71.235 -214.715 ;
        RECT -71.565 -216.405 -71.235 -216.075 ;
        RECT -71.565 -217.765 -71.235 -217.435 ;
        RECT -71.565 -219.125 -71.235 -218.795 ;
        RECT -71.565 -221.37 -71.235 -220.24 ;
        RECT -71.56 -221.485 -71.24 131.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -70.205 -65.445 -69.875 -65.115 ;
        RECT -70.205 -66.805 -69.875 -66.475 ;
        RECT -70.205 -68.165 -69.875 -67.835 ;
        RECT -70.205 -69.525 -69.875 -69.195 ;
        RECT -70.205 -70.885 -69.875 -70.555 ;
        RECT -70.205 -72.245 -69.875 -71.915 ;
        RECT -70.205 -73.605 -69.875 -73.275 ;
        RECT -70.205 -74.965 -69.875 -74.635 ;
        RECT -70.205 -76.325 -69.875 -75.995 ;
        RECT -70.205 -77.685 -69.875 -77.355 ;
        RECT -70.205 -79.045 -69.875 -78.715 ;
        RECT -70.205 -80.405 -69.875 -80.075 ;
        RECT -70.205 -81.765 -69.875 -81.435 ;
        RECT -70.205 -83.125 -69.875 -82.795 ;
        RECT -70.205 -84.485 -69.875 -84.155 ;
        RECT -70.205 -85.845 -69.875 -85.515 ;
        RECT -70.205 -87.205 -69.875 -86.875 ;
        RECT -70.205 -88.565 -69.875 -88.235 ;
        RECT -70.205 -89.925 -69.875 -89.595 ;
        RECT -70.205 -91.285 -69.875 -90.955 ;
        RECT -70.205 -92.645 -69.875 -92.315 ;
        RECT -70.205 -94.005 -69.875 -93.675 ;
        RECT -70.205 -95.365 -69.875 -95.035 ;
        RECT -70.205 -96.725 -69.875 -96.395 ;
        RECT -70.205 -98.085 -69.875 -97.755 ;
        RECT -70.205 -99.445 -69.875 -99.115 ;
        RECT -70.205 -100.805 -69.875 -100.475 ;
        RECT -70.205 -102.165 -69.875 -101.835 ;
        RECT -70.205 -103.525 -69.875 -103.195 ;
        RECT -70.205 -104.885 -69.875 -104.555 ;
        RECT -70.205 -106.245 -69.875 -105.915 ;
        RECT -70.205 -107.605 -69.875 -107.275 ;
        RECT -70.205 -108.965 -69.875 -108.635 ;
        RECT -70.205 -110.325 -69.875 -109.995 ;
        RECT -70.205 -111.685 -69.875 -111.355 ;
        RECT -70.205 -113.045 -69.875 -112.715 ;
        RECT -70.205 -114.405 -69.875 -114.075 ;
        RECT -70.205 -115.765 -69.875 -115.435 ;
        RECT -70.205 -117.125 -69.875 -116.795 ;
        RECT -70.205 -118.485 -69.875 -118.155 ;
        RECT -70.205 -119.845 -69.875 -119.515 ;
        RECT -70.205 -121.205 -69.875 -120.875 ;
        RECT -70.205 -122.565 -69.875 -122.235 ;
        RECT -70.205 -123.925 -69.875 -123.595 ;
        RECT -70.205 -125.285 -69.875 -124.955 ;
        RECT -70.205 -126.645 -69.875 -126.315 ;
        RECT -70.205 -128.005 -69.875 -127.675 ;
        RECT -70.205 -129.365 -69.875 -129.035 ;
        RECT -70.205 -130.725 -69.875 -130.395 ;
        RECT -70.205 -132.085 -69.875 -131.755 ;
        RECT -70.205 -133.445 -69.875 -133.115 ;
        RECT -70.205 -134.805 -69.875 -134.475 ;
        RECT -70.205 -136.165 -69.875 -135.835 ;
        RECT -70.205 -137.525 -69.875 -137.195 ;
        RECT -70.205 -138.885 -69.875 -138.555 ;
        RECT -70.205 -140.245 -69.875 -139.915 ;
        RECT -70.205 -141.605 -69.875 -141.275 ;
        RECT -70.205 -142.965 -69.875 -142.635 ;
        RECT -70.205 -144.325 -69.875 -143.995 ;
        RECT -70.205 -145.685 -69.875 -145.355 ;
        RECT -70.205 -147.045 -69.875 -146.715 ;
        RECT -70.205 -148.405 -69.875 -148.075 ;
        RECT -70.205 -149.765 -69.875 -149.435 ;
        RECT -70.205 -151.125 -69.875 -150.795 ;
        RECT -70.205 -152.485 -69.875 -152.155 ;
        RECT -70.205 -153.845 -69.875 -153.515 ;
        RECT -70.205 -155.205 -69.875 -154.875 ;
        RECT -70.205 -156.565 -69.875 -156.235 ;
        RECT -70.205 -157.925 -69.875 -157.595 ;
        RECT -70.205 -159.285 -69.875 -158.955 ;
        RECT -70.205 -160.645 -69.875 -160.315 ;
        RECT -70.205 -162.005 -69.875 -161.675 ;
        RECT -70.205 -163.365 -69.875 -163.035 ;
        RECT -70.205 -164.725 -69.875 -164.395 ;
        RECT -70.205 -166.085 -69.875 -165.755 ;
        RECT -70.205 -167.445 -69.875 -167.115 ;
        RECT -70.205 -168.805 -69.875 -168.475 ;
        RECT -70.205 -170.165 -69.875 -169.835 ;
        RECT -70.205 -171.525 -69.875 -171.195 ;
        RECT -70.205 -172.885 -69.875 -172.555 ;
        RECT -70.205 -174.245 -69.875 -173.915 ;
        RECT -70.205 -175.605 -69.875 -175.275 ;
        RECT -70.205 -176.965 -69.875 -176.635 ;
        RECT -70.205 -178.325 -69.875 -177.995 ;
        RECT -70.205 -179.685 -69.875 -179.355 ;
        RECT -70.205 -181.045 -69.875 -180.715 ;
        RECT -70.205 -182.405 -69.875 -182.075 ;
        RECT -70.205 -183.765 -69.875 -183.435 ;
        RECT -70.205 -185.125 -69.875 -184.795 ;
        RECT -70.205 -186.485 -69.875 -186.155 ;
        RECT -70.205 -187.845 -69.875 -187.515 ;
        RECT -70.205 -189.205 -69.875 -188.875 ;
        RECT -70.205 -190.565 -69.875 -190.235 ;
        RECT -70.205 -191.925 -69.875 -191.595 ;
        RECT -70.205 -193.285 -69.875 -192.955 ;
        RECT -70.205 -194.645 -69.875 -194.315 ;
        RECT -70.205 -196.005 -69.875 -195.675 ;
        RECT -70.205 -197.365 -69.875 -197.035 ;
        RECT -70.205 -198.725 -69.875 -198.395 ;
        RECT -70.205 -200.085 -69.875 -199.755 ;
        RECT -70.205 -201.445 -69.875 -201.115 ;
        RECT -70.205 -202.805 -69.875 -202.475 ;
        RECT -70.205 -204.165 -69.875 -203.835 ;
        RECT -70.205 -205.525 -69.875 -205.195 ;
        RECT -70.205 -206.885 -69.875 -206.555 ;
        RECT -70.205 -208.245 -69.875 -207.915 ;
        RECT -70.205 -209.605 -69.875 -209.275 ;
        RECT -70.205 -210.965 -69.875 -210.635 ;
        RECT -70.205 -212.325 -69.875 -211.995 ;
        RECT -70.205 -213.685 -69.875 -213.355 ;
        RECT -70.205 -215.045 -69.875 -214.715 ;
        RECT -70.205 -216.405 -69.875 -216.075 ;
        RECT -70.205 -217.765 -69.875 -217.435 ;
        RECT -70.205 -219.125 -69.875 -218.795 ;
        RECT -70.205 -221.37 -69.875 -220.24 ;
        RECT -70.2 -221.485 -69.88 131.045 ;
        RECT -70.205 129.8 -69.875 130.93 ;
        RECT -70.205 127.675 -69.875 128.005 ;
        RECT -70.205 126.315 -69.875 126.645 ;
        RECT -70.205 124.955 -69.875 125.285 ;
        RECT -70.205 123.595 -69.875 123.925 ;
        RECT -70.205 122.235 -69.875 122.565 ;
        RECT -70.205 120.875 -69.875 121.205 ;
        RECT -70.205 119.515 -69.875 119.845 ;
        RECT -70.205 118.155 -69.875 118.485 ;
        RECT -70.205 116.795 -69.875 117.125 ;
        RECT -70.205 115.435 -69.875 115.765 ;
        RECT -70.205 114.075 -69.875 114.405 ;
        RECT -70.205 112.715 -69.875 113.045 ;
        RECT -70.205 111.355 -69.875 111.685 ;
        RECT -70.205 109.995 -69.875 110.325 ;
        RECT -70.205 108.635 -69.875 108.965 ;
        RECT -70.205 107.275 -69.875 107.605 ;
        RECT -70.205 105.915 -69.875 106.245 ;
        RECT -70.205 104.555 -69.875 104.885 ;
        RECT -70.205 103.195 -69.875 103.525 ;
        RECT -70.205 101.835 -69.875 102.165 ;
        RECT -70.205 100.475 -69.875 100.805 ;
        RECT -70.205 99.115 -69.875 99.445 ;
        RECT -70.205 97.755 -69.875 98.085 ;
        RECT -70.205 96.395 -69.875 96.725 ;
        RECT -70.205 95.035 -69.875 95.365 ;
        RECT -70.205 93.675 -69.875 94.005 ;
        RECT -70.205 92.315 -69.875 92.645 ;
        RECT -70.205 90.955 -69.875 91.285 ;
        RECT -70.205 89.595 -69.875 89.925 ;
        RECT -70.205 88.235 -69.875 88.565 ;
        RECT -70.205 86.875 -69.875 87.205 ;
        RECT -70.205 85.515 -69.875 85.845 ;
        RECT -70.205 84.155 -69.875 84.485 ;
        RECT -70.205 82.795 -69.875 83.125 ;
        RECT -70.205 81.435 -69.875 81.765 ;
        RECT -70.205 80.075 -69.875 80.405 ;
        RECT -70.205 78.715 -69.875 79.045 ;
        RECT -70.205 77.355 -69.875 77.685 ;
        RECT -70.205 75.995 -69.875 76.325 ;
        RECT -70.205 74.635 -69.875 74.965 ;
        RECT -70.205 73.275 -69.875 73.605 ;
        RECT -70.205 71.915 -69.875 72.245 ;
        RECT -70.205 70.555 -69.875 70.885 ;
        RECT -70.205 69.195 -69.875 69.525 ;
        RECT -70.205 67.835 -69.875 68.165 ;
        RECT -70.205 66.475 -69.875 66.805 ;
        RECT -70.205 65.115 -69.875 65.445 ;
        RECT -70.205 63.755 -69.875 64.085 ;
        RECT -70.205 62.395 -69.875 62.725 ;
        RECT -70.205 61.035 -69.875 61.365 ;
        RECT -70.205 59.675 -69.875 60.005 ;
        RECT -70.205 58.315 -69.875 58.645 ;
        RECT -70.205 56.955 -69.875 57.285 ;
        RECT -70.205 55.595 -69.875 55.925 ;
        RECT -70.205 54.235 -69.875 54.565 ;
        RECT -70.205 52.875 -69.875 53.205 ;
        RECT -70.205 51.515 -69.875 51.845 ;
        RECT -70.205 50.155 -69.875 50.485 ;
        RECT -70.205 48.795 -69.875 49.125 ;
        RECT -70.205 47.435 -69.875 47.765 ;
        RECT -70.205 46.075 -69.875 46.405 ;
        RECT -70.205 44.715 -69.875 45.045 ;
        RECT -70.205 43.355 -69.875 43.685 ;
        RECT -70.205 41.995 -69.875 42.325 ;
        RECT -70.205 40.635 -69.875 40.965 ;
        RECT -70.205 39.275 -69.875 39.605 ;
        RECT -70.205 37.915 -69.875 38.245 ;
        RECT -70.205 36.555 -69.875 36.885 ;
        RECT -70.205 35.195 -69.875 35.525 ;
        RECT -70.205 33.835 -69.875 34.165 ;
        RECT -70.205 32.475 -69.875 32.805 ;
        RECT -70.205 31.115 -69.875 31.445 ;
        RECT -70.205 29.755 -69.875 30.085 ;
        RECT -70.205 28.395 -69.875 28.725 ;
        RECT -70.205 27.035 -69.875 27.365 ;
        RECT -70.205 25.675 -69.875 26.005 ;
        RECT -70.205 24.315 -69.875 24.645 ;
        RECT -70.205 22.955 -69.875 23.285 ;
        RECT -70.205 21.595 -69.875 21.925 ;
        RECT -70.205 20.235 -69.875 20.565 ;
        RECT -70.205 18.875 -69.875 19.205 ;
        RECT -70.205 17.515 -69.875 17.845 ;
        RECT -70.205 16.155 -69.875 16.485 ;
        RECT -70.205 14.795 -69.875 15.125 ;
        RECT -70.205 13.435 -69.875 13.765 ;
        RECT -70.205 12.075 -69.875 12.405 ;
        RECT -70.205 10.715 -69.875 11.045 ;
        RECT -70.205 9.355 -69.875 9.685 ;
        RECT -70.205 7.995 -69.875 8.325 ;
        RECT -70.205 6.635 -69.875 6.965 ;
        RECT -70.205 5.275 -69.875 5.605 ;
        RECT -70.205 3.915 -69.875 4.245 ;
        RECT -70.205 2.555 -69.875 2.885 ;
        RECT -70.205 1.195 -69.875 1.525 ;
        RECT -70.205 -0.165 -69.875 0.165 ;
        RECT -70.205 -1.525 -69.875 -1.195 ;
        RECT -70.205 -2.885 -69.875 -2.555 ;
        RECT -70.205 -4.245 -69.875 -3.915 ;
        RECT -70.205 -5.605 -69.875 -5.275 ;
        RECT -70.205 -6.965 -69.875 -6.635 ;
        RECT -70.205 -8.325 -69.875 -7.995 ;
        RECT -70.205 -9.685 -69.875 -9.355 ;
        RECT -70.205 -11.045 -69.875 -10.715 ;
        RECT -70.205 -12.405 -69.875 -12.075 ;
        RECT -70.205 -13.765 -69.875 -13.435 ;
        RECT -70.205 -15.125 -69.875 -14.795 ;
        RECT -70.205 -16.485 -69.875 -16.155 ;
        RECT -70.205 -17.845 -69.875 -17.515 ;
        RECT -70.205 -19.205 -69.875 -18.875 ;
        RECT -70.205 -20.565 -69.875 -20.235 ;
        RECT -70.205 -21.925 -69.875 -21.595 ;
        RECT -70.205 -23.285 -69.875 -22.955 ;
        RECT -70.205 -24.645 -69.875 -24.315 ;
        RECT -70.205 -26.005 -69.875 -25.675 ;
        RECT -70.205 -27.365 -69.875 -27.035 ;
        RECT -70.205 -28.725 -69.875 -28.395 ;
        RECT -70.205 -30.085 -69.875 -29.755 ;
        RECT -70.205 -31.445 -69.875 -31.115 ;
        RECT -70.205 -32.805 -69.875 -32.475 ;
        RECT -70.205 -34.165 -69.875 -33.835 ;
        RECT -70.205 -35.525 -69.875 -35.195 ;
        RECT -70.205 -36.885 -69.875 -36.555 ;
        RECT -70.205 -38.245 -69.875 -37.915 ;
        RECT -70.205 -39.605 -69.875 -39.275 ;
        RECT -70.205 -40.965 -69.875 -40.635 ;
        RECT -70.205 -42.325 -69.875 -41.995 ;
        RECT -70.205 -43.685 -69.875 -43.355 ;
        RECT -70.205 -45.045 -69.875 -44.715 ;
        RECT -70.205 -46.405 -69.875 -46.075 ;
        RECT -70.205 -47.765 -69.875 -47.435 ;
        RECT -70.205 -49.125 -69.875 -48.795 ;
        RECT -70.205 -50.485 -69.875 -50.155 ;
        RECT -70.205 -51.845 -69.875 -51.515 ;
        RECT -70.205 -53.205 -69.875 -52.875 ;
        RECT -70.205 -54.565 -69.875 -54.235 ;
        RECT -70.205 -55.925 -69.875 -55.595 ;
        RECT -70.205 -57.285 -69.875 -56.955 ;
        RECT -70.205 -58.645 -69.875 -58.315 ;
        RECT -70.205 -60.005 -69.875 -59.675 ;
        RECT -70.205 -61.365 -69.875 -61.035 ;
        RECT -70.205 -62.725 -69.875 -62.395 ;
        RECT -70.205 -64.085 -69.875 -63.755 ;
    END
  END vss
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -21.24 -224.365 -20.92 -224.045 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -28.04 -224.365 -27.72 -224.045 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -34.16 -224.365 -33.84 -224.045 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -40.28 -224.365 -39.96 -224.045 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -46.4 -224.365 -46.08 -224.045 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -52.52 -224.365 -52.2 -224.045 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -58.64 -224.365 -58.32 -224.045 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -64.76 -224.365 -64.44 -224.045 ;
    END
  END addr[7]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -9.68 -224.365 -9.36 -224.045 ;
    END
  END clk
  PIN din[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 5.6 -224.365 6 -223.965 ;
    END
  END din[0]
  PIN din[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 66.6 -224.365 67 -223.965 ;
    END
  END din[10]
  PIN din[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 72.7 -224.365 73.1 -223.965 ;
    END
  END din[11]
  PIN din[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 78.8 -224.365 79.2 -223.965 ;
    END
  END din[12]
  PIN din[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 84.9 -224.365 85.3 -223.965 ;
    END
  END din[13]
  PIN din[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91 -224.365 91.4 -223.965 ;
    END
  END din[14]
  PIN din[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 97.1 -224.365 97.5 -223.965 ;
    END
  END din[15]
  PIN din[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.2 -224.365 103.6 -223.965 ;
    END
  END din[16]
  PIN din[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.3 -224.365 109.7 -223.965 ;
    END
  END din[17]
  PIN din[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 115.4 -224.365 115.8 -223.965 ;
    END
  END din[18]
  PIN din[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.5 -224.365 121.9 -223.965 ;
    END
  END din[19]
  PIN din[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 11.7 -224.365 12.1 -223.965 ;
    END
  END din[1]
  PIN din[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 127.6 -224.365 128 -223.965 ;
    END
  END din[20]
  PIN din[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.7 -224.365 134.1 -223.965 ;
    END
  END din[21]
  PIN din[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 139.8 -224.365 140.2 -223.965 ;
    END
  END din[22]
  PIN din[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 145.9 -224.365 146.3 -223.965 ;
    END
  END din[23]
  PIN din[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 152 -224.365 152.4 -223.965 ;
    END
  END din[24]
  PIN din[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 158.1 -224.365 158.5 -223.965 ;
    END
  END din[25]
  PIN din[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 164.2 -224.365 164.6 -223.965 ;
    END
  END din[26]
  PIN din[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 170.3 -224.365 170.7 -223.965 ;
    END
  END din[27]
  PIN din[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.4 -224.365 176.8 -223.965 ;
    END
  END din[28]
  PIN din[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 182.5 -224.365 182.9 -223.965 ;
    END
  END din[29]
  PIN din[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 17.8 -224.365 18.2 -223.965 ;
    END
  END din[2]
  PIN din[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 188.6 -224.365 189 -223.965 ;
    END
  END din[30]
  PIN din[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 194.7 -224.365 195.1 -223.965 ;
    END
  END din[31]
  PIN din[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 23.9 -224.365 24.3 -223.965 ;
    END
  END din[3]
  PIN din[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 30 -224.365 30.4 -223.965 ;
    END
  END din[4]
  PIN din[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.1 -224.365 36.5 -223.965 ;
    END
  END din[5]
  PIN din[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 42.2 -224.365 42.6 -223.965 ;
    END
  END din[6]
  PIN din[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 48.3 -224.365 48.7 -223.965 ;
    END
  END din[7]
  PIN din[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 54.4 -224.365 54.8 -223.965 ;
    END
  END din[8]
  PIN din[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 60.5 -224.365 60.9 -223.965 ;
    END
  END din[9]
  PIN dout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 4 -224.365 4.4 -223.965 ;
    END
  END dout[0]
  PIN dout[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 65 -224.365 65.4 -223.965 ;
    END
  END dout[10]
  PIN dout[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.1 -224.365 71.5 -223.965 ;
    END
  END dout[11]
  PIN dout[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 77.2 -224.365 77.6 -223.965 ;
    END
  END dout[12]
  PIN dout[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.3 -224.365 83.7 -223.965 ;
    END
  END dout[13]
  PIN dout[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 89.4 -224.365 89.8 -223.965 ;
    END
  END dout[14]
  PIN dout[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 95.5 -224.365 95.9 -223.965 ;
    END
  END dout[15]
  PIN dout[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.6 -224.365 102 -223.965 ;
    END
  END dout[16]
  PIN dout[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 107.7 -224.365 108.1 -223.965 ;
    END
  END dout[17]
  PIN dout[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 113.8 -224.365 114.2 -223.965 ;
    END
  END dout[18]
  PIN dout[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.9 -224.365 120.3 -223.965 ;
    END
  END dout[19]
  PIN dout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 10.1 -224.365 10.5 -223.965 ;
    END
  END dout[1]
  PIN dout[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126 -224.365 126.4 -223.965 ;
    END
  END dout[20]
  PIN dout[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 132.1 -224.365 132.5 -223.965 ;
    END
  END dout[21]
  PIN dout[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.2 -224.365 138.6 -223.965 ;
    END
  END dout[22]
  PIN dout[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 144.3 -224.365 144.7 -223.965 ;
    END
  END dout[23]
  PIN dout[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 150.4 -224.365 150.8 -223.965 ;
    END
  END dout[24]
  PIN dout[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.5 -224.365 156.9 -223.965 ;
    END
  END dout[25]
  PIN dout[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 162.6 -224.365 163 -223.965 ;
    END
  END dout[26]
  PIN dout[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 168.7 -224.365 169.1 -223.965 ;
    END
  END dout[27]
  PIN dout[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 174.8 -224.365 175.2 -223.965 ;
    END
  END dout[28]
  PIN dout[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 180.9 -224.365 181.3 -223.965 ;
    END
  END dout[29]
  PIN dout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 16.2 -224.365 16.6 -223.965 ;
    END
  END dout[2]
  PIN dout[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 187 -224.365 187.4 -223.965 ;
    END
  END dout[30]
  PIN dout[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 193.1 -224.365 193.5 -223.965 ;
    END
  END dout[31]
  PIN dout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.3 -224.365 22.7 -223.965 ;
    END
  END dout[3]
  PIN dout[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.4 -224.365 28.8 -223.965 ;
    END
  END dout[4]
  PIN dout[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 34.5 -224.365 34.9 -223.965 ;
    END
  END dout[5]
  PIN dout[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 40.6 -224.365 41 -223.965 ;
    END
  END dout[6]
  PIN dout[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.7 -224.365 47.1 -223.965 ;
    END
  END dout[7]
  PIN dout[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 52.8 -224.365 53.2 -223.965 ;
    END
  END dout[8]
  PIN dout[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 58.9 -224.365 59.3 -223.965 ;
    END
  END dout[9]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -15.12 -224.365 -14.8 -224.045 ;
    END
  END we
  PIN wmask[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 6.4 -224.365 6.8 -223.965 ;
    END
  END wmask[0]
  PIN wmask[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 55.2 -224.365 55.6 -223.965 ;
    END
  END wmask[1]
  PIN wmask[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 104 -224.365 104.4 -223.965 ;
    END
  END wmask[2]
  PIN wmask[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 152.8 -224.365 153.2 -223.965 ;
    END
  END wmask[3]
  OBS
    LAYER met1 SPACING 0.14 ;
      RECT -76.825 -224.365 215.545 133.925 ;
    LAYER met2 SPACING 0.14 ;
      RECT -76.825 -224.365 215.545 133.925 ;
    LAYER met3 SPACING 0.3 ;
      RECT 1.195 -60.685 1.525 -60.355 ;
      RECT 1.2 -62.045 1.52 -60.355 ;
      RECT 1.195 -62.045 1.525 -61.715 ;
      RECT 0.515 -22.605 0.845 -22.275 ;
      RECT 0.52 -64.085 0.84 -22.275 ;
      RECT 0.515 -64.085 0.845 -63.755 ;
      RECT -0.165 -21.245 0.165 -20.915 ;
      RECT -0.16 -64.765 0.16 -20.915 ;
      RECT -0.165 -64.765 0.165 -64.435 ;
      RECT -9.005 -10.365 -8.675 -10.035 ;
      RECT -9 -141.605 -8.68 -10.035 ;
      RECT -9.005 -11.045 -8.675 -10.715 ;
      RECT -9.005 -141.605 -8.675 -141.275 ;
      RECT -9.685 -204.845 -9.355 -204.515 ;
      RECT -9.68 -223.555 -9.36 -204.515 ;
      RECT -9.685 -209.605 -9.355 -209.275 ;
      RECT -10.365 -205.525 -10.035 -205.195 ;
      RECT -10.36 -210.285 -10.04 -205.195 ;
      RECT -10.365 -210.285 -10.035 -209.955 ;
      RECT -12.405 -113.725 -12.075 -113.395 ;
      RECT -12.4 -196.685 -12.08 -113.395 ;
      RECT -12.405 -196.685 -12.075 -196.355 ;
      RECT -13.765 -67.485 -13.435 -67.155 ;
      RECT -13.76 -141.605 -13.44 -67.155 ;
      RECT -13.765 -141.605 -13.435 -141.275 ;
      RECT -14.445 -130.09 -14.115 -129.76 ;
      RECT -14.44 -208.925 -14.12 -129.76 ;
      RECT -14.445 -208.925 -14.115 -208.595 ;
      RECT -15.12 -223.555 -14.8 -210.51 ;
      RECT -15.125 -210.9 -14.795 -210.57 ;
      RECT -15.125 -130.57 -14.795 -130.24 ;
      RECT -15.12 -209.605 -14.8 -130.24 ;
      RECT -15.125 -209.605 -14.795 -209.275 ;
      RECT -15.805 -131.05 -15.475 -130.72 ;
      RECT -15.8 -208.245 -15.48 -130.72 ;
      RECT -15.805 -208.245 -15.475 -207.915 ;
      RECT -16.485 -208.245 -16.155 -207.915 ;
      RECT -16.48 -210.285 -16.16 -207.915 ;
      RECT -16.485 -210.285 -16.155 -209.955 ;
      RECT -16.485 -131.53 -16.155 -131.2 ;
      RECT -16.48 -207.565 -16.16 -131.2 ;
      RECT -16.485 -207.565 -16.155 -207.235 ;
      RECT -17.165 -207.565 -16.835 -207.235 ;
      RECT -17.16 -211.645 -16.84 -207.235 ;
      RECT -17.165 -211.645 -16.835 -211.315 ;
      RECT -18.525 -39.33 -18.195 -39 ;
      RECT -18.52 -108.285 -18.2 -39 ;
      RECT -18.525 -108.285 -18.195 -107.955 ;
      RECT -18.525 -18.15 -18.195 -17.82 ;
      RECT -18.52 -38.245 -18.2 -17.82 ;
      RECT -18.525 -38.245 -18.195 -37.915 ;
      RECT -19.205 -209.605 -18.875 -209.275 ;
      RECT -19.2 -211.645 -18.88 -209.275 ;
      RECT -19.205 -211.645 -18.875 -211.315 ;
      RECT -19.205 -39.81 -18.875 -39.48 ;
      RECT -19.2 -107.605 -18.88 -39.48 ;
      RECT -19.205 -107.605 -18.875 -107.275 ;
      RECT -19.205 -18.63 -18.875 -18.3 ;
      RECT -19.2 -36.205 -18.88 -18.3 ;
      RECT -19.205 -36.205 -18.875 -35.875 ;
      RECT -19.885 -204.845 -19.555 -204.515 ;
      RECT -19.88 -209.605 -19.56 -204.515 ;
      RECT -19.885 -209.605 -19.555 -209.275 ;
      RECT -19.885 -40.29 -19.555 -39.96 ;
      RECT -19.88 -106.925 -19.56 -39.96 ;
      RECT -19.885 -106.925 -19.555 -106.595 ;
      RECT -19.885 -19.11 -19.555 -18.78 ;
      RECT -19.88 -34.165 -19.56 -18.78 ;
      RECT -19.885 -34.165 -19.555 -33.835 ;
      RECT -20.565 -40.77 -20.235 -40.44 ;
      RECT -20.56 -104.885 -20.24 -40.44 ;
      RECT -20.565 -104.885 -20.235 -104.555 ;
      RECT -20.565 -19.59 -20.235 -19.26 ;
      RECT -20.56 -33.485 -20.24 -19.26 ;
      RECT -20.565 -33.485 -20.235 -33.155 ;
      RECT -21.24 -223.555 -20.92 -210.51 ;
      RECT -21.245 -210.9 -20.915 -210.57 ;
      RECT -21.245 -41.25 -20.915 -40.92 ;
      RECT -21.24 -106.245 -20.92 -40.92 ;
      RECT -21.245 -106.245 -20.915 -105.915 ;
      RECT -21.245 -20.07 -20.915 -19.74 ;
      RECT -21.24 -31.445 -20.92 -19.74 ;
      RECT -21.245 -31.445 -20.915 -31.115 ;
      RECT -21.925 -41.73 -21.595 -41.4 ;
      RECT -21.92 -105.565 -21.6 -41.4 ;
      RECT -21.925 -105.565 -21.595 -105.235 ;
      RECT -21.925 -20.55 -21.595 -20.22 ;
      RECT -21.92 -30.765 -21.6 -20.22 ;
      RECT -21.925 -30.765 -21.595 -30.435 ;
      RECT -23.285 -208.925 -22.955 -208.595 ;
      RECT -23.28 -210.285 -22.96 -208.595 ;
      RECT -23.285 -210.285 -22.955 -209.955 ;
      RECT -28.04 -223.555 -27.72 -210.51 ;
      RECT -28.045 -210.9 -27.715 -210.57 ;
      RECT -29.405 -132.765 -29.075 -132.435 ;
      RECT -29.4 -211.645 -29.08 -132.435 ;
      RECT -29.405 -211.645 -29.075 -211.315 ;
      RECT -30.085 -132.765 -29.755 -132.435 ;
      RECT -30.08 -210.285 -29.76 -132.435 ;
      RECT -30.085 -210.285 -29.755 -209.955 ;
      RECT -34.16 -223.555 -33.84 -210.51 ;
      RECT -34.165 -210.9 -33.835 -210.57 ;
      RECT -34.845 -133.445 -34.515 -133.115 ;
      RECT -34.84 -211.645 -34.52 -133.115 ;
      RECT -34.845 -211.645 -34.515 -211.315 ;
      RECT -35.525 -132.765 -35.195 -132.435 ;
      RECT -35.52 -210.285 -35.2 -132.435 ;
      RECT -35.525 -210.285 -35.195 -209.955 ;
      RECT -38.925 -132.765 -38.595 -132.435 ;
      RECT -38.92 -211.645 -38.6 -132.435 ;
      RECT -38.925 -211.645 -38.595 -211.315 ;
      RECT -40.28 -223.555 -39.96 -210.51 ;
      RECT -40.285 -210.9 -39.955 -210.57 ;
      RECT -41.645 -132.765 -41.315 -132.435 ;
      RECT -41.64 -210.285 -41.32 -132.435 ;
      RECT -41.645 -210.285 -41.315 -209.955 ;
      RECT -46 60.84 -44.72 61.43 ;
      RECT -45.04 -138.885 -44.72 61.43 ;
      RECT -45.045 -138.885 -44.715 -138.555 ;
      RECT -46.4 -223.555 -46.08 -210.51 ;
      RECT -46.405 -210.9 -46.075 -210.57 ;
      RECT -47.085 -132.765 -46.755 -132.435 ;
      RECT -47.08 -210.285 -46.76 -132.435 ;
      RECT -47.085 -210.285 -46.755 -209.955 ;
      RECT -48.445 -133.445 -48.115 -133.115 ;
      RECT -48.44 -211.645 -48.12 -133.115 ;
      RECT -48.445 -211.645 -48.115 -211.315 ;
      RECT -51.845 37.915 -51.515 38.245 ;
      RECT -51.84 -10.365 -51.52 38.245 ;
      RECT -51.845 -10.365 -51.515 -10.035 ;
      RECT -52.52 -223.555 -52.2 -210.51 ;
      RECT -52.525 -210.9 -52.195 -210.57 ;
      RECT -52.525 37.235 -52.195 37.565 ;
      RECT -52.52 -141.605 -52.2 37.565 ;
      RECT -52.525 -141.605 -52.195 -141.275 ;
      RECT -53.205 -132.765 -52.875 -132.435 ;
      RECT -53.2 -210.285 -52.88 -132.435 ;
      RECT -53.205 -210.285 -52.875 -209.955 ;
      RECT -54.565 -134.125 -54.235 -133.795 ;
      RECT -54.56 -211.645 -54.24 -133.795 ;
      RECT -54.565 -211.645 -54.235 -211.315 ;
      RECT -56.605 -132.085 -56.275 -131.755 ;
      RECT -56.6 -140.925 -56.28 -131.755 ;
      RECT -56.605 -140.925 -56.275 -140.595 ;
      RECT -58.64 -223.555 -58.32 -210.51 ;
      RECT -58.645 -210.9 -58.315 -210.57 ;
      RECT -60.005 -132.765 -59.675 -132.435 ;
      RECT -60 -210.285 -59.68 -132.435 ;
      RECT -60.005 -210.285 -59.675 -209.955 ;
      RECT -60.685 -133.445 -60.355 -133.115 ;
      RECT -60.68 -211.645 -60.36 -133.115 ;
      RECT -60.685 -211.645 -60.355 -211.315 ;
      RECT -64.76 -223.555 -64.44 -210.51 ;
      RECT -64.765 -210.9 -64.435 -210.57 ;
      RECT 196.3 -107.675 196.7 -22.12 ;
      RECT 195.5 -106.815 195.9 -22.12 ;
      RECT 194.7 -223.475 195.1 -106.905 ;
      RECT 193.9 -90.96 194.3 -76.365 ;
      RECT 193.9 -72.54 194.3 -17.24 ;
      RECT 193.1 -223.475 193.5 -101.065 ;
      RECT 193.1 -91.46 193.5 -76.82 ;
      RECT 193.1 -72.97 193.5 -12.97 ;
      RECT 190.2 -107.675 190.6 -22.12 ;
      RECT 189.4 -106.815 189.8 -22.12 ;
      RECT 188.6 -223.475 189 -106.905 ;
      RECT 187.8 -90.96 188.2 -76.365 ;
      RECT 187.8 -72.54 188.2 -17.24 ;
      RECT 187 -223.475 187.4 -101.065 ;
      RECT 187 -91.46 187.4 -76.82 ;
      RECT 187 -72.97 187.4 -12.97 ;
      RECT 184.1 -107.675 184.5 -22.12 ;
      RECT 183.3 -106.815 183.7 -22.12 ;
      RECT 182.5 -223.475 182.9 -106.905 ;
      RECT 181.7 -90.96 182.1 -76.365 ;
      RECT 181.7 -72.54 182.1 -17.24 ;
      RECT 180.9 -223.475 181.3 -101.065 ;
      RECT 180.9 -91.46 181.3 -76.82 ;
      RECT 180.9 -72.97 181.3 -12.97 ;
      RECT 178 -107.675 178.4 -22.12 ;
      RECT 177.2 -106.815 177.6 -22.12 ;
      RECT 176.4 -223.475 176.8 -106.905 ;
      RECT 175.6 -90.96 176 -76.365 ;
      RECT 175.6 -72.54 176 -17.24 ;
      RECT 174.8 -223.475 175.2 -101.065 ;
      RECT 174.8 -91.46 175.2 -76.82 ;
      RECT 174.8 -72.97 175.2 -12.97 ;
      RECT 171.9 -107.675 172.3 -22.12 ;
      RECT 171.1 -106.815 171.5 -22.12 ;
      RECT 170.3 -223.475 170.7 -106.905 ;
      RECT 169.5 -90.96 169.9 -76.365 ;
      RECT 169.5 -72.54 169.9 -17.24 ;
      RECT 168.7 -223.475 169.1 -101.065 ;
      RECT 168.7 -91.46 169.1 -76.82 ;
      RECT 168.7 -72.97 169.1 -12.97 ;
      RECT 165.8 -107.675 166.2 -22.12 ;
      RECT 165 -106.815 165.4 -22.12 ;
      RECT 164.2 -223.475 164.6 -106.905 ;
      RECT 163.4 -90.96 163.8 -76.365 ;
      RECT 163.4 -72.54 163.8 -17.24 ;
      RECT 162.6 -223.475 163 -101.065 ;
      RECT 162.6 -91.46 163 -76.82 ;
      RECT 162.6 -72.97 163 -12.97 ;
      RECT 159.7 -107.675 160.1 -22.12 ;
      RECT 158.9 -106.815 159.3 -22.12 ;
      RECT 158.1 -223.475 158.5 -106.905 ;
      RECT 157.3 -90.96 157.7 -76.365 ;
      RECT 157.3 -72.54 157.7 -17.24 ;
      RECT 156.5 -223.475 156.9 -101.065 ;
      RECT 156.5 -91.46 156.9 -76.82 ;
      RECT 156.5 -72.97 156.9 -12.97 ;
      RECT 154.4 -114.52 154.8 -22.12 ;
      RECT 153.6 -107.675 154 -22.12 ;
      RECT 152.8 -223.475 153.2 -114.61 ;
      RECT 152.8 -106.815 153.2 -22.12 ;
      RECT 152 -223.475 152.4 -106.905 ;
      RECT 151.2 -90.96 151.6 -76.365 ;
      RECT 151.2 -72.54 151.6 -17.24 ;
      RECT 150.4 -223.475 150.8 -101.065 ;
      RECT 150.4 -91.46 150.8 -76.82 ;
      RECT 150.4 -72.97 150.8 -12.97 ;
      RECT 147.5 -107.675 147.9 -22.12 ;
      RECT 146.7 -106.815 147.1 -22.12 ;
      RECT 145.9 -223.475 146.3 -106.905 ;
      RECT 145.1 -90.96 145.5 -76.365 ;
      RECT 145.1 -72.54 145.5 -17.24 ;
      RECT 144.3 -223.475 144.7 -101.065 ;
      RECT 144.3 -91.46 144.7 -76.82 ;
      RECT 144.3 -72.97 144.7 -12.97 ;
      RECT 141.4 -107.675 141.8 -22.12 ;
      RECT 140.6 -106.815 141 -22.12 ;
      RECT 139.8 -223.475 140.2 -106.905 ;
      RECT 139 -90.96 139.4 -76.365 ;
      RECT 139 -72.54 139.4 -17.24 ;
      RECT 138.2 -223.475 138.6 -101.065 ;
      RECT 138.2 -91.46 138.6 -76.82 ;
      RECT 138.2 -72.97 138.6 -12.97 ;
      RECT 135.3 -107.675 135.7 -22.12 ;
      RECT 134.5 -106.815 134.9 -22.12 ;
      RECT 133.7 -223.475 134.1 -106.905 ;
      RECT 132.9 -90.96 133.3 -76.365 ;
      RECT 132.9 -72.54 133.3 -17.24 ;
      RECT 132.1 -223.475 132.5 -101.065 ;
      RECT 132.1 -91.46 132.5 -76.82 ;
      RECT 132.1 -72.97 132.5 -12.97 ;
      RECT 129.2 -107.675 129.6 -22.12 ;
      RECT 128.4 -106.815 128.8 -22.12 ;
      RECT 127.6 -223.475 128 -106.905 ;
      RECT 126.8 -90.96 127.2 -76.365 ;
      RECT 126.8 -72.54 127.2 -17.24 ;
      RECT 126 -223.475 126.4 -101.065 ;
      RECT 126 -91.46 126.4 -76.82 ;
      RECT 126 -72.97 126.4 -12.97 ;
      RECT 123.1 -107.675 123.5 -22.12 ;
      RECT 122.3 -106.815 122.7 -22.12 ;
      RECT 121.5 -223.475 121.9 -106.905 ;
      RECT 120.7 -90.96 121.1 -76.365 ;
      RECT 120.7 -72.54 121.1 -17.24 ;
      RECT 119.9 -223.475 120.3 -101.065 ;
      RECT 119.9 -91.46 120.3 -76.82 ;
      RECT 119.9 -72.97 120.3 -12.97 ;
      RECT 117 -107.675 117.4 -22.12 ;
      RECT 116.2 -106.815 116.6 -22.12 ;
      RECT 115.4 -223.475 115.8 -106.905 ;
      RECT 114.6 -90.96 115 -76.365 ;
      RECT 114.6 -72.54 115 -17.24 ;
      RECT 113.8 -223.475 114.2 -101.065 ;
      RECT 113.8 -91.46 114.2 -76.82 ;
      RECT 113.8 -72.97 114.2 -12.97 ;
      RECT 110.9 -107.675 111.3 -22.12 ;
      RECT 110.1 -106.815 110.5 -22.12 ;
      RECT 109.3 -223.475 109.7 -106.905 ;
      RECT 108.5 -90.96 108.9 -76.365 ;
      RECT 108.5 -72.54 108.9 -17.24 ;
      RECT 107.7 -223.475 108.1 -101.065 ;
      RECT 107.7 -91.46 108.1 -76.82 ;
      RECT 107.7 -72.97 108.1 -12.97 ;
      RECT 105.6 -114.52 106 -22.12 ;
      RECT 104.8 -107.675 105.2 -22.12 ;
      RECT 104 -223.475 104.4 -114.61 ;
      RECT 104 -106.815 104.4 -22.12 ;
      RECT 103.2 -223.475 103.6 -106.905 ;
      RECT 102.4 -90.96 102.8 -76.365 ;
      RECT 102.4 -72.54 102.8 -17.24 ;
      RECT 101.6 -223.475 102 -101.065 ;
      RECT 101.6 -91.46 102 -76.82 ;
      RECT 101.6 -72.97 102 -12.97 ;
      RECT 98.7 -107.675 99.1 -22.12 ;
      RECT 97.9 -106.815 98.3 -22.12 ;
      RECT 97.1 -223.475 97.5 -106.905 ;
      RECT 96.3 -90.96 96.7 -76.365 ;
      RECT 96.3 -72.54 96.7 -17.24 ;
      RECT 95.5 -223.475 95.9 -101.065 ;
      RECT 95.5 -91.46 95.9 -76.82 ;
      RECT 95.5 -72.97 95.9 -12.97 ;
      RECT 92.6 -107.675 93 -22.12 ;
      RECT 91.8 -106.815 92.2 -22.12 ;
      RECT 91 -223.475 91.4 -106.905 ;
      RECT 90.2 -90.96 90.6 -76.365 ;
      RECT 90.2 -72.54 90.6 -17.24 ;
      RECT 89.4 -223.475 89.8 -101.065 ;
      RECT 89.4 -91.46 89.8 -76.82 ;
      RECT 89.4 -72.97 89.8 -12.97 ;
      RECT 86.5 -107.675 86.9 -22.12 ;
      RECT 85.7 -106.815 86.1 -22.12 ;
      RECT 84.9 -223.475 85.3 -106.905 ;
      RECT 84.1 -90.96 84.5 -76.365 ;
      RECT 84.1 -72.54 84.5 -17.24 ;
      RECT 83.3 -223.475 83.7 -101.065 ;
      RECT 83.3 -91.46 83.7 -76.82 ;
      RECT 83.3 -72.97 83.7 -12.97 ;
      RECT 80.4 -107.675 80.8 -22.12 ;
      RECT 79.6 -106.815 80 -22.12 ;
      RECT 78.8 -223.475 79.2 -106.905 ;
      RECT 78 -90.96 78.4 -76.365 ;
      RECT 78 -72.54 78.4 -17.24 ;
      RECT 77.2 -223.475 77.6 -101.065 ;
      RECT 77.2 -91.46 77.6 -76.82 ;
      RECT 77.2 -72.97 77.6 -12.97 ;
      RECT 74.3 -107.675 74.7 -22.12 ;
      RECT 73.5 -106.815 73.9 -22.12 ;
      RECT 72.7 -223.475 73.1 -106.905 ;
      RECT 71.9 -90.96 72.3 -76.365 ;
      RECT 71.9 -72.54 72.3 -17.24 ;
      RECT 71.1 -223.475 71.5 -101.065 ;
      RECT 71.1 -91.46 71.5 -76.82 ;
      RECT 71.1 -72.97 71.5 -12.97 ;
      RECT 68.2 -107.675 68.6 -22.12 ;
      RECT 67.4 -106.815 67.8 -22.12 ;
      RECT 66.6 -223.475 67 -106.905 ;
      RECT 65.8 -90.96 66.2 -76.365 ;
      RECT 65.8 -72.54 66.2 -17.24 ;
      RECT 65 -223.475 65.4 -101.065 ;
      RECT 65 -91.46 65.4 -76.82 ;
      RECT 65 -72.97 65.4 -12.97 ;
      RECT 62.1 -107.675 62.5 -22.12 ;
      RECT 61.3 -106.815 61.7 -22.12 ;
      RECT 60.5 -223.475 60.9 -106.905 ;
      RECT 59.7 -90.96 60.1 -76.365 ;
      RECT 59.7 -72.54 60.1 -17.24 ;
      RECT 58.9 -223.475 59.3 -101.065 ;
      RECT 58.9 -91.46 59.3 -76.82 ;
      RECT 58.9 -72.97 59.3 -12.97 ;
      RECT 56.8 -114.52 57.2 -22.12 ;
      RECT 56 -107.675 56.4 -22.12 ;
      RECT 55.2 -223.475 55.6 -114.61 ;
      RECT 55.2 -106.815 55.6 -22.12 ;
      RECT 54.4 -223.475 54.8 -106.905 ;
      RECT 53.6 -90.96 54 -76.365 ;
      RECT 53.6 -72.54 54 -17.24 ;
      RECT 52.8 -223.475 53.2 -101.065 ;
      RECT 52.8 -91.46 53.2 -76.82 ;
      RECT 52.8 -72.97 53.2 -12.97 ;
      RECT 49.9 -107.675 50.3 -22.12 ;
      RECT 49.1 -106.815 49.5 -22.12 ;
      RECT 48.3 -223.475 48.7 -106.905 ;
      RECT 47.5 -90.96 47.9 -76.365 ;
      RECT 47.5 -72.54 47.9 -17.24 ;
      RECT 46.7 -223.475 47.1 -101.065 ;
      RECT 46.7 -91.46 47.1 -76.82 ;
      RECT 46.7 -72.97 47.1 -12.97 ;
      RECT 43.8 -107.675 44.2 -22.12 ;
      RECT 43 -106.815 43.4 -22.12 ;
      RECT 42.2 -223.475 42.6 -106.905 ;
      RECT 41.4 -90.96 41.8 -76.365 ;
      RECT 41.4 -72.54 41.8 -17.24 ;
      RECT 40.6 -223.475 41 -101.065 ;
      RECT 40.6 -91.46 41 -76.82 ;
      RECT 40.6 -72.97 41 -12.97 ;
      RECT 37.7 -107.675 38.1 -22.12 ;
      RECT 36.9 -106.815 37.3 -22.12 ;
      RECT 36.1 -223.475 36.5 -106.905 ;
      RECT 35.3 -90.96 35.7 -76.365 ;
      RECT 35.3 -72.54 35.7 -17.24 ;
      RECT 34.5 -223.475 34.9 -101.065 ;
      RECT 34.5 -91.46 34.9 -76.82 ;
      RECT 34.5 -72.97 34.9 -12.97 ;
      RECT 31.6 -107.675 32 -22.12 ;
      RECT 30.8 -106.815 31.2 -22.12 ;
      RECT 30 -223.475 30.4 -106.905 ;
      RECT 29.2 -90.96 29.6 -76.365 ;
      RECT 29.2 -72.54 29.6 -17.24 ;
      RECT 28.4 -223.475 28.8 -101.065 ;
      RECT 28.4 -91.46 28.8 -76.82 ;
      RECT 28.4 -72.97 28.8 -12.97 ;
      RECT 25.5 -107.675 25.9 -22.12 ;
      RECT 24.7 -106.815 25.1 -22.12 ;
      RECT 23.9 -223.475 24.3 -106.905 ;
      RECT 23.1 -90.96 23.5 -76.365 ;
      RECT 23.1 -72.54 23.5 -17.24 ;
      RECT 22.3 -223.475 22.7 -101.065 ;
      RECT 22.3 -91.46 22.7 -76.82 ;
      RECT 22.3 -72.97 22.7 -12.97 ;
      RECT 19.4 -107.675 19.8 -22.12 ;
      RECT 18.6 -106.815 19 -22.12 ;
      RECT 17.8 -223.475 18.2 -106.905 ;
      RECT 17 -90.96 17.4 -76.365 ;
      RECT 17 -72.54 17.4 -17.24 ;
      RECT 16.2 -223.475 16.6 -101.065 ;
      RECT 16.2 -91.46 16.6 -76.82 ;
      RECT 16.2 -72.97 16.6 -12.97 ;
      RECT 13.3 -107.675 13.7 -22.12 ;
      RECT 12.5 -106.815 12.9 -22.12 ;
      RECT 11.7 -223.475 12.1 -106.905 ;
      RECT 10.9 -90.96 11.3 -76.365 ;
      RECT 10.9 -72.54 11.3 -17.24 ;
      RECT 10.1 -223.475 10.5 -101.065 ;
      RECT 10.1 -91.46 10.5 -76.82 ;
      RECT 10.1 -72.97 10.5 -12.97 ;
      RECT 8 -114.52 8.4 -22.12 ;
      RECT 7.2 -107.675 7.6 -22.12 ;
      RECT 6.4 -223.475 6.8 -114.61 ;
      RECT 6.4 -106.815 6.8 -22.12 ;
      RECT 5.6 -223.475 6 -106.905 ;
      RECT 4.8 -90.96 5.2 -76.365 ;
      RECT 4.8 -72.54 5.2 -17.24 ;
      RECT 4 -223.475 4.4 -101.065 ;
      RECT 4 -91.46 4.4 -76.82 ;
      RECT 4 -72.97 4.4 -12.97 ;
  END
END sram22_256x32m4w8

END LIBRARY
