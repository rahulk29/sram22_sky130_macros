* Substrate SPICE library
* This is a generated file. Be careful when editing manually: this file may be overwritten.


.SUBCKT mos_w700_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.700


.ENDS mos_w700_l150_m1_nf1_id1

.SUBCKT mos_w700_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.700


.ENDS mos_w700_l150_m1_nf1_id0

.SUBCKT multi_finger_inv_10 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_10

.SUBCKT mos_w7050_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=7.050


.ENDS mos_w7050_l150_m1_nf1_id1

.SUBCKT mos_w900_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.900


.ENDS mos_w900_l150_m1_nf1_id0

.SUBCKT multi_finger_inv_8 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP19 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP20 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP21 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP22 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP23 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP24 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP25 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP26 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP27 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP28 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP29 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP30 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP31 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN7 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN8 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN9 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN10 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN11 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN12 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_8

.SUBCKT mos_w1250_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.250


.ENDS mos_w1250_l150_m1_nf1_id1

.SUBCKT mos_w500_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.500


.ENDS mos_w500_l150_m1_nf1_id0

.SUBCKT folded_inv vdd vss a y

  XMP0 y a vdd vdd mos_w1250_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w500_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w1250_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w500_l150_m1_nf1_id0

.ENDS folded_inv

.SUBCKT multi_finger_inv_5 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_5

.SUBCKT decoder_stage_4 vdd vss y y_b predecode_0_0

  Xgate_0_0_0 vdd vss predecode_0_0 y_b folded_inv
  Xgate_1_0_0 vdd vss y_b y multi_finger_inv_5
  Xgate_1_0_1 vdd vss y_b y multi_finger_inv_5

.ENDS decoder_stage_4

.SUBCKT sram_sp_cell_replica BL BR VSS VDD VPB VNB WL

  X0 VDD WL BR VNB sky130_fd_pr__special_nfet_pass l=0.150 nf=1 w=0.140

  X1 Q VDD VSS VNB sky130_fd_pr__special_nfet_latch l=0.150 nf=1 w=0.210

  X2 BL WL Q VNB sky130_fd_pr__special_nfet_pass l=0.150 nf=1 w=0.140

  X3 Q WL Q VPB sky130_fd_pr__special_pfet_pass l=0.025 nf=1 w=0.140

  X4 VDD WL VDD VPB sky130_fd_pr__special_pfet_pass l=0.025 nf=1 w=0.140

  X5 VDD Q VDD VPB sky130_fd_pr__special_pfet_pass l=0.150 nf=1 w=0.140

  X6 Q VDD VDD VPB sky130_fd_pr__special_pfet_pass l=0.150 nf=1 w=0.140

  X7 VSS Q VDD VNB sky130_fd_pr__special_nfet_latch l=0.150 nf=1 w=0.210


.ENDS sram_sp_cell_replica

.SUBCKT sram_sp_cell_replica_wrapper BL BR VSS VDD VPB VNB WL

  X0 BL BR VSS VDD VPB VNB WL sram_sp_cell_replica

.ENDS sram_sp_cell_replica_wrapper

.SUBCKT multi_finger_inv vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv

.SUBCKT sky130_fd_sc_hs__dfrbp_2 CLK D RESET_B VGND VNB VPB VPWR Q Q_N

  X0 a_1800_291# a_1586_149# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X1 VGND CLK a_728_331# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X2 Q a_2363_352# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X3 VPWR CLK a_728_331# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X4 a_1499_149# a_728_331# a_1586_149# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X5 a_536_81# a_331_392# a_614_81# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X6 a_156_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X7 a_298_294# a_818_418# a_614_81# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X8 a_70_74# a_728_331# a_298_294# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X9 a_331_392# a_728_331# a_1586_149# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X10 a_70_74# D a_156_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X11 a_818_418# a_728_331# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X12 a_818_418# a_728_331# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X13 a_1586_149# a_818_418# a_1755_389# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X14 Q_N a_1586_149# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X15 a_298_294# a_818_418# a_70_74# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X16 VGND RESET_B a_536_81# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X17 a_1755_389# a_1800_291# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X18 a_1586_149# a_818_418# a_331_392# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X19 Q a_2363_352# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X20 VGND a_1586_149# Q_N VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X21 VGND a_1586_149# a_2363_352# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X22 VPWR a_298_294# a_331_392# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X23 a_298_294# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X24 a_1499_149# a_1800_291# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X25 VPWR a_331_392# a_683_485# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X26 VPWR D a_70_74# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X27 VPWR RESET_B a_1800_291# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X28 a_1974_74# a_1586_149# a_1800_291# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X29 a_70_74# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X30 Q_N a_1586_149# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X31 VPWR a_1586_149# a_2363_352# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X32 VGND a_2363_352# Q VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X33 VPWR a_1586_149# Q_N VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X34 VGND RESET_B a_1974_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X35 a_683_485# a_728_331# a_298_294# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X36 VGND a_298_294# a_331_392# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X37 VPWR a_2363_352# Q VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120


.ENDS sky130_fd_sc_hs__dfrbp_2

.SUBCKT sky130_fd_sc_hs__dfrbp_2_wrapper CLK D RESET_B VGND VNB VPB VPWR Q Q_N

  X0 CLK D RESET_B VGND VNB VPB VPWR Q Q_N sky130_fd_sc_hs__dfrbp_2

.ENDS sky130_fd_sc_hs__dfrbp_2_wrapper

.SUBCKT dff_array_12 vdd vss clk rb d[0] d[1] d[2] d[3] d[4] d[5] d[6] d[7] d[8] d[9] d[10] d[11] q[0] q[1] q[2] q[3] q[4] q[5] q[6] q[7] q[8] q[9] q[10] q[11] qn[0] qn[1] qn[2] qn[3] qn[4] qn[5] qn[6] qn[7] qn[8] qn[9] qn[10] qn[11]

  Xdff_0 clk d[0] rb vss vss vdd vdd q[0] qn[0] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_1 clk d[1] rb vss vss vdd vdd q[1] qn[1] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_2 clk d[2] rb vss vss vdd vdd q[2] qn[2] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_3 clk d[3] rb vss vss vdd vdd q[3] qn[3] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_4 clk d[4] rb vss vss vdd vdd q[4] qn[4] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_5 clk d[5] rb vss vss vdd vdd q[5] qn[5] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_6 clk d[6] rb vss vss vdd vdd q[6] qn[6] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_7 clk d[7] rb vss vss vdd vdd q[7] qn[7] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_8 clk d[8] rb vss vss vdd vdd q[8] qn[8] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_9 clk d[9] rb vss vss vdd vdd q[9] qn[9] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_10 clk d[10] rb vss vss vdd vdd q[10] qn[10] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_11 clk d[11] rb vss vss vdd vdd q[11] qn[11] sky130_fd_sc_hs__dfrbp_2_wrapper

.ENDS dff_array_12

.SUBCKT sky130_fd_sc_hs__buf_16 A VGND VNB VPB VPWR X

  X0 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X3 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X4 VPWR A a_83_260# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X5 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X6 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X7 VPWR A a_83_260# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X8 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X9 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 VPWR A a_83_260# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X11 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X12 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X13 a_83_260# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X14 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X15 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X16 VGND A a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X17 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X18 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X19 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X20 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X21 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X22 VGND A a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X23 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X24 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X25 a_83_260# A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X26 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X27 a_83_260# A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X28 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X29 a_83_260# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X30 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X31 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X32 a_83_260# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X33 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X34 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X35 a_83_260# A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X36 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X37 VGND A a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X38 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X39 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X40 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X41 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X42 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X43 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__buf_16

.SUBCKT sky130_fd_sc_hs__buf_16_wrapper A VGND VNB VPB VPWR X

  X0 A VGND VNB VPB VPWR X sky130_fd_sc_hs__buf_16

.ENDS sky130_fd_sc_hs__buf_16_wrapper

.SUBCKT sramgen_svt_inv_2 A VGND VNB VPB VPWR Y

  X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740

  X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740


.ENDS sramgen_svt_inv_2

.SUBCKT mos_w2000_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=2.000


.ENDS mos_w2000_l150_m1_nf1_id0

.SUBCKT mos_w2500_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.500


.ENDS mos_w2500_l150_m1_nf1_id1

.SUBCKT nand2_1 vdd vss a b y

  Xn1 x a vss vss mos_w2000_l150_m1_nf1_id0
  Xn2 y b x vss mos_w2000_l150_m1_nf1_id0
  Xp1 y a vdd vdd mos_w2500_l150_m1_nf1_id1
  Xp2 y b vdd vdd mos_w2500_l150_m1_nf1_id1

.ENDS nand2_1

.SUBCKT mos_w3200_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=3.200


.ENDS mos_w3200_l150_m1_nf1_id1

.SUBCKT mos_w1280_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.280


.ENDS mos_w1280_l150_m1_nf1_id0

.SUBCKT folded_inv_8 vdd vss a y

  XMP0 y a vdd vdd mos_w3200_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w1280_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w3200_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w1280_l150_m1_nf1_id0

.ENDS folded_inv_8

.SUBCKT decoder_stage_10 vdd vss y[0] y[1] y[2] y[3] y_b[0] y_b[1] y_b[2] y_b[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1

  Xgate_0_0_0 vdd vss predecode_0_0 predecode_1_0 y_b[0] nand2_1
  Xgate_0_1_0 vdd vss predecode_0_1 predecode_1_0 y_b[1] nand2_1
  Xgate_0_2_0 vdd vss predecode_0_0 predecode_1_1 y_b[2] nand2_1
  Xgate_0_3_0 vdd vss predecode_0_1 predecode_1_1 y_b[3] nand2_1
  Xgate_1_0_0 vdd vss y_b[0] y[0] folded_inv_8
  Xgate_1_1_0 vdd vss y_b[1] y[1] folded_inv_8
  Xgate_1_2_0 vdd vss y_b[2] y[2] folded_inv_8
  Xgate_1_3_0 vdd vss y_b[3] y[3] folded_inv_8

.ENDS decoder_stage_10

.SUBCKT multi_finger_inv_1 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_1

.SUBCKT multi_finger_inv_2 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_2

.SUBCKT decoder_stage_1 vdd vss y y_b predecode_0_0

  Xgate_0_0_0 vdd vss predecode_0_0 x_0 folded_inv
  Xgate_1_0_0 vdd vss x_0 x_1 multi_finger_inv
  Xgate_1_0_1 vdd vss x_0 x_1 multi_finger_inv
  Xgate_2_0_0 vdd vss x_1 y_b multi_finger_inv_1
  Xgate_2_0_1 vdd vss x_1 y_b multi_finger_inv_1
  Xgate_2_0_2 vdd vss x_1 y_b multi_finger_inv_1
  Xgate_2_0_3 vdd vss x_1 y_b multi_finger_inv_1
  Xgate_2_0_4 vdd vss x_1 y_b multi_finger_inv_1
  Xgate_2_0_5 vdd vss x_1 y_b multi_finger_inv_1
  Xgate_2_0_6 vdd vss x_1 y_b multi_finger_inv_1
  Xgate_3_0_0 vdd vss y_b y multi_finger_inv_2
  Xgate_3_0_1 vdd vss y_b y multi_finger_inv_2
  Xgate_3_0_2 vdd vss y_b y multi_finger_inv_2
  Xgate_3_0_3 vdd vss y_b y multi_finger_inv_2
  Xgate_3_0_4 vdd vss y_b y multi_finger_inv_2
  Xgate_3_0_5 vdd vss y_b y multi_finger_inv_2
  Xgate_3_0_6 vdd vss y_b y multi_finger_inv_2
  Xgate_3_0_7 vdd vss y_b y multi_finger_inv_2
  Xgate_3_0_8 vdd vss y_b y multi_finger_inv_2
  Xgate_3_0_9 vdd vss y_b y multi_finger_inv_2
  Xgate_3_0_10 vdd vss y_b y multi_finger_inv_2
  Xgate_3_0_11 vdd vss y_b y multi_finger_inv_2
  Xgate_3_0_12 vdd vss y_b y multi_finger_inv_2

.ENDS decoder_stage_1

.SUBCKT mos_w800_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.800


.ENDS mos_w800_l150_m1_nf1_id0

.SUBCKT mos_w1950_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.950


.ENDS mos_w1950_l150_m1_nf1_id0

.SUBCKT mos_w2850_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.850


.ENDS mos_w2850_l150_m1_nf1_id1

.SUBCKT column_mos vdd vss bl

  Xgate_nmos vss bl vss vss mos_w800_l150_m1_nf1_id0
  Xdrain_nmos bl vss vss vss mos_w1950_l150_m1_nf1_id0
  Xdrain_pmos bl vdd vdd vdd mos_w2850_l150_m1_nf1_id1

.ENDS column_mos

.SUBCKT mos_w3000_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=3.000


.ENDS mos_w3000_l150_m1_nf1_id0

.SUBCKT nand3 vdd vss a b c y

  Xn1 x1 a vss vss mos_w3000_l150_m1_nf1_id0
  Xn2 x2 b x1 vss mos_w3000_l150_m1_nf1_id0
  Xn3 y c x2 vss mos_w3000_l150_m1_nf1_id0
  Xp1 y a vdd vdd mos_w2500_l150_m1_nf1_id1
  Xp2 y b vdd vdd mos_w2500_l150_m1_nf1_id1
  Xp3 y c vdd vdd mos_w2500_l150_m1_nf1_id1

.ENDS nand3

.SUBCKT mos_w2690_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.690


.ENDS mos_w2690_l150_m1_nf1_id1

.SUBCKT mos_w1080_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.080


.ENDS mos_w1080_l150_m1_nf1_id0

.SUBCKT folded_inv_5 vdd vss a y

  XMP0 y a vdd vdd mos_w2690_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w1080_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w2690_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w1080_l150_m1_nf1_id0

.ENDS folded_inv_5

.SUBCKT decoder_stage_9 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 predecode_2_0 predecode_2_1

  Xgate_0_0_0 vdd vss predecode_0_0 predecode_1_0 predecode_2_0 y_b[0] nand3
  Xgate_0_1_0 vdd vss predecode_0_1 predecode_1_0 predecode_2_0 y_b[1] nand3
  Xgate_0_2_0 vdd vss predecode_0_0 predecode_1_1 predecode_2_0 y_b[2] nand3
  Xgate_0_3_0 vdd vss predecode_0_1 predecode_1_1 predecode_2_0 y_b[3] nand3
  Xgate_0_4_0 vdd vss predecode_0_0 predecode_1_0 predecode_2_1 y_b[4] nand3
  Xgate_0_5_0 vdd vss predecode_0_1 predecode_1_0 predecode_2_1 y_b[5] nand3
  Xgate_0_6_0 vdd vss predecode_0_0 predecode_1_1 predecode_2_1 y_b[6] nand3
  Xgate_0_7_0 vdd vss predecode_0_1 predecode_1_1 predecode_2_1 y_b[7] nand3
  Xgate_1_0_0 vdd vss y_b[0] y[0] folded_inv_5
  Xgate_1_0_1 vdd vss y_b[0] y[0] folded_inv_5
  Xgate_1_1_0 vdd vss y_b[1] y[1] folded_inv_5
  Xgate_1_1_1 vdd vss y_b[1] y[1] folded_inv_5
  Xgate_1_2_0 vdd vss y_b[2] y[2] folded_inv_5
  Xgate_1_2_1 vdd vss y_b[2] y[2] folded_inv_5
  Xgate_1_3_0 vdd vss y_b[3] y[3] folded_inv_5
  Xgate_1_3_1 vdd vss y_b[3] y[3] folded_inv_5
  Xgate_1_4_0 vdd vss y_b[4] y[4] folded_inv_5
  Xgate_1_4_1 vdd vss y_b[4] y[4] folded_inv_5
  Xgate_1_5_0 vdd vss y_b[5] y[5] folded_inv_5
  Xgate_1_5_1 vdd vss y_b[5] y[5] folded_inv_5
  Xgate_1_6_0 vdd vss y_b[6] y[6] folded_inv_5
  Xgate_1_6_1 vdd vss y_b[6] y[6] folded_inv_5
  Xgate_1_7_0 vdd vss y_b[7] y[7] folded_inv_5
  Xgate_1_7_1 vdd vss y_b[7] y[7] folded_inv_5

.ENDS decoder_stage_9

.SUBCKT mos_w2270_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.270


.ENDS mos_w2270_l150_m1_nf1_id1

.SUBCKT folded_inv_4 vdd vss a y

  XMP0 y a vdd vdd mos_w2270_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w900_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w2270_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w900_l150_m1_nf1_id0

.ENDS folded_inv_4

.SUBCKT sky130_fd_sc_hs__inv_2 A VGND VNB VPB VPWR Y

  X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X3 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__inv_2

.SUBCKT sky130_fd_sc_hs__inv_2_wrapper A VGND VNB VPB VPWR Y

  X0 A VGND VNB VPB VPWR Y sky130_fd_sc_hs__inv_2

.ENDS sky130_fd_sc_hs__inv_2_wrapper

.SUBCKT sky130_fd_sc_hs__inv_4 A VGND VNB VPB VPWR Y

  X0 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X4 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X7 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__inv_4

.SUBCKT sky130_fd_sc_hs__inv_4_wrapper A VGND VNB VPB VPWR Y

  X0 A VGND VNB VPB VPWR Y sky130_fd_sc_hs__inv_4

.ENDS sky130_fd_sc_hs__inv_4_wrapper

.SUBCKT inv_chain_3 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sky130_fd_sc_hs__inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_3

.SUBCKT mos_w5000_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=5.000


.ENDS mos_w5000_l150_m1_nf1_id1

.SUBCKT column_mos_1 vdd vss bl

  Xdrain_nmos bl vss vss vss mos_w1950_l150_m1_nf1_id0
  Xdrain_pmos bl vdd vdd vdd mos_w2850_l150_m1_nf1_id1

.ENDS column_mos_1

.SUBCKT column_mos_2 vdd vss bl

  Xdrain_nmos bl vss vss vss mos_w1950_l150_m1_nf1_id0

.ENDS column_mos_2

.SUBCKT replica_column_mos vdd vss bl

  Xunit0 vdd vss bl column_mos
  Xunit1 vdd vss bl column_mos_1
  Xunit2 vdd vss bl column_mos_1
  Xunit3 vdd vss bl column_mos_1
  Xunit4 vdd vss bl column_mos_2

.ENDS replica_column_mos

.SUBCKT mos_w600_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.600


.ENDS mos_w600_l150_m1_nf1_id0

.SUBCKT mos_w2100_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.100


.ENDS mos_w2100_l150_m1_nf1_id1

.SUBCKT mos_w850_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.850


.ENDS mos_w850_l150_m1_nf1_id0

.SUBCKT folded_inv_6 vdd vss a y

  XMP0 y a vdd vdd mos_w2100_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w850_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w2100_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w850_l150_m1_nf1_id0

.ENDS folded_inv_6

.SUBCKT sky130_fd_sc_hs__and2_4 A B VGND VNB VPB VPWR X

  X0 VPWR a_83_269# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 VPWR B a_83_269# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.840

  X2 VPWR a_83_269# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 a_504_119# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X4 a_83_269# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.840

  X5 VGND B a_504_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X6 VGND a_83_269# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X7 a_83_269# B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.840

  X8 X a_83_269# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 VGND a_83_269# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 X a_83_269# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X11 X a_83_269# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X12 a_504_119# A a_83_269# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X13 a_83_269# A a_504_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X14 VPWR A a_83_269# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.840

  X15 X a_83_269# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__and2_4

.SUBCKT sky130_fd_sc_hs__and2_4_wrapper A B VGND VNB VPB VPWR X

  X0 A B VGND VNB VPB VPWR X sky130_fd_sc_hs__and2_4

.ENDS sky130_fd_sc_hs__and2_4_wrapper

.SUBCKT sky130_fd_sc_hs__mux2_4 A0 A1 S VGND VNB VPB VPWR X

  X0 a_27_368# S VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X1 a_722_391# A0 a_193_241# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X2 a_722_391# S VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X3 VGND a_27_368# a_937_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X4 a_193_241# A1 a_936_391# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X5 a_709_119# S VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X6 a_709_119# A1 a_193_241# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X7 X a_193_241# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X8 X a_193_241# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 VPWR a_27_368# a_936_391# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X10 X a_193_241# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X11 a_193_241# A0 a_722_391# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X12 a_937_119# A0 a_193_241# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X13 a_936_391# a_27_368# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X14 VGND a_193_241# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X15 VPWR a_193_241# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X16 VPWR S a_722_391# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X17 a_936_391# A1 a_193_241# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X18 a_193_241# A0 a_937_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X19 a_193_241# A1 a_709_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X20 X a_193_241# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X21 VGND a_193_241# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X22 a_27_368# S VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X23 a_937_119# a_27_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X24 VPWR a_193_241# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X25 VGND S a_709_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640


.ENDS sky130_fd_sc_hs__mux2_4

.SUBCKT sky130_fd_sc_hs__mux2_4_wrapper A0 A1 S VGND VNB VPB VPWR X

  X0 A0 A1 S VGND VNB VPB VPWR X sky130_fd_sc_hs__mux2_4

.ENDS sky130_fd_sc_hs__mux2_4_wrapper

.SUBCKT mos_w2000_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.000


.ENDS mos_w2000_l150_m1_nf1_id1

.SUBCKT folded_inv_2 vdd vss a y

  XMP0 y a vdd vdd mos_w2000_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w800_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w2000_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w800_l150_m1_nf1_id0

.ENDS folded_inv_2

.SUBCKT mos_w4700_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=4.700


.ENDS mos_w4700_l150_m1_nf1_id0

.SUBCKT tgate_mux sel_b sel bl br bl_out br_out vdd vss

  XMPBL bl_out sel_b bl vdd mos_w7050_l150_m1_nf1_id1
  XMPBR br_out sel_b br vdd mos_w7050_l150_m1_nf1_id1
  XMNBL bl_out sel bl vss mos_w4700_l150_m1_nf1_id0
  XMNBR br_out sel br vss mos_w4700_l150_m1_nf1_id0

.ENDS tgate_mux

.SUBCKT multi_finger_inv_3 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_3

.SUBCKT sram_sp_colend BR VDD VSS BL VNB VPB

  X0 BR VNB BR VNB sky130_fd_pr__special_nfet_pass l=0.140 nf=1 w=0.140


.ENDS sram_sp_colend

.SUBCKT sram_sp_colend_wrapper BR VDD VSS BL VNB VPB

  X0 BR VDD VSS BL VNB VPB sram_sp_colend

.ENDS sram_sp_colend_wrapper

.SUBCKT nand2 vdd vss a b y

  Xn1 x a vss vss mos_w2000_l150_m1_nf1_id0
  Xn2 y b x vss mos_w2000_l150_m1_nf1_id0
  Xp1 y a vdd vdd mos_w2500_l150_m1_nf1_id1
  Xp2 y b vdd vdd mos_w2500_l150_m1_nf1_id1

.ENDS nand2

.SUBCKT and2_1 vdd a b y yb vss

  X0 vdd vss a b yb nand2
  X0_1 vdd vss yb y folded_inv_6

.ENDS and2_1

.SUBCKT sky130_fd_sc_hs__nand2_8 A B VGND VNB VPB VPWR Y

  X0 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X1 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X2 Y B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X4 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X5 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X6 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X7 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X11 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X12 VPWR B Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X13 VPWR B Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X14 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X16 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X17 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X18 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X19 Y B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X20 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X21 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X22 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X23 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120


.ENDS sky130_fd_sc_hs__nand2_8

.SUBCKT sky130_fd_sc_hs__nand2_8_wrapper A B VGND VNB VPB VPWR Y

  X0 A B VGND VNB VPB VPWR Y sky130_fd_sc_hs__nand2_8

.ENDS sky130_fd_sc_hs__nand2_8_wrapper

.SUBCKT sr_latch sb rb q qb vdd vss

  Xnand_set q0b sb vss vss vdd vdd q0 sky130_fd_sc_hs__nand2_8_wrapper
  Xnand_reset q0 rb vss vss vdd vdd q0b sky130_fd_sc_hs__nand2_8_wrapper
  Xqb_inv q0 vss vss vdd vdd qb sky130_fd_sc_hs__inv_2_wrapper
  Xq_inv q0b vss vss vdd vdd q sky130_fd_sc_hs__inv_2_wrapper

.ENDS sr_latch

.SUBCKT mos_w3000_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=3.000


.ENDS mos_w3000_l150_m1_nf1_id1

.SUBCKT precharge_1 vdd bl br en_b

  Xbl_pull_up bl en_b vdd vdd mos_w5000_l150_m1_nf1_id1
  Xbr_pull_up br en_b vdd vdd mos_w5000_l150_m1_nf1_id1
  Xequalizer bl en_b br vdd mos_w3000_l150_m1_nf1_id1

.ENDS precharge_1

.SUBCKT sram_sp_hstrap BR VDD VSS BL VNB VPB

  X0 BL VNB BL VNB sky130_fd_pr__special_nfet_pass l=0.140 nf=1 w=0.140

  X1 BL VNB BL VNB sky130_fd_pr__special_nfet_pass l=0.140 nf=1 w=0.140


.ENDS sram_sp_hstrap

.SUBCKT folded_inv_1 vdd vss a y

  XMP0 y a vdd vdd mos_w5000_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w2000_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w5000_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w2000_l150_m1_nf1_id0

.ENDS folded_inv_1

.SUBCKT and2 vdd a b y yb vss

  X0 vdd vss a b yb nand2
  X0_1 vdd vss yb y folded_inv_1

.ENDS and2

.SUBCKT decoder_stage vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y[12] y[13] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] y_b[12] y_b[13] wl_en in[0] in[1] in[2] in[3] in[4] in[5] in[6] in[7] in[8] in[9] in[10] in[11] in[12] in[13]

  Xgate_0_0_0 vdd wl_en in[0] y[0] y_b[0] vss and2
  Xgate_0_1_0 vdd wl_en in[1] y[1] y_b[1] vss and2
  Xgate_0_2_0 vdd wl_en in[2] y[2] y_b[2] vss and2
  Xgate_0_3_0 vdd wl_en in[3] y[3] y_b[3] vss and2
  Xgate_0_4_0 vdd wl_en in[4] y[4] y_b[4] vss and2
  Xgate_0_5_0 vdd wl_en in[5] y[5] y_b[5] vss and2
  Xgate_0_6_0 vdd wl_en in[6] y[6] y_b[6] vss and2
  Xgate_0_7_0 vdd wl_en in[7] y[7] y_b[7] vss and2
  Xgate_0_8_0 vdd wl_en in[8] y[8] y_b[8] vss and2
  Xgate_0_9_0 vdd wl_en in[9] y[9] y_b[9] vss and2
  Xgate_0_10_0 vdd wl_en in[10] y[10] y_b[10] vss and2
  Xgate_0_11_0 vdd wl_en in[11] y[11] y_b[11] vss and2
  Xgate_0_12_0 vdd wl_en in[12] y[12] y_b[12] vss and2
  Xgate_0_13_0 vdd wl_en in[13] y[13] y_b[13] vss and2

.ENDS decoder_stage

.SUBCKT decoder_4 vdd vss y[0] y[1] y[2] y[3] y_b[0] y_b[1] y_b[2] y_b[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1

  X0 vdd vss y[0] y[1] y[2] y[3] y_b[0] y_b[1] y_b[2] y_b[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 decoder_stage_10

.ENDS decoder_4

.SUBCKT mos_w2850_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=2.850


.ENDS mos_w2850_l150_m1_nf1_id0

.SUBCKT mos_w3550_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=3.550


.ENDS mos_w3550_l150_m1_nf1_id1

.SUBCKT nand2_2 vdd vss a b y

  Xn1 x a vss vss mos_w2850_l150_m1_nf1_id0
  Xn2 y b x vss mos_w2850_l150_m1_nf1_id0
  Xp1 y a vdd vdd mos_w3550_l150_m1_nf1_id1
  Xp2 y b vdd vdd mos_w3550_l150_m1_nf1_id1

.ENDS nand2_2

.SUBCKT decoder_stage_8 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y[12] y[13] y[14] y[15] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] y_b[12] y_b[13] y_b[14] y_b[15] predecode_0_0 predecode_0_1 predecode_0_2 predecode_0_3 predecode_1_0 predecode_1_1 predecode_1_2 predecode_1_3

  Xgate_0_0_0 vdd vss predecode_0_0 predecode_1_0 y_b[0] nand2_2
  Xgate_0_1_0 vdd vss predecode_0_1 predecode_1_0 y_b[1] nand2_2
  Xgate_0_2_0 vdd vss predecode_0_2 predecode_1_0 y_b[2] nand2_2
  Xgate_0_3_0 vdd vss predecode_0_3 predecode_1_0 y_b[3] nand2_2
  Xgate_0_4_0 vdd vss predecode_0_0 predecode_1_1 y_b[4] nand2_2
  Xgate_0_5_0 vdd vss predecode_0_1 predecode_1_1 y_b[5] nand2_2
  Xgate_0_6_0 vdd vss predecode_0_2 predecode_1_1 y_b[6] nand2_2
  Xgate_0_7_0 vdd vss predecode_0_3 predecode_1_1 y_b[7] nand2_2
  Xgate_0_8_0 vdd vss predecode_0_0 predecode_1_2 y_b[8] nand2_2
  Xgate_0_9_0 vdd vss predecode_0_1 predecode_1_2 y_b[9] nand2_2
  Xgate_0_10_0 vdd vss predecode_0_2 predecode_1_2 y_b[10] nand2_2
  Xgate_0_11_0 vdd vss predecode_0_3 predecode_1_2 y_b[11] nand2_2
  Xgate_0_12_0 vdd vss predecode_0_0 predecode_1_3 y_b[12] nand2_2
  Xgate_0_13_0 vdd vss predecode_0_1 predecode_1_3 y_b[13] nand2_2
  Xgate_0_14_0 vdd vss predecode_0_2 predecode_1_3 y_b[14] nand2_2
  Xgate_0_15_0 vdd vss predecode_0_3 predecode_1_3 y_b[15] nand2_2
  Xgate_1_0_0 vdd vss y_b[0] y[0] folded_inv_4
  Xgate_1_0_1 vdd vss y_b[0] y[0] folded_inv_4
  Xgate_1_1_0 vdd vss y_b[1] y[1] folded_inv_4
  Xgate_1_1_1 vdd vss y_b[1] y[1] folded_inv_4
  Xgate_1_2_0 vdd vss y_b[2] y[2] folded_inv_4
  Xgate_1_2_1 vdd vss y_b[2] y[2] folded_inv_4
  Xgate_1_3_0 vdd vss y_b[3] y[3] folded_inv_4
  Xgate_1_3_1 vdd vss y_b[3] y[3] folded_inv_4
  Xgate_1_4_0 vdd vss y_b[4] y[4] folded_inv_4
  Xgate_1_4_1 vdd vss y_b[4] y[4] folded_inv_4
  Xgate_1_5_0 vdd vss y_b[5] y[5] folded_inv_4
  Xgate_1_5_1 vdd vss y_b[5] y[5] folded_inv_4
  Xgate_1_6_0 vdd vss y_b[6] y[6] folded_inv_4
  Xgate_1_6_1 vdd vss y_b[6] y[6] folded_inv_4
  Xgate_1_7_0 vdd vss y_b[7] y[7] folded_inv_4
  Xgate_1_7_1 vdd vss y_b[7] y[7] folded_inv_4
  Xgate_1_8_0 vdd vss y_b[8] y[8] folded_inv_4
  Xgate_1_8_1 vdd vss y_b[8] y[8] folded_inv_4
  Xgate_1_9_0 vdd vss y_b[9] y[9] folded_inv_4
  Xgate_1_9_1 vdd vss y_b[9] y[9] folded_inv_4
  Xgate_1_10_0 vdd vss y_b[10] y[10] folded_inv_4
  Xgate_1_10_1 vdd vss y_b[10] y[10] folded_inv_4
  Xgate_1_11_0 vdd vss y_b[11] y[11] folded_inv_4
  Xgate_1_11_1 vdd vss y_b[11] y[11] folded_inv_4
  Xgate_1_12_0 vdd vss y_b[12] y[12] folded_inv_4
  Xgate_1_12_1 vdd vss y_b[12] y[12] folded_inv_4
  Xgate_1_13_0 vdd vss y_b[13] y[13] folded_inv_4
  Xgate_1_13_1 vdd vss y_b[13] y[13] folded_inv_4
  Xgate_1_14_0 vdd vss y_b[14] y[14] folded_inv_4
  Xgate_1_14_1 vdd vss y_b[14] y[14] folded_inv_4
  Xgate_1_15_0 vdd vss y_b[15] y[15] folded_inv_4
  Xgate_1_15_1 vdd vss y_b[15] y[15] folded_inv_4

.ENDS decoder_stage_8

.SUBCKT decoder_2 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y[12] y[13] y[14] y[15] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] y_b[12] y_b[13] y_b[14] y_b[15] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 predecode_2_0 predecode_2_1 predecode_3_0 predecode_3_1

  X0 vdd vss child_conn_0[0] child_conn_0[1] child_conn_0[2] child_conn_0[3] child_noconn_0[0] child_noconn_0[1] child_noconn_0[2] child_noconn_0[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 decoder_4
  X0_1 vdd vss child_conn_1[0] child_conn_1[1] child_conn_1[2] child_conn_1[3] child_noconn_1[0] child_noconn_1[1] child_noconn_1[2] child_noconn_1[3] predecode_2_0 predecode_2_1 predecode_3_0 predecode_3_1 decoder_4
  X0_2 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y[12] y[13] y[14] y[15] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] y_b[12] y_b[13] y_b[14] y_b[15] child_conn_0[0] child_conn_0[1] child_conn_0[2] child_conn_0[3] child_conn_1[0] child_conn_1[1] child_conn_1[2] child_conn_1[3] decoder_stage_8

.ENDS decoder_2

.SUBCKT decoder_3 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 predecode_2_0 predecode_2_1

  X0 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 predecode_2_0 predecode_2_1 decoder_stage_9

.ENDS decoder_3

.SUBCKT multi_finger_inv_6 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_6

.SUBCKT multi_finger_inv_7 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_7

.SUBCKT multi_finger_inv_9 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP19 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP20 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP21 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP22 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP23 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP24 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP25 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP26 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP27 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP28 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP29 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP30 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP31 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP32 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP33 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP34 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP35 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP36 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP37 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP38 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP39 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP40 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP41 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP42 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP43 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP44 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP45 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP46 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP47 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP48 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP49 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP50 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP51 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP52 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP53 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP54 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP55 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP56 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN7 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN8 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN9 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN10 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN11 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN12 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN13 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN14 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN15 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN16 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN17 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN18 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN19 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN20 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN21 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN22 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_9

.SUBCKT decoder_stage_5 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y[12] y[13] y[14] y[15] y[16] y[17] y[18] y[19] y[20] y[21] y[22] y[23] y[24] y[25] y[26] y[27] y[28] y[29] y[30] y[31] y[32] y[33] y[34] y[35] y[36] y[37] y[38] y[39] y[40] y[41] y[42] y[43] y[44] y[45] y[46] y[47] y[48] y[49] y[50] y[51] y[52] y[53] y[54] y[55] y[56] y[57] y[58] y[59] y[60] y[61] y[62] y[63] y[64] y[65] y[66] y[67] y[68] y[69] y[70] y[71] y[72] y[73] y[74] y[75] y[76] y[77] y[78] y[79] y[80] y[81] y[82] y[83] y[84] y[85] y[86] y[87] y[88] y[89] y[90] y[91] y[92] y[93] y[94] y[95] y[96] y[97] y[98] y[99] y[100] y[101] y[102] y[103] y[104] y[105] y[106] y[107] y[108] y[109] y[110] y[111] y[112] y[113] y[114] y[115] y[116] y[117] y[118] y[119] y[120] y[121] y[122] y[123] y[124] y[125] y[126] y[127] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] y_b[12] y_b[13] y_b[14] y_b[15] y_b[16] y_b[17] y_b[18] y_b[19] y_b[20] y_b[21] y_b[22] y_b[23] y_b[24] y_b[25] y_b[26] y_b[27] y_b[28] y_b[29] y_b[30] y_b[31] y_b[32] y_b[33] y_b[34] y_b[35] y_b[36] y_b[37] y_b[38] y_b[39] y_b[40] y_b[41] y_b[42] y_b[43] y_b[44] y_b[45] y_b[46] y_b[47] y_b[48] y_b[49] y_b[50] y_b[51] y_b[52] y_b[53] y_b[54] y_b[55] y_b[56] y_b[57] y_b[58] y_b[59] y_b[60] y_b[61] y_b[62] y_b[63] y_b[64] y_b[65] y_b[66] y_b[67] y_b[68] y_b[69] y_b[70] y_b[71] y_b[72] y_b[73] y_b[74] y_b[75] y_b[76] y_b[77] y_b[78] y_b[79] y_b[80] y_b[81] y_b[82] y_b[83] y_b[84] y_b[85] y_b[86] y_b[87] y_b[88] y_b[89] y_b[90] y_b[91] y_b[92] y_b[93] y_b[94] y_b[95] y_b[96] y_b[97] y_b[98] y_b[99] y_b[100] y_b[101] y_b[102] y_b[103] y_b[104] y_b[105] y_b[106] y_b[107] y_b[108] y_b[109] y_b[110] y_b[111] y_b[112] y_b[113] y_b[114] y_b[115] y_b[116] y_b[117] y_b[118] y_b[119] y_b[120] y_b[121] y_b[122] y_b[123] y_b[124] y_b[125] y_b[126] y_b[127] predecode_0_0 predecode_0_1 predecode_0_2 predecode_0_3 predecode_0_4 predecode_0_5 predecode_0_6 predecode_0_7 predecode_0_8 predecode_0_9 predecode_0_10 predecode_0_11 predecode_0_12 predecode_0_13 predecode_0_14 predecode_0_15 predecode_1_0 predecode_1_1 predecode_1_2 predecode_1_3 predecode_1_4 predecode_1_5 predecode_1_6 predecode_1_7

  Xgate_0_0_0 vdd predecode_0_0 predecode_1_0 x_0[0] y_b_noconn_0_0_0 vss and2_1
  Xgate_0_1_0 vdd predecode_0_1 predecode_1_0 x_0[1] y_b_noconn_0_1_0 vss and2_1
  Xgate_0_2_0 vdd predecode_0_2 predecode_1_0 x_0[2] y_b_noconn_0_2_0 vss and2_1
  Xgate_0_3_0 vdd predecode_0_3 predecode_1_0 x_0[3] y_b_noconn_0_3_0 vss and2_1
  Xgate_0_4_0 vdd predecode_0_4 predecode_1_0 x_0[4] y_b_noconn_0_4_0 vss and2_1
  Xgate_0_5_0 vdd predecode_0_5 predecode_1_0 x_0[5] y_b_noconn_0_5_0 vss and2_1
  Xgate_0_6_0 vdd predecode_0_6 predecode_1_0 x_0[6] y_b_noconn_0_6_0 vss and2_1
  Xgate_0_7_0 vdd predecode_0_7 predecode_1_0 x_0[7] y_b_noconn_0_7_0 vss and2_1
  Xgate_0_8_0 vdd predecode_0_8 predecode_1_0 x_0[8] y_b_noconn_0_8_0 vss and2_1
  Xgate_0_9_0 vdd predecode_0_9 predecode_1_0 x_0[9] y_b_noconn_0_9_0 vss and2_1
  Xgate_0_10_0 vdd predecode_0_10 predecode_1_0 x_0[10] y_b_noconn_0_10_0 vss and2_1
  Xgate_0_11_0 vdd predecode_0_11 predecode_1_0 x_0[11] y_b_noconn_0_11_0 vss and2_1
  Xgate_0_12_0 vdd predecode_0_12 predecode_1_0 x_0[12] y_b_noconn_0_12_0 vss and2_1
  Xgate_0_13_0 vdd predecode_0_13 predecode_1_0 x_0[13] y_b_noconn_0_13_0 vss and2_1
  Xgate_0_14_0 vdd predecode_0_14 predecode_1_0 x_0[14] y_b_noconn_0_14_0 vss and2_1
  Xgate_0_15_0 vdd predecode_0_15 predecode_1_0 x_0[15] y_b_noconn_0_15_0 vss and2_1
  Xgate_0_16_0 vdd predecode_0_0 predecode_1_1 x_0[16] y_b_noconn_0_16_0 vss and2_1
  Xgate_0_17_0 vdd predecode_0_1 predecode_1_1 x_0[17] y_b_noconn_0_17_0 vss and2_1
  Xgate_0_18_0 vdd predecode_0_2 predecode_1_1 x_0[18] y_b_noconn_0_18_0 vss and2_1
  Xgate_0_19_0 vdd predecode_0_3 predecode_1_1 x_0[19] y_b_noconn_0_19_0 vss and2_1
  Xgate_0_20_0 vdd predecode_0_4 predecode_1_1 x_0[20] y_b_noconn_0_20_0 vss and2_1
  Xgate_0_21_0 vdd predecode_0_5 predecode_1_1 x_0[21] y_b_noconn_0_21_0 vss and2_1
  Xgate_0_22_0 vdd predecode_0_6 predecode_1_1 x_0[22] y_b_noconn_0_22_0 vss and2_1
  Xgate_0_23_0 vdd predecode_0_7 predecode_1_1 x_0[23] y_b_noconn_0_23_0 vss and2_1
  Xgate_0_24_0 vdd predecode_0_8 predecode_1_1 x_0[24] y_b_noconn_0_24_0 vss and2_1
  Xgate_0_25_0 vdd predecode_0_9 predecode_1_1 x_0[25] y_b_noconn_0_25_0 vss and2_1
  Xgate_0_26_0 vdd predecode_0_10 predecode_1_1 x_0[26] y_b_noconn_0_26_0 vss and2_1
  Xgate_0_27_0 vdd predecode_0_11 predecode_1_1 x_0[27] y_b_noconn_0_27_0 vss and2_1
  Xgate_0_28_0 vdd predecode_0_12 predecode_1_1 x_0[28] y_b_noconn_0_28_0 vss and2_1
  Xgate_0_29_0 vdd predecode_0_13 predecode_1_1 x_0[29] y_b_noconn_0_29_0 vss and2_1
  Xgate_0_30_0 vdd predecode_0_14 predecode_1_1 x_0[30] y_b_noconn_0_30_0 vss and2_1
  Xgate_0_31_0 vdd predecode_0_15 predecode_1_1 x_0[31] y_b_noconn_0_31_0 vss and2_1
  Xgate_0_32_0 vdd predecode_0_0 predecode_1_2 x_0[32] y_b_noconn_0_32_0 vss and2_1
  Xgate_0_33_0 vdd predecode_0_1 predecode_1_2 x_0[33] y_b_noconn_0_33_0 vss and2_1
  Xgate_0_34_0 vdd predecode_0_2 predecode_1_2 x_0[34] y_b_noconn_0_34_0 vss and2_1
  Xgate_0_35_0 vdd predecode_0_3 predecode_1_2 x_0[35] y_b_noconn_0_35_0 vss and2_1
  Xgate_0_36_0 vdd predecode_0_4 predecode_1_2 x_0[36] y_b_noconn_0_36_0 vss and2_1
  Xgate_0_37_0 vdd predecode_0_5 predecode_1_2 x_0[37] y_b_noconn_0_37_0 vss and2_1
  Xgate_0_38_0 vdd predecode_0_6 predecode_1_2 x_0[38] y_b_noconn_0_38_0 vss and2_1
  Xgate_0_39_0 vdd predecode_0_7 predecode_1_2 x_0[39] y_b_noconn_0_39_0 vss and2_1
  Xgate_0_40_0 vdd predecode_0_8 predecode_1_2 x_0[40] y_b_noconn_0_40_0 vss and2_1
  Xgate_0_41_0 vdd predecode_0_9 predecode_1_2 x_0[41] y_b_noconn_0_41_0 vss and2_1
  Xgate_0_42_0 vdd predecode_0_10 predecode_1_2 x_0[42] y_b_noconn_0_42_0 vss and2_1
  Xgate_0_43_0 vdd predecode_0_11 predecode_1_2 x_0[43] y_b_noconn_0_43_0 vss and2_1
  Xgate_0_44_0 vdd predecode_0_12 predecode_1_2 x_0[44] y_b_noconn_0_44_0 vss and2_1
  Xgate_0_45_0 vdd predecode_0_13 predecode_1_2 x_0[45] y_b_noconn_0_45_0 vss and2_1
  Xgate_0_46_0 vdd predecode_0_14 predecode_1_2 x_0[46] y_b_noconn_0_46_0 vss and2_1
  Xgate_0_47_0 vdd predecode_0_15 predecode_1_2 x_0[47] y_b_noconn_0_47_0 vss and2_1
  Xgate_0_48_0 vdd predecode_0_0 predecode_1_3 x_0[48] y_b_noconn_0_48_0 vss and2_1
  Xgate_0_49_0 vdd predecode_0_1 predecode_1_3 x_0[49] y_b_noconn_0_49_0 vss and2_1
  Xgate_0_50_0 vdd predecode_0_2 predecode_1_3 x_0[50] y_b_noconn_0_50_0 vss and2_1
  Xgate_0_51_0 vdd predecode_0_3 predecode_1_3 x_0[51] y_b_noconn_0_51_0 vss and2_1
  Xgate_0_52_0 vdd predecode_0_4 predecode_1_3 x_0[52] y_b_noconn_0_52_0 vss and2_1
  Xgate_0_53_0 vdd predecode_0_5 predecode_1_3 x_0[53] y_b_noconn_0_53_0 vss and2_1
  Xgate_0_54_0 vdd predecode_0_6 predecode_1_3 x_0[54] y_b_noconn_0_54_0 vss and2_1
  Xgate_0_55_0 vdd predecode_0_7 predecode_1_3 x_0[55] y_b_noconn_0_55_0 vss and2_1
  Xgate_0_56_0 vdd predecode_0_8 predecode_1_3 x_0[56] y_b_noconn_0_56_0 vss and2_1
  Xgate_0_57_0 vdd predecode_0_9 predecode_1_3 x_0[57] y_b_noconn_0_57_0 vss and2_1
  Xgate_0_58_0 vdd predecode_0_10 predecode_1_3 x_0[58] y_b_noconn_0_58_0 vss and2_1
  Xgate_0_59_0 vdd predecode_0_11 predecode_1_3 x_0[59] y_b_noconn_0_59_0 vss and2_1
  Xgate_0_60_0 vdd predecode_0_12 predecode_1_3 x_0[60] y_b_noconn_0_60_0 vss and2_1
  Xgate_0_61_0 vdd predecode_0_13 predecode_1_3 x_0[61] y_b_noconn_0_61_0 vss and2_1
  Xgate_0_62_0 vdd predecode_0_14 predecode_1_3 x_0[62] y_b_noconn_0_62_0 vss and2_1
  Xgate_0_63_0 vdd predecode_0_15 predecode_1_3 x_0[63] y_b_noconn_0_63_0 vss and2_1
  Xgate_0_64_0 vdd predecode_0_0 predecode_1_4 x_0[64] y_b_noconn_0_64_0 vss and2_1
  Xgate_0_65_0 vdd predecode_0_1 predecode_1_4 x_0[65] y_b_noconn_0_65_0 vss and2_1
  Xgate_0_66_0 vdd predecode_0_2 predecode_1_4 x_0[66] y_b_noconn_0_66_0 vss and2_1
  Xgate_0_67_0 vdd predecode_0_3 predecode_1_4 x_0[67] y_b_noconn_0_67_0 vss and2_1
  Xgate_0_68_0 vdd predecode_0_4 predecode_1_4 x_0[68] y_b_noconn_0_68_0 vss and2_1
  Xgate_0_69_0 vdd predecode_0_5 predecode_1_4 x_0[69] y_b_noconn_0_69_0 vss and2_1
  Xgate_0_70_0 vdd predecode_0_6 predecode_1_4 x_0[70] y_b_noconn_0_70_0 vss and2_1
  Xgate_0_71_0 vdd predecode_0_7 predecode_1_4 x_0[71] y_b_noconn_0_71_0 vss and2_1
  Xgate_0_72_0 vdd predecode_0_8 predecode_1_4 x_0[72] y_b_noconn_0_72_0 vss and2_1
  Xgate_0_73_0 vdd predecode_0_9 predecode_1_4 x_0[73] y_b_noconn_0_73_0 vss and2_1
  Xgate_0_74_0 vdd predecode_0_10 predecode_1_4 x_0[74] y_b_noconn_0_74_0 vss and2_1
  Xgate_0_75_0 vdd predecode_0_11 predecode_1_4 x_0[75] y_b_noconn_0_75_0 vss and2_1
  Xgate_0_76_0 vdd predecode_0_12 predecode_1_4 x_0[76] y_b_noconn_0_76_0 vss and2_1
  Xgate_0_77_0 vdd predecode_0_13 predecode_1_4 x_0[77] y_b_noconn_0_77_0 vss and2_1
  Xgate_0_78_0 vdd predecode_0_14 predecode_1_4 x_0[78] y_b_noconn_0_78_0 vss and2_1
  Xgate_0_79_0 vdd predecode_0_15 predecode_1_4 x_0[79] y_b_noconn_0_79_0 vss and2_1
  Xgate_0_80_0 vdd predecode_0_0 predecode_1_5 x_0[80] y_b_noconn_0_80_0 vss and2_1
  Xgate_0_81_0 vdd predecode_0_1 predecode_1_5 x_0[81] y_b_noconn_0_81_0 vss and2_1
  Xgate_0_82_0 vdd predecode_0_2 predecode_1_5 x_0[82] y_b_noconn_0_82_0 vss and2_1
  Xgate_0_83_0 vdd predecode_0_3 predecode_1_5 x_0[83] y_b_noconn_0_83_0 vss and2_1
  Xgate_0_84_0 vdd predecode_0_4 predecode_1_5 x_0[84] y_b_noconn_0_84_0 vss and2_1
  Xgate_0_85_0 vdd predecode_0_5 predecode_1_5 x_0[85] y_b_noconn_0_85_0 vss and2_1
  Xgate_0_86_0 vdd predecode_0_6 predecode_1_5 x_0[86] y_b_noconn_0_86_0 vss and2_1
  Xgate_0_87_0 vdd predecode_0_7 predecode_1_5 x_0[87] y_b_noconn_0_87_0 vss and2_1
  Xgate_0_88_0 vdd predecode_0_8 predecode_1_5 x_0[88] y_b_noconn_0_88_0 vss and2_1
  Xgate_0_89_0 vdd predecode_0_9 predecode_1_5 x_0[89] y_b_noconn_0_89_0 vss and2_1
  Xgate_0_90_0 vdd predecode_0_10 predecode_1_5 x_0[90] y_b_noconn_0_90_0 vss and2_1
  Xgate_0_91_0 vdd predecode_0_11 predecode_1_5 x_0[91] y_b_noconn_0_91_0 vss and2_1
  Xgate_0_92_0 vdd predecode_0_12 predecode_1_5 x_0[92] y_b_noconn_0_92_0 vss and2_1
  Xgate_0_93_0 vdd predecode_0_13 predecode_1_5 x_0[93] y_b_noconn_0_93_0 vss and2_1
  Xgate_0_94_0 vdd predecode_0_14 predecode_1_5 x_0[94] y_b_noconn_0_94_0 vss and2_1
  Xgate_0_95_0 vdd predecode_0_15 predecode_1_5 x_0[95] y_b_noconn_0_95_0 vss and2_1
  Xgate_0_96_0 vdd predecode_0_0 predecode_1_6 x_0[96] y_b_noconn_0_96_0 vss and2_1
  Xgate_0_97_0 vdd predecode_0_1 predecode_1_6 x_0[97] y_b_noconn_0_97_0 vss and2_1
  Xgate_0_98_0 vdd predecode_0_2 predecode_1_6 x_0[98] y_b_noconn_0_98_0 vss and2_1
  Xgate_0_99_0 vdd predecode_0_3 predecode_1_6 x_0[99] y_b_noconn_0_99_0 vss and2_1
  Xgate_0_100_0 vdd predecode_0_4 predecode_1_6 x_0[100] y_b_noconn_0_100_0 vss and2_1
  Xgate_0_101_0 vdd predecode_0_5 predecode_1_6 x_0[101] y_b_noconn_0_101_0 vss and2_1
  Xgate_0_102_0 vdd predecode_0_6 predecode_1_6 x_0[102] y_b_noconn_0_102_0 vss and2_1
  Xgate_0_103_0 vdd predecode_0_7 predecode_1_6 x_0[103] y_b_noconn_0_103_0 vss and2_1
  Xgate_0_104_0 vdd predecode_0_8 predecode_1_6 x_0[104] y_b_noconn_0_104_0 vss and2_1
  Xgate_0_105_0 vdd predecode_0_9 predecode_1_6 x_0[105] y_b_noconn_0_105_0 vss and2_1
  Xgate_0_106_0 vdd predecode_0_10 predecode_1_6 x_0[106] y_b_noconn_0_106_0 vss and2_1
  Xgate_0_107_0 vdd predecode_0_11 predecode_1_6 x_0[107] y_b_noconn_0_107_0 vss and2_1
  Xgate_0_108_0 vdd predecode_0_12 predecode_1_6 x_0[108] y_b_noconn_0_108_0 vss and2_1
  Xgate_0_109_0 vdd predecode_0_13 predecode_1_6 x_0[109] y_b_noconn_0_109_0 vss and2_1
  Xgate_0_110_0 vdd predecode_0_14 predecode_1_6 x_0[110] y_b_noconn_0_110_0 vss and2_1
  Xgate_0_111_0 vdd predecode_0_15 predecode_1_6 x_0[111] y_b_noconn_0_111_0 vss and2_1
  Xgate_0_112_0 vdd predecode_0_0 predecode_1_7 x_0[112] y_b_noconn_0_112_0 vss and2_1
  Xgate_0_113_0 vdd predecode_0_1 predecode_1_7 x_0[113] y_b_noconn_0_113_0 vss and2_1
  Xgate_0_114_0 vdd predecode_0_2 predecode_1_7 x_0[114] y_b_noconn_0_114_0 vss and2_1
  Xgate_0_115_0 vdd predecode_0_3 predecode_1_7 x_0[115] y_b_noconn_0_115_0 vss and2_1
  Xgate_0_116_0 vdd predecode_0_4 predecode_1_7 x_0[116] y_b_noconn_0_116_0 vss and2_1
  Xgate_0_117_0 vdd predecode_0_5 predecode_1_7 x_0[117] y_b_noconn_0_117_0 vss and2_1
  Xgate_0_118_0 vdd predecode_0_6 predecode_1_7 x_0[118] y_b_noconn_0_118_0 vss and2_1
  Xgate_0_119_0 vdd predecode_0_7 predecode_1_7 x_0[119] y_b_noconn_0_119_0 vss and2_1
  Xgate_0_120_0 vdd predecode_0_8 predecode_1_7 x_0[120] y_b_noconn_0_120_0 vss and2_1
  Xgate_0_121_0 vdd predecode_0_9 predecode_1_7 x_0[121] y_b_noconn_0_121_0 vss and2_1
  Xgate_0_122_0 vdd predecode_0_10 predecode_1_7 x_0[122] y_b_noconn_0_122_0 vss and2_1
  Xgate_0_123_0 vdd predecode_0_11 predecode_1_7 x_0[123] y_b_noconn_0_123_0 vss and2_1
  Xgate_0_124_0 vdd predecode_0_12 predecode_1_7 x_0[124] y_b_noconn_0_124_0 vss and2_1
  Xgate_0_125_0 vdd predecode_0_13 predecode_1_7 x_0[125] y_b_noconn_0_125_0 vss and2_1
  Xgate_0_126_0 vdd predecode_0_14 predecode_1_7 x_0[126] y_b_noconn_0_126_0 vss and2_1
  Xgate_0_127_0 vdd predecode_0_15 predecode_1_7 x_0[127] y_b_noconn_0_127_0 vss and2_1
  Xgate_1_0_0 vdd vss x_0[0] x_1[0] multi_finger_inv_6
  Xgate_1_1_0 vdd vss x_0[1] x_1[1] multi_finger_inv_6
  Xgate_1_2_0 vdd vss x_0[2] x_1[2] multi_finger_inv_6
  Xgate_1_3_0 vdd vss x_0[3] x_1[3] multi_finger_inv_6
  Xgate_1_4_0 vdd vss x_0[4] x_1[4] multi_finger_inv_6
  Xgate_1_5_0 vdd vss x_0[5] x_1[5] multi_finger_inv_6
  Xgate_1_6_0 vdd vss x_0[6] x_1[6] multi_finger_inv_6
  Xgate_1_7_0 vdd vss x_0[7] x_1[7] multi_finger_inv_6
  Xgate_1_8_0 vdd vss x_0[8] x_1[8] multi_finger_inv_6
  Xgate_1_9_0 vdd vss x_0[9] x_1[9] multi_finger_inv_6
  Xgate_1_10_0 vdd vss x_0[10] x_1[10] multi_finger_inv_6
  Xgate_1_11_0 vdd vss x_0[11] x_1[11] multi_finger_inv_6
  Xgate_1_12_0 vdd vss x_0[12] x_1[12] multi_finger_inv_6
  Xgate_1_13_0 vdd vss x_0[13] x_1[13] multi_finger_inv_6
  Xgate_1_14_0 vdd vss x_0[14] x_1[14] multi_finger_inv_6
  Xgate_1_15_0 vdd vss x_0[15] x_1[15] multi_finger_inv_6
  Xgate_1_16_0 vdd vss x_0[16] x_1[16] multi_finger_inv_6
  Xgate_1_17_0 vdd vss x_0[17] x_1[17] multi_finger_inv_6
  Xgate_1_18_0 vdd vss x_0[18] x_1[18] multi_finger_inv_6
  Xgate_1_19_0 vdd vss x_0[19] x_1[19] multi_finger_inv_6
  Xgate_1_20_0 vdd vss x_0[20] x_1[20] multi_finger_inv_6
  Xgate_1_21_0 vdd vss x_0[21] x_1[21] multi_finger_inv_6
  Xgate_1_22_0 vdd vss x_0[22] x_1[22] multi_finger_inv_6
  Xgate_1_23_0 vdd vss x_0[23] x_1[23] multi_finger_inv_6
  Xgate_1_24_0 vdd vss x_0[24] x_1[24] multi_finger_inv_6
  Xgate_1_25_0 vdd vss x_0[25] x_1[25] multi_finger_inv_6
  Xgate_1_26_0 vdd vss x_0[26] x_1[26] multi_finger_inv_6
  Xgate_1_27_0 vdd vss x_0[27] x_1[27] multi_finger_inv_6
  Xgate_1_28_0 vdd vss x_0[28] x_1[28] multi_finger_inv_6
  Xgate_1_29_0 vdd vss x_0[29] x_1[29] multi_finger_inv_6
  Xgate_1_30_0 vdd vss x_0[30] x_1[30] multi_finger_inv_6
  Xgate_1_31_0 vdd vss x_0[31] x_1[31] multi_finger_inv_6
  Xgate_1_32_0 vdd vss x_0[32] x_1[32] multi_finger_inv_6
  Xgate_1_33_0 vdd vss x_0[33] x_1[33] multi_finger_inv_6
  Xgate_1_34_0 vdd vss x_0[34] x_1[34] multi_finger_inv_6
  Xgate_1_35_0 vdd vss x_0[35] x_1[35] multi_finger_inv_6
  Xgate_1_36_0 vdd vss x_0[36] x_1[36] multi_finger_inv_6
  Xgate_1_37_0 vdd vss x_0[37] x_1[37] multi_finger_inv_6
  Xgate_1_38_0 vdd vss x_0[38] x_1[38] multi_finger_inv_6
  Xgate_1_39_0 vdd vss x_0[39] x_1[39] multi_finger_inv_6
  Xgate_1_40_0 vdd vss x_0[40] x_1[40] multi_finger_inv_6
  Xgate_1_41_0 vdd vss x_0[41] x_1[41] multi_finger_inv_6
  Xgate_1_42_0 vdd vss x_0[42] x_1[42] multi_finger_inv_6
  Xgate_1_43_0 vdd vss x_0[43] x_1[43] multi_finger_inv_6
  Xgate_1_44_0 vdd vss x_0[44] x_1[44] multi_finger_inv_6
  Xgate_1_45_0 vdd vss x_0[45] x_1[45] multi_finger_inv_6
  Xgate_1_46_0 vdd vss x_0[46] x_1[46] multi_finger_inv_6
  Xgate_1_47_0 vdd vss x_0[47] x_1[47] multi_finger_inv_6
  Xgate_1_48_0 vdd vss x_0[48] x_1[48] multi_finger_inv_6
  Xgate_1_49_0 vdd vss x_0[49] x_1[49] multi_finger_inv_6
  Xgate_1_50_0 vdd vss x_0[50] x_1[50] multi_finger_inv_6
  Xgate_1_51_0 vdd vss x_0[51] x_1[51] multi_finger_inv_6
  Xgate_1_52_0 vdd vss x_0[52] x_1[52] multi_finger_inv_6
  Xgate_1_53_0 vdd vss x_0[53] x_1[53] multi_finger_inv_6
  Xgate_1_54_0 vdd vss x_0[54] x_1[54] multi_finger_inv_6
  Xgate_1_55_0 vdd vss x_0[55] x_1[55] multi_finger_inv_6
  Xgate_1_56_0 vdd vss x_0[56] x_1[56] multi_finger_inv_6
  Xgate_1_57_0 vdd vss x_0[57] x_1[57] multi_finger_inv_6
  Xgate_1_58_0 vdd vss x_0[58] x_1[58] multi_finger_inv_6
  Xgate_1_59_0 vdd vss x_0[59] x_1[59] multi_finger_inv_6
  Xgate_1_60_0 vdd vss x_0[60] x_1[60] multi_finger_inv_6
  Xgate_1_61_0 vdd vss x_0[61] x_1[61] multi_finger_inv_6
  Xgate_1_62_0 vdd vss x_0[62] x_1[62] multi_finger_inv_6
  Xgate_1_63_0 vdd vss x_0[63] x_1[63] multi_finger_inv_6
  Xgate_1_64_0 vdd vss x_0[64] x_1[64] multi_finger_inv_6
  Xgate_1_65_0 vdd vss x_0[65] x_1[65] multi_finger_inv_6
  Xgate_1_66_0 vdd vss x_0[66] x_1[66] multi_finger_inv_6
  Xgate_1_67_0 vdd vss x_0[67] x_1[67] multi_finger_inv_6
  Xgate_1_68_0 vdd vss x_0[68] x_1[68] multi_finger_inv_6
  Xgate_1_69_0 vdd vss x_0[69] x_1[69] multi_finger_inv_6
  Xgate_1_70_0 vdd vss x_0[70] x_1[70] multi_finger_inv_6
  Xgate_1_71_0 vdd vss x_0[71] x_1[71] multi_finger_inv_6
  Xgate_1_72_0 vdd vss x_0[72] x_1[72] multi_finger_inv_6
  Xgate_1_73_0 vdd vss x_0[73] x_1[73] multi_finger_inv_6
  Xgate_1_74_0 vdd vss x_0[74] x_1[74] multi_finger_inv_6
  Xgate_1_75_0 vdd vss x_0[75] x_1[75] multi_finger_inv_6
  Xgate_1_76_0 vdd vss x_0[76] x_1[76] multi_finger_inv_6
  Xgate_1_77_0 vdd vss x_0[77] x_1[77] multi_finger_inv_6
  Xgate_1_78_0 vdd vss x_0[78] x_1[78] multi_finger_inv_6
  Xgate_1_79_0 vdd vss x_0[79] x_1[79] multi_finger_inv_6
  Xgate_1_80_0 vdd vss x_0[80] x_1[80] multi_finger_inv_6
  Xgate_1_81_0 vdd vss x_0[81] x_1[81] multi_finger_inv_6
  Xgate_1_82_0 vdd vss x_0[82] x_1[82] multi_finger_inv_6
  Xgate_1_83_0 vdd vss x_0[83] x_1[83] multi_finger_inv_6
  Xgate_1_84_0 vdd vss x_0[84] x_1[84] multi_finger_inv_6
  Xgate_1_85_0 vdd vss x_0[85] x_1[85] multi_finger_inv_6
  Xgate_1_86_0 vdd vss x_0[86] x_1[86] multi_finger_inv_6
  Xgate_1_87_0 vdd vss x_0[87] x_1[87] multi_finger_inv_6
  Xgate_1_88_0 vdd vss x_0[88] x_1[88] multi_finger_inv_6
  Xgate_1_89_0 vdd vss x_0[89] x_1[89] multi_finger_inv_6
  Xgate_1_90_0 vdd vss x_0[90] x_1[90] multi_finger_inv_6
  Xgate_1_91_0 vdd vss x_0[91] x_1[91] multi_finger_inv_6
  Xgate_1_92_0 vdd vss x_0[92] x_1[92] multi_finger_inv_6
  Xgate_1_93_0 vdd vss x_0[93] x_1[93] multi_finger_inv_6
  Xgate_1_94_0 vdd vss x_0[94] x_1[94] multi_finger_inv_6
  Xgate_1_95_0 vdd vss x_0[95] x_1[95] multi_finger_inv_6
  Xgate_1_96_0 vdd vss x_0[96] x_1[96] multi_finger_inv_6
  Xgate_1_97_0 vdd vss x_0[97] x_1[97] multi_finger_inv_6
  Xgate_1_98_0 vdd vss x_0[98] x_1[98] multi_finger_inv_6
  Xgate_1_99_0 vdd vss x_0[99] x_1[99] multi_finger_inv_6
  Xgate_1_100_0 vdd vss x_0[100] x_1[100] multi_finger_inv_6
  Xgate_1_101_0 vdd vss x_0[101] x_1[101] multi_finger_inv_6
  Xgate_1_102_0 vdd vss x_0[102] x_1[102] multi_finger_inv_6
  Xgate_1_103_0 vdd vss x_0[103] x_1[103] multi_finger_inv_6
  Xgate_1_104_0 vdd vss x_0[104] x_1[104] multi_finger_inv_6
  Xgate_1_105_0 vdd vss x_0[105] x_1[105] multi_finger_inv_6
  Xgate_1_106_0 vdd vss x_0[106] x_1[106] multi_finger_inv_6
  Xgate_1_107_0 vdd vss x_0[107] x_1[107] multi_finger_inv_6
  Xgate_1_108_0 vdd vss x_0[108] x_1[108] multi_finger_inv_6
  Xgate_1_109_0 vdd vss x_0[109] x_1[109] multi_finger_inv_6
  Xgate_1_110_0 vdd vss x_0[110] x_1[110] multi_finger_inv_6
  Xgate_1_111_0 vdd vss x_0[111] x_1[111] multi_finger_inv_6
  Xgate_1_112_0 vdd vss x_0[112] x_1[112] multi_finger_inv_6
  Xgate_1_113_0 vdd vss x_0[113] x_1[113] multi_finger_inv_6
  Xgate_1_114_0 vdd vss x_0[114] x_1[114] multi_finger_inv_6
  Xgate_1_115_0 vdd vss x_0[115] x_1[115] multi_finger_inv_6
  Xgate_1_116_0 vdd vss x_0[116] x_1[116] multi_finger_inv_6
  Xgate_1_117_0 vdd vss x_0[117] x_1[117] multi_finger_inv_6
  Xgate_1_118_0 vdd vss x_0[118] x_1[118] multi_finger_inv_6
  Xgate_1_119_0 vdd vss x_0[119] x_1[119] multi_finger_inv_6
  Xgate_1_120_0 vdd vss x_0[120] x_1[120] multi_finger_inv_6
  Xgate_1_121_0 vdd vss x_0[121] x_1[121] multi_finger_inv_6
  Xgate_1_122_0 vdd vss x_0[122] x_1[122] multi_finger_inv_6
  Xgate_1_123_0 vdd vss x_0[123] x_1[123] multi_finger_inv_6
  Xgate_1_124_0 vdd vss x_0[124] x_1[124] multi_finger_inv_6
  Xgate_1_125_0 vdd vss x_0[125] x_1[125] multi_finger_inv_6
  Xgate_1_126_0 vdd vss x_0[126] x_1[126] multi_finger_inv_6
  Xgate_1_127_0 vdd vss x_0[127] x_1[127] multi_finger_inv_6
  Xgate_2_0_0 vdd vss x_1[0] x_2[0] multi_finger_inv_7
  Xgate_2_1_0 vdd vss x_1[1] x_2[1] multi_finger_inv_7
  Xgate_2_2_0 vdd vss x_1[2] x_2[2] multi_finger_inv_7
  Xgate_2_3_0 vdd vss x_1[3] x_2[3] multi_finger_inv_7
  Xgate_2_4_0 vdd vss x_1[4] x_2[4] multi_finger_inv_7
  Xgate_2_5_0 vdd vss x_1[5] x_2[5] multi_finger_inv_7
  Xgate_2_6_0 vdd vss x_1[6] x_2[6] multi_finger_inv_7
  Xgate_2_7_0 vdd vss x_1[7] x_2[7] multi_finger_inv_7
  Xgate_2_8_0 vdd vss x_1[8] x_2[8] multi_finger_inv_7
  Xgate_2_9_0 vdd vss x_1[9] x_2[9] multi_finger_inv_7
  Xgate_2_10_0 vdd vss x_1[10] x_2[10] multi_finger_inv_7
  Xgate_2_11_0 vdd vss x_1[11] x_2[11] multi_finger_inv_7
  Xgate_2_12_0 vdd vss x_1[12] x_2[12] multi_finger_inv_7
  Xgate_2_13_0 vdd vss x_1[13] x_2[13] multi_finger_inv_7
  Xgate_2_14_0 vdd vss x_1[14] x_2[14] multi_finger_inv_7
  Xgate_2_15_0 vdd vss x_1[15] x_2[15] multi_finger_inv_7
  Xgate_2_16_0 vdd vss x_1[16] x_2[16] multi_finger_inv_7
  Xgate_2_17_0 vdd vss x_1[17] x_2[17] multi_finger_inv_7
  Xgate_2_18_0 vdd vss x_1[18] x_2[18] multi_finger_inv_7
  Xgate_2_19_0 vdd vss x_1[19] x_2[19] multi_finger_inv_7
  Xgate_2_20_0 vdd vss x_1[20] x_2[20] multi_finger_inv_7
  Xgate_2_21_0 vdd vss x_1[21] x_2[21] multi_finger_inv_7
  Xgate_2_22_0 vdd vss x_1[22] x_2[22] multi_finger_inv_7
  Xgate_2_23_0 vdd vss x_1[23] x_2[23] multi_finger_inv_7
  Xgate_2_24_0 vdd vss x_1[24] x_2[24] multi_finger_inv_7
  Xgate_2_25_0 vdd vss x_1[25] x_2[25] multi_finger_inv_7
  Xgate_2_26_0 vdd vss x_1[26] x_2[26] multi_finger_inv_7
  Xgate_2_27_0 vdd vss x_1[27] x_2[27] multi_finger_inv_7
  Xgate_2_28_0 vdd vss x_1[28] x_2[28] multi_finger_inv_7
  Xgate_2_29_0 vdd vss x_1[29] x_2[29] multi_finger_inv_7
  Xgate_2_30_0 vdd vss x_1[30] x_2[30] multi_finger_inv_7
  Xgate_2_31_0 vdd vss x_1[31] x_2[31] multi_finger_inv_7
  Xgate_2_32_0 vdd vss x_1[32] x_2[32] multi_finger_inv_7
  Xgate_2_33_0 vdd vss x_1[33] x_2[33] multi_finger_inv_7
  Xgate_2_34_0 vdd vss x_1[34] x_2[34] multi_finger_inv_7
  Xgate_2_35_0 vdd vss x_1[35] x_2[35] multi_finger_inv_7
  Xgate_2_36_0 vdd vss x_1[36] x_2[36] multi_finger_inv_7
  Xgate_2_37_0 vdd vss x_1[37] x_2[37] multi_finger_inv_7
  Xgate_2_38_0 vdd vss x_1[38] x_2[38] multi_finger_inv_7
  Xgate_2_39_0 vdd vss x_1[39] x_2[39] multi_finger_inv_7
  Xgate_2_40_0 vdd vss x_1[40] x_2[40] multi_finger_inv_7
  Xgate_2_41_0 vdd vss x_1[41] x_2[41] multi_finger_inv_7
  Xgate_2_42_0 vdd vss x_1[42] x_2[42] multi_finger_inv_7
  Xgate_2_43_0 vdd vss x_1[43] x_2[43] multi_finger_inv_7
  Xgate_2_44_0 vdd vss x_1[44] x_2[44] multi_finger_inv_7
  Xgate_2_45_0 vdd vss x_1[45] x_2[45] multi_finger_inv_7
  Xgate_2_46_0 vdd vss x_1[46] x_2[46] multi_finger_inv_7
  Xgate_2_47_0 vdd vss x_1[47] x_2[47] multi_finger_inv_7
  Xgate_2_48_0 vdd vss x_1[48] x_2[48] multi_finger_inv_7
  Xgate_2_49_0 vdd vss x_1[49] x_2[49] multi_finger_inv_7
  Xgate_2_50_0 vdd vss x_1[50] x_2[50] multi_finger_inv_7
  Xgate_2_51_0 vdd vss x_1[51] x_2[51] multi_finger_inv_7
  Xgate_2_52_0 vdd vss x_1[52] x_2[52] multi_finger_inv_7
  Xgate_2_53_0 vdd vss x_1[53] x_2[53] multi_finger_inv_7
  Xgate_2_54_0 vdd vss x_1[54] x_2[54] multi_finger_inv_7
  Xgate_2_55_0 vdd vss x_1[55] x_2[55] multi_finger_inv_7
  Xgate_2_56_0 vdd vss x_1[56] x_2[56] multi_finger_inv_7
  Xgate_2_57_0 vdd vss x_1[57] x_2[57] multi_finger_inv_7
  Xgate_2_58_0 vdd vss x_1[58] x_2[58] multi_finger_inv_7
  Xgate_2_59_0 vdd vss x_1[59] x_2[59] multi_finger_inv_7
  Xgate_2_60_0 vdd vss x_1[60] x_2[60] multi_finger_inv_7
  Xgate_2_61_0 vdd vss x_1[61] x_2[61] multi_finger_inv_7
  Xgate_2_62_0 vdd vss x_1[62] x_2[62] multi_finger_inv_7
  Xgate_2_63_0 vdd vss x_1[63] x_2[63] multi_finger_inv_7
  Xgate_2_64_0 vdd vss x_1[64] x_2[64] multi_finger_inv_7
  Xgate_2_65_0 vdd vss x_1[65] x_2[65] multi_finger_inv_7
  Xgate_2_66_0 vdd vss x_1[66] x_2[66] multi_finger_inv_7
  Xgate_2_67_0 vdd vss x_1[67] x_2[67] multi_finger_inv_7
  Xgate_2_68_0 vdd vss x_1[68] x_2[68] multi_finger_inv_7
  Xgate_2_69_0 vdd vss x_1[69] x_2[69] multi_finger_inv_7
  Xgate_2_70_0 vdd vss x_1[70] x_2[70] multi_finger_inv_7
  Xgate_2_71_0 vdd vss x_1[71] x_2[71] multi_finger_inv_7
  Xgate_2_72_0 vdd vss x_1[72] x_2[72] multi_finger_inv_7
  Xgate_2_73_0 vdd vss x_1[73] x_2[73] multi_finger_inv_7
  Xgate_2_74_0 vdd vss x_1[74] x_2[74] multi_finger_inv_7
  Xgate_2_75_0 vdd vss x_1[75] x_2[75] multi_finger_inv_7
  Xgate_2_76_0 vdd vss x_1[76] x_2[76] multi_finger_inv_7
  Xgate_2_77_0 vdd vss x_1[77] x_2[77] multi_finger_inv_7
  Xgate_2_78_0 vdd vss x_1[78] x_2[78] multi_finger_inv_7
  Xgate_2_79_0 vdd vss x_1[79] x_2[79] multi_finger_inv_7
  Xgate_2_80_0 vdd vss x_1[80] x_2[80] multi_finger_inv_7
  Xgate_2_81_0 vdd vss x_1[81] x_2[81] multi_finger_inv_7
  Xgate_2_82_0 vdd vss x_1[82] x_2[82] multi_finger_inv_7
  Xgate_2_83_0 vdd vss x_1[83] x_2[83] multi_finger_inv_7
  Xgate_2_84_0 vdd vss x_1[84] x_2[84] multi_finger_inv_7
  Xgate_2_85_0 vdd vss x_1[85] x_2[85] multi_finger_inv_7
  Xgate_2_86_0 vdd vss x_1[86] x_2[86] multi_finger_inv_7
  Xgate_2_87_0 vdd vss x_1[87] x_2[87] multi_finger_inv_7
  Xgate_2_88_0 vdd vss x_1[88] x_2[88] multi_finger_inv_7
  Xgate_2_89_0 vdd vss x_1[89] x_2[89] multi_finger_inv_7
  Xgate_2_90_0 vdd vss x_1[90] x_2[90] multi_finger_inv_7
  Xgate_2_91_0 vdd vss x_1[91] x_2[91] multi_finger_inv_7
  Xgate_2_92_0 vdd vss x_1[92] x_2[92] multi_finger_inv_7
  Xgate_2_93_0 vdd vss x_1[93] x_2[93] multi_finger_inv_7
  Xgate_2_94_0 vdd vss x_1[94] x_2[94] multi_finger_inv_7
  Xgate_2_95_0 vdd vss x_1[95] x_2[95] multi_finger_inv_7
  Xgate_2_96_0 vdd vss x_1[96] x_2[96] multi_finger_inv_7
  Xgate_2_97_0 vdd vss x_1[97] x_2[97] multi_finger_inv_7
  Xgate_2_98_0 vdd vss x_1[98] x_2[98] multi_finger_inv_7
  Xgate_2_99_0 vdd vss x_1[99] x_2[99] multi_finger_inv_7
  Xgate_2_100_0 vdd vss x_1[100] x_2[100] multi_finger_inv_7
  Xgate_2_101_0 vdd vss x_1[101] x_2[101] multi_finger_inv_7
  Xgate_2_102_0 vdd vss x_1[102] x_2[102] multi_finger_inv_7
  Xgate_2_103_0 vdd vss x_1[103] x_2[103] multi_finger_inv_7
  Xgate_2_104_0 vdd vss x_1[104] x_2[104] multi_finger_inv_7
  Xgate_2_105_0 vdd vss x_1[105] x_2[105] multi_finger_inv_7
  Xgate_2_106_0 vdd vss x_1[106] x_2[106] multi_finger_inv_7
  Xgate_2_107_0 vdd vss x_1[107] x_2[107] multi_finger_inv_7
  Xgate_2_108_0 vdd vss x_1[108] x_2[108] multi_finger_inv_7
  Xgate_2_109_0 vdd vss x_1[109] x_2[109] multi_finger_inv_7
  Xgate_2_110_0 vdd vss x_1[110] x_2[110] multi_finger_inv_7
  Xgate_2_111_0 vdd vss x_1[111] x_2[111] multi_finger_inv_7
  Xgate_2_112_0 vdd vss x_1[112] x_2[112] multi_finger_inv_7
  Xgate_2_113_0 vdd vss x_1[113] x_2[113] multi_finger_inv_7
  Xgate_2_114_0 vdd vss x_1[114] x_2[114] multi_finger_inv_7
  Xgate_2_115_0 vdd vss x_1[115] x_2[115] multi_finger_inv_7
  Xgate_2_116_0 vdd vss x_1[116] x_2[116] multi_finger_inv_7
  Xgate_2_117_0 vdd vss x_1[117] x_2[117] multi_finger_inv_7
  Xgate_2_118_0 vdd vss x_1[118] x_2[118] multi_finger_inv_7
  Xgate_2_119_0 vdd vss x_1[119] x_2[119] multi_finger_inv_7
  Xgate_2_120_0 vdd vss x_1[120] x_2[120] multi_finger_inv_7
  Xgate_2_121_0 vdd vss x_1[121] x_2[121] multi_finger_inv_7
  Xgate_2_122_0 vdd vss x_1[122] x_2[122] multi_finger_inv_7
  Xgate_2_123_0 vdd vss x_1[123] x_2[123] multi_finger_inv_7
  Xgate_2_124_0 vdd vss x_1[124] x_2[124] multi_finger_inv_7
  Xgate_2_125_0 vdd vss x_1[125] x_2[125] multi_finger_inv_7
  Xgate_2_126_0 vdd vss x_1[126] x_2[126] multi_finger_inv_7
  Xgate_2_127_0 vdd vss x_1[127] x_2[127] multi_finger_inv_7
  Xgate_3_0_0 vdd vss x_2[0] y_b[0] multi_finger_inv_8
  Xgate_3_1_0 vdd vss x_2[1] y_b[1] multi_finger_inv_8
  Xgate_3_2_0 vdd vss x_2[2] y_b[2] multi_finger_inv_8
  Xgate_3_3_0 vdd vss x_2[3] y_b[3] multi_finger_inv_8
  Xgate_3_4_0 vdd vss x_2[4] y_b[4] multi_finger_inv_8
  Xgate_3_5_0 vdd vss x_2[5] y_b[5] multi_finger_inv_8
  Xgate_3_6_0 vdd vss x_2[6] y_b[6] multi_finger_inv_8
  Xgate_3_7_0 vdd vss x_2[7] y_b[7] multi_finger_inv_8
  Xgate_3_8_0 vdd vss x_2[8] y_b[8] multi_finger_inv_8
  Xgate_3_9_0 vdd vss x_2[9] y_b[9] multi_finger_inv_8
  Xgate_3_10_0 vdd vss x_2[10] y_b[10] multi_finger_inv_8
  Xgate_3_11_0 vdd vss x_2[11] y_b[11] multi_finger_inv_8
  Xgate_3_12_0 vdd vss x_2[12] y_b[12] multi_finger_inv_8
  Xgate_3_13_0 vdd vss x_2[13] y_b[13] multi_finger_inv_8
  Xgate_3_14_0 vdd vss x_2[14] y_b[14] multi_finger_inv_8
  Xgate_3_15_0 vdd vss x_2[15] y_b[15] multi_finger_inv_8
  Xgate_3_16_0 vdd vss x_2[16] y_b[16] multi_finger_inv_8
  Xgate_3_17_0 vdd vss x_2[17] y_b[17] multi_finger_inv_8
  Xgate_3_18_0 vdd vss x_2[18] y_b[18] multi_finger_inv_8
  Xgate_3_19_0 vdd vss x_2[19] y_b[19] multi_finger_inv_8
  Xgate_3_20_0 vdd vss x_2[20] y_b[20] multi_finger_inv_8
  Xgate_3_21_0 vdd vss x_2[21] y_b[21] multi_finger_inv_8
  Xgate_3_22_0 vdd vss x_2[22] y_b[22] multi_finger_inv_8
  Xgate_3_23_0 vdd vss x_2[23] y_b[23] multi_finger_inv_8
  Xgate_3_24_0 vdd vss x_2[24] y_b[24] multi_finger_inv_8
  Xgate_3_25_0 vdd vss x_2[25] y_b[25] multi_finger_inv_8
  Xgate_3_26_0 vdd vss x_2[26] y_b[26] multi_finger_inv_8
  Xgate_3_27_0 vdd vss x_2[27] y_b[27] multi_finger_inv_8
  Xgate_3_28_0 vdd vss x_2[28] y_b[28] multi_finger_inv_8
  Xgate_3_29_0 vdd vss x_2[29] y_b[29] multi_finger_inv_8
  Xgate_3_30_0 vdd vss x_2[30] y_b[30] multi_finger_inv_8
  Xgate_3_31_0 vdd vss x_2[31] y_b[31] multi_finger_inv_8
  Xgate_3_32_0 vdd vss x_2[32] y_b[32] multi_finger_inv_8
  Xgate_3_33_0 vdd vss x_2[33] y_b[33] multi_finger_inv_8
  Xgate_3_34_0 vdd vss x_2[34] y_b[34] multi_finger_inv_8
  Xgate_3_35_0 vdd vss x_2[35] y_b[35] multi_finger_inv_8
  Xgate_3_36_0 vdd vss x_2[36] y_b[36] multi_finger_inv_8
  Xgate_3_37_0 vdd vss x_2[37] y_b[37] multi_finger_inv_8
  Xgate_3_38_0 vdd vss x_2[38] y_b[38] multi_finger_inv_8
  Xgate_3_39_0 vdd vss x_2[39] y_b[39] multi_finger_inv_8
  Xgate_3_40_0 vdd vss x_2[40] y_b[40] multi_finger_inv_8
  Xgate_3_41_0 vdd vss x_2[41] y_b[41] multi_finger_inv_8
  Xgate_3_42_0 vdd vss x_2[42] y_b[42] multi_finger_inv_8
  Xgate_3_43_0 vdd vss x_2[43] y_b[43] multi_finger_inv_8
  Xgate_3_44_0 vdd vss x_2[44] y_b[44] multi_finger_inv_8
  Xgate_3_45_0 vdd vss x_2[45] y_b[45] multi_finger_inv_8
  Xgate_3_46_0 vdd vss x_2[46] y_b[46] multi_finger_inv_8
  Xgate_3_47_0 vdd vss x_2[47] y_b[47] multi_finger_inv_8
  Xgate_3_48_0 vdd vss x_2[48] y_b[48] multi_finger_inv_8
  Xgate_3_49_0 vdd vss x_2[49] y_b[49] multi_finger_inv_8
  Xgate_3_50_0 vdd vss x_2[50] y_b[50] multi_finger_inv_8
  Xgate_3_51_0 vdd vss x_2[51] y_b[51] multi_finger_inv_8
  Xgate_3_52_0 vdd vss x_2[52] y_b[52] multi_finger_inv_8
  Xgate_3_53_0 vdd vss x_2[53] y_b[53] multi_finger_inv_8
  Xgate_3_54_0 vdd vss x_2[54] y_b[54] multi_finger_inv_8
  Xgate_3_55_0 vdd vss x_2[55] y_b[55] multi_finger_inv_8
  Xgate_3_56_0 vdd vss x_2[56] y_b[56] multi_finger_inv_8
  Xgate_3_57_0 vdd vss x_2[57] y_b[57] multi_finger_inv_8
  Xgate_3_58_0 vdd vss x_2[58] y_b[58] multi_finger_inv_8
  Xgate_3_59_0 vdd vss x_2[59] y_b[59] multi_finger_inv_8
  Xgate_3_60_0 vdd vss x_2[60] y_b[60] multi_finger_inv_8
  Xgate_3_61_0 vdd vss x_2[61] y_b[61] multi_finger_inv_8
  Xgate_3_62_0 vdd vss x_2[62] y_b[62] multi_finger_inv_8
  Xgate_3_63_0 vdd vss x_2[63] y_b[63] multi_finger_inv_8
  Xgate_3_64_0 vdd vss x_2[64] y_b[64] multi_finger_inv_8
  Xgate_3_65_0 vdd vss x_2[65] y_b[65] multi_finger_inv_8
  Xgate_3_66_0 vdd vss x_2[66] y_b[66] multi_finger_inv_8
  Xgate_3_67_0 vdd vss x_2[67] y_b[67] multi_finger_inv_8
  Xgate_3_68_0 vdd vss x_2[68] y_b[68] multi_finger_inv_8
  Xgate_3_69_0 vdd vss x_2[69] y_b[69] multi_finger_inv_8
  Xgate_3_70_0 vdd vss x_2[70] y_b[70] multi_finger_inv_8
  Xgate_3_71_0 vdd vss x_2[71] y_b[71] multi_finger_inv_8
  Xgate_3_72_0 vdd vss x_2[72] y_b[72] multi_finger_inv_8
  Xgate_3_73_0 vdd vss x_2[73] y_b[73] multi_finger_inv_8
  Xgate_3_74_0 vdd vss x_2[74] y_b[74] multi_finger_inv_8
  Xgate_3_75_0 vdd vss x_2[75] y_b[75] multi_finger_inv_8
  Xgate_3_76_0 vdd vss x_2[76] y_b[76] multi_finger_inv_8
  Xgate_3_77_0 vdd vss x_2[77] y_b[77] multi_finger_inv_8
  Xgate_3_78_0 vdd vss x_2[78] y_b[78] multi_finger_inv_8
  Xgate_3_79_0 vdd vss x_2[79] y_b[79] multi_finger_inv_8
  Xgate_3_80_0 vdd vss x_2[80] y_b[80] multi_finger_inv_8
  Xgate_3_81_0 vdd vss x_2[81] y_b[81] multi_finger_inv_8
  Xgate_3_82_0 vdd vss x_2[82] y_b[82] multi_finger_inv_8
  Xgate_3_83_0 vdd vss x_2[83] y_b[83] multi_finger_inv_8
  Xgate_3_84_0 vdd vss x_2[84] y_b[84] multi_finger_inv_8
  Xgate_3_85_0 vdd vss x_2[85] y_b[85] multi_finger_inv_8
  Xgate_3_86_0 vdd vss x_2[86] y_b[86] multi_finger_inv_8
  Xgate_3_87_0 vdd vss x_2[87] y_b[87] multi_finger_inv_8
  Xgate_3_88_0 vdd vss x_2[88] y_b[88] multi_finger_inv_8
  Xgate_3_89_0 vdd vss x_2[89] y_b[89] multi_finger_inv_8
  Xgate_3_90_0 vdd vss x_2[90] y_b[90] multi_finger_inv_8
  Xgate_3_91_0 vdd vss x_2[91] y_b[91] multi_finger_inv_8
  Xgate_3_92_0 vdd vss x_2[92] y_b[92] multi_finger_inv_8
  Xgate_3_93_0 vdd vss x_2[93] y_b[93] multi_finger_inv_8
  Xgate_3_94_0 vdd vss x_2[94] y_b[94] multi_finger_inv_8
  Xgate_3_95_0 vdd vss x_2[95] y_b[95] multi_finger_inv_8
  Xgate_3_96_0 vdd vss x_2[96] y_b[96] multi_finger_inv_8
  Xgate_3_97_0 vdd vss x_2[97] y_b[97] multi_finger_inv_8
  Xgate_3_98_0 vdd vss x_2[98] y_b[98] multi_finger_inv_8
  Xgate_3_99_0 vdd vss x_2[99] y_b[99] multi_finger_inv_8
  Xgate_3_100_0 vdd vss x_2[100] y_b[100] multi_finger_inv_8
  Xgate_3_101_0 vdd vss x_2[101] y_b[101] multi_finger_inv_8
  Xgate_3_102_0 vdd vss x_2[102] y_b[102] multi_finger_inv_8
  Xgate_3_103_0 vdd vss x_2[103] y_b[103] multi_finger_inv_8
  Xgate_3_104_0 vdd vss x_2[104] y_b[104] multi_finger_inv_8
  Xgate_3_105_0 vdd vss x_2[105] y_b[105] multi_finger_inv_8
  Xgate_3_106_0 vdd vss x_2[106] y_b[106] multi_finger_inv_8
  Xgate_3_107_0 vdd vss x_2[107] y_b[107] multi_finger_inv_8
  Xgate_3_108_0 vdd vss x_2[108] y_b[108] multi_finger_inv_8
  Xgate_3_109_0 vdd vss x_2[109] y_b[109] multi_finger_inv_8
  Xgate_3_110_0 vdd vss x_2[110] y_b[110] multi_finger_inv_8
  Xgate_3_111_0 vdd vss x_2[111] y_b[111] multi_finger_inv_8
  Xgate_3_112_0 vdd vss x_2[112] y_b[112] multi_finger_inv_8
  Xgate_3_113_0 vdd vss x_2[113] y_b[113] multi_finger_inv_8
  Xgate_3_114_0 vdd vss x_2[114] y_b[114] multi_finger_inv_8
  Xgate_3_115_0 vdd vss x_2[115] y_b[115] multi_finger_inv_8
  Xgate_3_116_0 vdd vss x_2[116] y_b[116] multi_finger_inv_8
  Xgate_3_117_0 vdd vss x_2[117] y_b[117] multi_finger_inv_8
  Xgate_3_118_0 vdd vss x_2[118] y_b[118] multi_finger_inv_8
  Xgate_3_119_0 vdd vss x_2[119] y_b[119] multi_finger_inv_8
  Xgate_3_120_0 vdd vss x_2[120] y_b[120] multi_finger_inv_8
  Xgate_3_121_0 vdd vss x_2[121] y_b[121] multi_finger_inv_8
  Xgate_3_122_0 vdd vss x_2[122] y_b[122] multi_finger_inv_8
  Xgate_3_123_0 vdd vss x_2[123] y_b[123] multi_finger_inv_8
  Xgate_3_124_0 vdd vss x_2[124] y_b[124] multi_finger_inv_8
  Xgate_3_125_0 vdd vss x_2[125] y_b[125] multi_finger_inv_8
  Xgate_3_126_0 vdd vss x_2[126] y_b[126] multi_finger_inv_8
  Xgate_3_127_0 vdd vss x_2[127] y_b[127] multi_finger_inv_8
  Xgate_4_0_0 vdd vss y_b[0] y[0] multi_finger_inv_9
  Xgate_4_1_0 vdd vss y_b[1] y[1] multi_finger_inv_9
  Xgate_4_2_0 vdd vss y_b[2] y[2] multi_finger_inv_9
  Xgate_4_3_0 vdd vss y_b[3] y[3] multi_finger_inv_9
  Xgate_4_4_0 vdd vss y_b[4] y[4] multi_finger_inv_9
  Xgate_4_5_0 vdd vss y_b[5] y[5] multi_finger_inv_9
  Xgate_4_6_0 vdd vss y_b[6] y[6] multi_finger_inv_9
  Xgate_4_7_0 vdd vss y_b[7] y[7] multi_finger_inv_9
  Xgate_4_8_0 vdd vss y_b[8] y[8] multi_finger_inv_9
  Xgate_4_9_0 vdd vss y_b[9] y[9] multi_finger_inv_9
  Xgate_4_10_0 vdd vss y_b[10] y[10] multi_finger_inv_9
  Xgate_4_11_0 vdd vss y_b[11] y[11] multi_finger_inv_9
  Xgate_4_12_0 vdd vss y_b[12] y[12] multi_finger_inv_9
  Xgate_4_13_0 vdd vss y_b[13] y[13] multi_finger_inv_9
  Xgate_4_14_0 vdd vss y_b[14] y[14] multi_finger_inv_9
  Xgate_4_15_0 vdd vss y_b[15] y[15] multi_finger_inv_9
  Xgate_4_16_0 vdd vss y_b[16] y[16] multi_finger_inv_9
  Xgate_4_17_0 vdd vss y_b[17] y[17] multi_finger_inv_9
  Xgate_4_18_0 vdd vss y_b[18] y[18] multi_finger_inv_9
  Xgate_4_19_0 vdd vss y_b[19] y[19] multi_finger_inv_9
  Xgate_4_20_0 vdd vss y_b[20] y[20] multi_finger_inv_9
  Xgate_4_21_0 vdd vss y_b[21] y[21] multi_finger_inv_9
  Xgate_4_22_0 vdd vss y_b[22] y[22] multi_finger_inv_9
  Xgate_4_23_0 vdd vss y_b[23] y[23] multi_finger_inv_9
  Xgate_4_24_0 vdd vss y_b[24] y[24] multi_finger_inv_9
  Xgate_4_25_0 vdd vss y_b[25] y[25] multi_finger_inv_9
  Xgate_4_26_0 vdd vss y_b[26] y[26] multi_finger_inv_9
  Xgate_4_27_0 vdd vss y_b[27] y[27] multi_finger_inv_9
  Xgate_4_28_0 vdd vss y_b[28] y[28] multi_finger_inv_9
  Xgate_4_29_0 vdd vss y_b[29] y[29] multi_finger_inv_9
  Xgate_4_30_0 vdd vss y_b[30] y[30] multi_finger_inv_9
  Xgate_4_31_0 vdd vss y_b[31] y[31] multi_finger_inv_9
  Xgate_4_32_0 vdd vss y_b[32] y[32] multi_finger_inv_9
  Xgate_4_33_0 vdd vss y_b[33] y[33] multi_finger_inv_9
  Xgate_4_34_0 vdd vss y_b[34] y[34] multi_finger_inv_9
  Xgate_4_35_0 vdd vss y_b[35] y[35] multi_finger_inv_9
  Xgate_4_36_0 vdd vss y_b[36] y[36] multi_finger_inv_9
  Xgate_4_37_0 vdd vss y_b[37] y[37] multi_finger_inv_9
  Xgate_4_38_0 vdd vss y_b[38] y[38] multi_finger_inv_9
  Xgate_4_39_0 vdd vss y_b[39] y[39] multi_finger_inv_9
  Xgate_4_40_0 vdd vss y_b[40] y[40] multi_finger_inv_9
  Xgate_4_41_0 vdd vss y_b[41] y[41] multi_finger_inv_9
  Xgate_4_42_0 vdd vss y_b[42] y[42] multi_finger_inv_9
  Xgate_4_43_0 vdd vss y_b[43] y[43] multi_finger_inv_9
  Xgate_4_44_0 vdd vss y_b[44] y[44] multi_finger_inv_9
  Xgate_4_45_0 vdd vss y_b[45] y[45] multi_finger_inv_9
  Xgate_4_46_0 vdd vss y_b[46] y[46] multi_finger_inv_9
  Xgate_4_47_0 vdd vss y_b[47] y[47] multi_finger_inv_9
  Xgate_4_48_0 vdd vss y_b[48] y[48] multi_finger_inv_9
  Xgate_4_49_0 vdd vss y_b[49] y[49] multi_finger_inv_9
  Xgate_4_50_0 vdd vss y_b[50] y[50] multi_finger_inv_9
  Xgate_4_51_0 vdd vss y_b[51] y[51] multi_finger_inv_9
  Xgate_4_52_0 vdd vss y_b[52] y[52] multi_finger_inv_9
  Xgate_4_53_0 vdd vss y_b[53] y[53] multi_finger_inv_9
  Xgate_4_54_0 vdd vss y_b[54] y[54] multi_finger_inv_9
  Xgate_4_55_0 vdd vss y_b[55] y[55] multi_finger_inv_9
  Xgate_4_56_0 vdd vss y_b[56] y[56] multi_finger_inv_9
  Xgate_4_57_0 vdd vss y_b[57] y[57] multi_finger_inv_9
  Xgate_4_58_0 vdd vss y_b[58] y[58] multi_finger_inv_9
  Xgate_4_59_0 vdd vss y_b[59] y[59] multi_finger_inv_9
  Xgate_4_60_0 vdd vss y_b[60] y[60] multi_finger_inv_9
  Xgate_4_61_0 vdd vss y_b[61] y[61] multi_finger_inv_9
  Xgate_4_62_0 vdd vss y_b[62] y[62] multi_finger_inv_9
  Xgate_4_63_0 vdd vss y_b[63] y[63] multi_finger_inv_9
  Xgate_4_64_0 vdd vss y_b[64] y[64] multi_finger_inv_9
  Xgate_4_65_0 vdd vss y_b[65] y[65] multi_finger_inv_9
  Xgate_4_66_0 vdd vss y_b[66] y[66] multi_finger_inv_9
  Xgate_4_67_0 vdd vss y_b[67] y[67] multi_finger_inv_9
  Xgate_4_68_0 vdd vss y_b[68] y[68] multi_finger_inv_9
  Xgate_4_69_0 vdd vss y_b[69] y[69] multi_finger_inv_9
  Xgate_4_70_0 vdd vss y_b[70] y[70] multi_finger_inv_9
  Xgate_4_71_0 vdd vss y_b[71] y[71] multi_finger_inv_9
  Xgate_4_72_0 vdd vss y_b[72] y[72] multi_finger_inv_9
  Xgate_4_73_0 vdd vss y_b[73] y[73] multi_finger_inv_9
  Xgate_4_74_0 vdd vss y_b[74] y[74] multi_finger_inv_9
  Xgate_4_75_0 vdd vss y_b[75] y[75] multi_finger_inv_9
  Xgate_4_76_0 vdd vss y_b[76] y[76] multi_finger_inv_9
  Xgate_4_77_0 vdd vss y_b[77] y[77] multi_finger_inv_9
  Xgate_4_78_0 vdd vss y_b[78] y[78] multi_finger_inv_9
  Xgate_4_79_0 vdd vss y_b[79] y[79] multi_finger_inv_9
  Xgate_4_80_0 vdd vss y_b[80] y[80] multi_finger_inv_9
  Xgate_4_81_0 vdd vss y_b[81] y[81] multi_finger_inv_9
  Xgate_4_82_0 vdd vss y_b[82] y[82] multi_finger_inv_9
  Xgate_4_83_0 vdd vss y_b[83] y[83] multi_finger_inv_9
  Xgate_4_84_0 vdd vss y_b[84] y[84] multi_finger_inv_9
  Xgate_4_85_0 vdd vss y_b[85] y[85] multi_finger_inv_9
  Xgate_4_86_0 vdd vss y_b[86] y[86] multi_finger_inv_9
  Xgate_4_87_0 vdd vss y_b[87] y[87] multi_finger_inv_9
  Xgate_4_88_0 vdd vss y_b[88] y[88] multi_finger_inv_9
  Xgate_4_89_0 vdd vss y_b[89] y[89] multi_finger_inv_9
  Xgate_4_90_0 vdd vss y_b[90] y[90] multi_finger_inv_9
  Xgate_4_91_0 vdd vss y_b[91] y[91] multi_finger_inv_9
  Xgate_4_92_0 vdd vss y_b[92] y[92] multi_finger_inv_9
  Xgate_4_93_0 vdd vss y_b[93] y[93] multi_finger_inv_9
  Xgate_4_94_0 vdd vss y_b[94] y[94] multi_finger_inv_9
  Xgate_4_95_0 vdd vss y_b[95] y[95] multi_finger_inv_9
  Xgate_4_96_0 vdd vss y_b[96] y[96] multi_finger_inv_9
  Xgate_4_97_0 vdd vss y_b[97] y[97] multi_finger_inv_9
  Xgate_4_98_0 vdd vss y_b[98] y[98] multi_finger_inv_9
  Xgate_4_99_0 vdd vss y_b[99] y[99] multi_finger_inv_9
  Xgate_4_100_0 vdd vss y_b[100] y[100] multi_finger_inv_9
  Xgate_4_101_0 vdd vss y_b[101] y[101] multi_finger_inv_9
  Xgate_4_102_0 vdd vss y_b[102] y[102] multi_finger_inv_9
  Xgate_4_103_0 vdd vss y_b[103] y[103] multi_finger_inv_9
  Xgate_4_104_0 vdd vss y_b[104] y[104] multi_finger_inv_9
  Xgate_4_105_0 vdd vss y_b[105] y[105] multi_finger_inv_9
  Xgate_4_106_0 vdd vss y_b[106] y[106] multi_finger_inv_9
  Xgate_4_107_0 vdd vss y_b[107] y[107] multi_finger_inv_9
  Xgate_4_108_0 vdd vss y_b[108] y[108] multi_finger_inv_9
  Xgate_4_109_0 vdd vss y_b[109] y[109] multi_finger_inv_9
  Xgate_4_110_0 vdd vss y_b[110] y[110] multi_finger_inv_9
  Xgate_4_111_0 vdd vss y_b[111] y[111] multi_finger_inv_9
  Xgate_4_112_0 vdd vss y_b[112] y[112] multi_finger_inv_9
  Xgate_4_113_0 vdd vss y_b[113] y[113] multi_finger_inv_9
  Xgate_4_114_0 vdd vss y_b[114] y[114] multi_finger_inv_9
  Xgate_4_115_0 vdd vss y_b[115] y[115] multi_finger_inv_9
  Xgate_4_116_0 vdd vss y_b[116] y[116] multi_finger_inv_9
  Xgate_4_117_0 vdd vss y_b[117] y[117] multi_finger_inv_9
  Xgate_4_118_0 vdd vss y_b[118] y[118] multi_finger_inv_9
  Xgate_4_119_0 vdd vss y_b[119] y[119] multi_finger_inv_9
  Xgate_4_120_0 vdd vss y_b[120] y[120] multi_finger_inv_9
  Xgate_4_121_0 vdd vss y_b[121] y[121] multi_finger_inv_9
  Xgate_4_122_0 vdd vss y_b[122] y[122] multi_finger_inv_9
  Xgate_4_123_0 vdd vss y_b[123] y[123] multi_finger_inv_9
  Xgate_4_124_0 vdd vss y_b[124] y[124] multi_finger_inv_9
  Xgate_4_125_0 vdd vss y_b[125] y[125] multi_finger_inv_9
  Xgate_4_126_0 vdd vss y_b[126] y[126] multi_finger_inv_9
  Xgate_4_127_0 vdd vss y_b[127] y[127] multi_finger_inv_9

.ENDS decoder_stage_5

.SUBCKT decoder vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y[12] y[13] y[14] y[15] y[16] y[17] y[18] y[19] y[20] y[21] y[22] y[23] y[24] y[25] y[26] y[27] y[28] y[29] y[30] y[31] y[32] y[33] y[34] y[35] y[36] y[37] y[38] y[39] y[40] y[41] y[42] y[43] y[44] y[45] y[46] y[47] y[48] y[49] y[50] y[51] y[52] y[53] y[54] y[55] y[56] y[57] y[58] y[59] y[60] y[61] y[62] y[63] y[64] y[65] y[66] y[67] y[68] y[69] y[70] y[71] y[72] y[73] y[74] y[75] y[76] y[77] y[78] y[79] y[80] y[81] y[82] y[83] y[84] y[85] y[86] y[87] y[88] y[89] y[90] y[91] y[92] y[93] y[94] y[95] y[96] y[97] y[98] y[99] y[100] y[101] y[102] y[103] y[104] y[105] y[106] y[107] y[108] y[109] y[110] y[111] y[112] y[113] y[114] y[115] y[116] y[117] y[118] y[119] y[120] y[121] y[122] y[123] y[124] y[125] y[126] y[127] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] y_b[12] y_b[13] y_b[14] y_b[15] y_b[16] y_b[17] y_b[18] y_b[19] y_b[20] y_b[21] y_b[22] y_b[23] y_b[24] y_b[25] y_b[26] y_b[27] y_b[28] y_b[29] y_b[30] y_b[31] y_b[32] y_b[33] y_b[34] y_b[35] y_b[36] y_b[37] y_b[38] y_b[39] y_b[40] y_b[41] y_b[42] y_b[43] y_b[44] y_b[45] y_b[46] y_b[47] y_b[48] y_b[49] y_b[50] y_b[51] y_b[52] y_b[53] y_b[54] y_b[55] y_b[56] y_b[57] y_b[58] y_b[59] y_b[60] y_b[61] y_b[62] y_b[63] y_b[64] y_b[65] y_b[66] y_b[67] y_b[68] y_b[69] y_b[70] y_b[71] y_b[72] y_b[73] y_b[74] y_b[75] y_b[76] y_b[77] y_b[78] y_b[79] y_b[80] y_b[81] y_b[82] y_b[83] y_b[84] y_b[85] y_b[86] y_b[87] y_b[88] y_b[89] y_b[90] y_b[91] y_b[92] y_b[93] y_b[94] y_b[95] y_b[96] y_b[97] y_b[98] y_b[99] y_b[100] y_b[101] y_b[102] y_b[103] y_b[104] y_b[105] y_b[106] y_b[107] y_b[108] y_b[109] y_b[110] y_b[111] y_b[112] y_b[113] y_b[114] y_b[115] y_b[116] y_b[117] y_b[118] y_b[119] y_b[120] y_b[121] y_b[122] y_b[123] y_b[124] y_b[125] y_b[126] y_b[127] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 predecode_2_0 predecode_2_1 predecode_3_0 predecode_3_1 predecode_4_0 predecode_4_1 predecode_5_0 predecode_5_1 predecode_6_0 predecode_6_1

  X0 vdd vss child_conn_0[0] child_conn_0[1] child_conn_0[2] child_conn_0[3] child_conn_0[4] child_conn_0[5] child_conn_0[6] child_conn_0[7] child_conn_0[8] child_conn_0[9] child_conn_0[10] child_conn_0[11] child_conn_0[12] child_conn_0[13] child_conn_0[14] child_conn_0[15] child_noconn_0[0] child_noconn_0[1] child_noconn_0[2] child_noconn_0[3] child_noconn_0[4] child_noconn_0[5] child_noconn_0[6] child_noconn_0[7] child_noconn_0[8] child_noconn_0[9] child_noconn_0[10] child_noconn_0[11] child_noconn_0[12] child_noconn_0[13] child_noconn_0[14] child_noconn_0[15] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 predecode_2_0 predecode_2_1 predecode_3_0 predecode_3_1 decoder_2
  X0_1 vdd vss child_conn_1[0] child_conn_1[1] child_conn_1[2] child_conn_1[3] child_conn_1[4] child_conn_1[5] child_conn_1[6] child_conn_1[7] child_noconn_1[0] child_noconn_1[1] child_noconn_1[2] child_noconn_1[3] child_noconn_1[4] child_noconn_1[5] child_noconn_1[6] child_noconn_1[7] predecode_4_0 predecode_4_1 predecode_5_0 predecode_5_1 predecode_6_0 predecode_6_1 decoder_3
  X0_2 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y[12] y[13] y[14] y[15] y[16] y[17] y[18] y[19] y[20] y[21] y[22] y[23] y[24] y[25] y[26] y[27] y[28] y[29] y[30] y[31] y[32] y[33] y[34] y[35] y[36] y[37] y[38] y[39] y[40] y[41] y[42] y[43] y[44] y[45] y[46] y[47] y[48] y[49] y[50] y[51] y[52] y[53] y[54] y[55] y[56] y[57] y[58] y[59] y[60] y[61] y[62] y[63] y[64] y[65] y[66] y[67] y[68] y[69] y[70] y[71] y[72] y[73] y[74] y[75] y[76] y[77] y[78] y[79] y[80] y[81] y[82] y[83] y[84] y[85] y[86] y[87] y[88] y[89] y[90] y[91] y[92] y[93] y[94] y[95] y[96] y[97] y[98] y[99] y[100] y[101] y[102] y[103] y[104] y[105] y[106] y[107] y[108] y[109] y[110] y[111] y[112] y[113] y[114] y[115] y[116] y[117] y[118] y[119] y[120] y[121] y[122] y[123] y[124] y[125] y[126] y[127] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] y_b[12] y_b[13] y_b[14] y_b[15] y_b[16] y_b[17] y_b[18] y_b[19] y_b[20] y_b[21] y_b[22] y_b[23] y_b[24] y_b[25] y_b[26] y_b[27] y_b[28] y_b[29] y_b[30] y_b[31] y_b[32] y_b[33] y_b[34] y_b[35] y_b[36] y_b[37] y_b[38] y_b[39] y_b[40] y_b[41] y_b[42] y_b[43] y_b[44] y_b[45] y_b[46] y_b[47] y_b[48] y_b[49] y_b[50] y_b[51] y_b[52] y_b[53] y_b[54] y_b[55] y_b[56] y_b[57] y_b[58] y_b[59] y_b[60] y_b[61] y_b[62] y_b[63] y_b[64] y_b[65] y_b[66] y_b[67] y_b[68] y_b[69] y_b[70] y_b[71] y_b[72] y_b[73] y_b[74] y_b[75] y_b[76] y_b[77] y_b[78] y_b[79] y_b[80] y_b[81] y_b[82] y_b[83] y_b[84] y_b[85] y_b[86] y_b[87] y_b[88] y_b[89] y_b[90] y_b[91] y_b[92] y_b[93] y_b[94] y_b[95] y_b[96] y_b[97] y_b[98] y_b[99] y_b[100] y_b[101] y_b[102] y_b[103] y_b[104] y_b[105] y_b[106] y_b[107] y_b[108] y_b[109] y_b[110] y_b[111] y_b[112] y_b[113] y_b[114] y_b[115] y_b[116] y_b[117] y_b[118] y_b[119] y_b[120] y_b[121] y_b[122] y_b[123] y_b[124] y_b[125] y_b[126] y_b[127] child_conn_0[0] child_conn_0[1] child_conn_0[2] child_conn_0[3] child_conn_0[4] child_conn_0[5] child_conn_0[6] child_conn_0[7] child_conn_0[8] child_conn_0[9] child_conn_0[10] child_conn_0[11] child_conn_0[12] child_conn_0[13] child_conn_0[14] child_conn_0[15] child_conn_1[0] child_conn_1[1] child_conn_1[2] child_conn_1[3] child_conn_1[4] child_conn_1[5] child_conn_1[6] child_conn_1[7] decoder_stage_5

.ENDS decoder

.SUBCKT multi_finger_inv_11 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_11

.SUBCKT multi_finger_inv_12 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN7 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_12

.SUBCKT decoder_stage_6 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 predecode_2_0 predecode_2_1

  Xgate_0_0_0 vdd vss predecode_0_0 predecode_1_0 predecode_2_0 x_0[0] nand3
  Xgate_0_1_0 vdd vss predecode_0_1 predecode_1_0 predecode_2_0 x_0[1] nand3
  Xgate_0_2_0 vdd vss predecode_0_0 predecode_1_1 predecode_2_0 x_0[2] nand3
  Xgate_0_3_0 vdd vss predecode_0_1 predecode_1_1 predecode_2_0 x_0[3] nand3
  Xgate_0_4_0 vdd vss predecode_0_0 predecode_1_0 predecode_2_1 x_0[4] nand3
  Xgate_0_5_0 vdd vss predecode_0_1 predecode_1_0 predecode_2_1 x_0[5] nand3
  Xgate_0_6_0 vdd vss predecode_0_0 predecode_1_1 predecode_2_1 x_0[6] nand3
  Xgate_0_7_0 vdd vss predecode_0_1 predecode_1_1 predecode_2_1 x_0[7] nand3
  Xgate_1_0_0 vdd vss x_0[0] x_1[0] multi_finger_inv_10
  Xgate_1_1_0 vdd vss x_0[1] x_1[1] multi_finger_inv_10
  Xgate_1_2_0 vdd vss x_0[2] x_1[2] multi_finger_inv_10
  Xgate_1_3_0 vdd vss x_0[3] x_1[3] multi_finger_inv_10
  Xgate_1_4_0 vdd vss x_0[4] x_1[4] multi_finger_inv_10
  Xgate_1_5_0 vdd vss x_0[5] x_1[5] multi_finger_inv_10
  Xgate_1_6_0 vdd vss x_0[6] x_1[6] multi_finger_inv_10
  Xgate_1_7_0 vdd vss x_0[7] x_1[7] multi_finger_inv_10
  Xgate_2_0_0 vdd vss x_1[0] y_b[0] multi_finger_inv_11
  Xgate_2_0_1 vdd vss x_1[0] y_b[0] multi_finger_inv_11
  Xgate_2_0_2 vdd vss x_1[0] y_b[0] multi_finger_inv_11
  Xgate_2_1_0 vdd vss x_1[1] y_b[1] multi_finger_inv_11
  Xgate_2_1_1 vdd vss x_1[1] y_b[1] multi_finger_inv_11
  Xgate_2_1_2 vdd vss x_1[1] y_b[1] multi_finger_inv_11
  Xgate_2_2_0 vdd vss x_1[2] y_b[2] multi_finger_inv_11
  Xgate_2_2_1 vdd vss x_1[2] y_b[2] multi_finger_inv_11
  Xgate_2_2_2 vdd vss x_1[2] y_b[2] multi_finger_inv_11
  Xgate_2_3_0 vdd vss x_1[3] y_b[3] multi_finger_inv_11
  Xgate_2_3_1 vdd vss x_1[3] y_b[3] multi_finger_inv_11
  Xgate_2_3_2 vdd vss x_1[3] y_b[3] multi_finger_inv_11
  Xgate_2_4_0 vdd vss x_1[4] y_b[4] multi_finger_inv_11
  Xgate_2_4_1 vdd vss x_1[4] y_b[4] multi_finger_inv_11
  Xgate_2_4_2 vdd vss x_1[4] y_b[4] multi_finger_inv_11
  Xgate_2_5_0 vdd vss x_1[5] y_b[5] multi_finger_inv_11
  Xgate_2_5_1 vdd vss x_1[5] y_b[5] multi_finger_inv_11
  Xgate_2_5_2 vdd vss x_1[5] y_b[5] multi_finger_inv_11
  Xgate_2_6_0 vdd vss x_1[6] y_b[6] multi_finger_inv_11
  Xgate_2_6_1 vdd vss x_1[6] y_b[6] multi_finger_inv_11
  Xgate_2_6_2 vdd vss x_1[6] y_b[6] multi_finger_inv_11
  Xgate_2_7_0 vdd vss x_1[7] y_b[7] multi_finger_inv_11
  Xgate_2_7_1 vdd vss x_1[7] y_b[7] multi_finger_inv_11
  Xgate_2_7_2 vdd vss x_1[7] y_b[7] multi_finger_inv_11
  Xgate_3_0_0 vdd vss y_b[0] y[0] multi_finger_inv_12
  Xgate_3_0_1 vdd vss y_b[0] y[0] multi_finger_inv_12
  Xgate_3_0_2 vdd vss y_b[0] y[0] multi_finger_inv_12
  Xgate_3_1_0 vdd vss y_b[1] y[1] multi_finger_inv_12
  Xgate_3_1_1 vdd vss y_b[1] y[1] multi_finger_inv_12
  Xgate_3_1_2 vdd vss y_b[1] y[1] multi_finger_inv_12
  Xgate_3_2_0 vdd vss y_b[2] y[2] multi_finger_inv_12
  Xgate_3_2_1 vdd vss y_b[2] y[2] multi_finger_inv_12
  Xgate_3_2_2 vdd vss y_b[2] y[2] multi_finger_inv_12
  Xgate_3_3_0 vdd vss y_b[3] y[3] multi_finger_inv_12
  Xgate_3_3_1 vdd vss y_b[3] y[3] multi_finger_inv_12
  Xgate_3_3_2 vdd vss y_b[3] y[3] multi_finger_inv_12
  Xgate_3_4_0 vdd vss y_b[4] y[4] multi_finger_inv_12
  Xgate_3_4_1 vdd vss y_b[4] y[4] multi_finger_inv_12
  Xgate_3_4_2 vdd vss y_b[4] y[4] multi_finger_inv_12
  Xgate_3_5_0 vdd vss y_b[5] y[5] multi_finger_inv_12
  Xgate_3_5_1 vdd vss y_b[5] y[5] multi_finger_inv_12
  Xgate_3_5_2 vdd vss y_b[5] y[5] multi_finger_inv_12
  Xgate_3_6_0 vdd vss y_b[6] y[6] multi_finger_inv_12
  Xgate_3_6_1 vdd vss y_b[6] y[6] multi_finger_inv_12
  Xgate_3_6_2 vdd vss y_b[6] y[6] multi_finger_inv_12
  Xgate_3_7_0 vdd vss y_b[7] y[7] multi_finger_inv_12
  Xgate_3_7_1 vdd vss y_b[7] y[7] multi_finger_inv_12
  Xgate_3_7_2 vdd vss y_b[7] y[7] multi_finger_inv_12

.ENDS decoder_stage_6

.SUBCKT decoder_1 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 predecode_2_0 predecode_2_1

  X0 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 predecode_2_0 predecode_2_1 decoder_stage_6

.ENDS decoder_1

.SUBCKT sky130_fd_sc_hs__inv_16 A VGND VNB VPB VPWR Y

  X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X5 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X7 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X11 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X13 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X14 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X15 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X16 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X17 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X18 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X19 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X20 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X21 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X22 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X23 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X24 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X25 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X26 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X27 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X28 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X30 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X31 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120


.ENDS sky130_fd_sc_hs__inv_16

.SUBCKT sky130_fd_sc_hs__inv_16_wrapper A VGND VNB VPB VPWR Y

  X0 A VGND VNB VPB VPWR Y sky130_fd_sc_hs__inv_16

.ENDS sky130_fd_sc_hs__inv_16_wrapper

.SUBCKT inv_chain_12 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sky130_fd_sc_hs__inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd x[2] sky130_fd_sc_hs__inv_2_wrapper
  Xinv3 x[2] vss vss vdd vdd x[3] sky130_fd_sc_hs__inv_2_wrapper
  Xinv4 x[3] vss vss vdd vdd x[4] sky130_fd_sc_hs__inv_2_wrapper
  Xinv5 x[4] vss vss vdd vdd x[5] sky130_fd_sc_hs__inv_2_wrapper
  Xinv6 x[5] vss vss vdd vdd x[6] sky130_fd_sc_hs__inv_2_wrapper
  Xinv7 x[6] vss vss vdd vdd x[7] sky130_fd_sc_hs__inv_2_wrapper
  Xinv8 x[7] vss vss vdd vdd x[8] sky130_fd_sc_hs__inv_2_wrapper
  Xinv9 x[8] vss vss vdd vdd x[9] sky130_fd_sc_hs__inv_2_wrapper
  Xinv10 x[9] vss vss vdd vdd x[10] sky130_fd_sc_hs__inv_2_wrapper
  Xinv11 x[10] vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_12

.SUBCKT sky130_fd_sc_hs__and2_2 A B VGND VNB VPB VPWR X

  X0 a_31_74# B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X1 X a_31_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X2 X a_31_74# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 a_118_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X4 a_31_74# A a_118_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X5 VPWR A a_31_74# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X6 VPWR a_31_74# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X7 VGND a_31_74# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__and2_2

.SUBCKT sky130_fd_sc_hs__and2_2_wrapper A B VGND VNB VPB VPWR X

  X0 A B VGND VNB VPB VPWR X sky130_fd_sc_hs__and2_2

.ENDS sky130_fd_sc_hs__and2_2_wrapper

.SUBCKT inv_chain_9 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sky130_fd_sc_hs__inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd x[2] sky130_fd_sc_hs__inv_2_wrapper
  Xinv3 x[2] vss vss vdd vdd x[3] sky130_fd_sc_hs__inv_2_wrapper
  Xinv4 x[3] vss vss vdd vdd x[4] sky130_fd_sc_hs__inv_2_wrapper
  Xinv5 x[4] vss vss vdd vdd x[5] sky130_fd_sc_hs__inv_2_wrapper
  Xinv6 x[5] vss vss vdd vdd x[6] sky130_fd_sc_hs__inv_2_wrapper
  Xinv7 x[6] vss vss vdd vdd x[7] sky130_fd_sc_hs__inv_2_wrapper
  Xinv8 x[7] vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_9

.SUBCKT edge_detector din dout vdd vss

  Xdelay_chain din delayed vdd vss inv_chain_9
  Xand din delayed vss vss vdd vdd dout sky130_fd_sc_hs__and2_4_wrapper

.ENDS edge_detector

.SUBCKT inv_chain_15 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sky130_fd_sc_hs__inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd x[2] sky130_fd_sc_hs__inv_2_wrapper
  Xinv3 x[2] vss vss vdd vdd x[3] sky130_fd_sc_hs__inv_2_wrapper
  Xinv4 x[3] vss vss vdd vdd x[4] sky130_fd_sc_hs__inv_2_wrapper
  Xinv5 x[4] vss vss vdd vdd x[5] sky130_fd_sc_hs__inv_2_wrapper
  Xinv6 x[5] vss vss vdd vdd x[6] sky130_fd_sc_hs__inv_2_wrapper
  Xinv7 x[6] vss vss vdd vdd x[7] sky130_fd_sc_hs__inv_2_wrapper
  Xinv8 x[7] vss vss vdd vdd x[8] sky130_fd_sc_hs__inv_2_wrapper
  Xinv9 x[8] vss vss vdd vdd x[9] sky130_fd_sc_hs__inv_2_wrapper
  Xinv10 x[9] vss vss vdd vdd x[10] sky130_fd_sc_hs__inv_2_wrapper
  Xinv11 x[10] vss vss vdd vdd x[11] sky130_fd_sc_hs__inv_2_wrapper
  Xinv12 x[11] vss vss vdd vdd x[12] sky130_fd_sc_hs__inv_2_wrapper
  Xinv13 x[12] vss vss vdd vdd x[13] sky130_fd_sc_hs__inv_2_wrapper
  Xinv14 x[13] vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_15

.SUBCKT sramgen_svt_inv_2_wrapper A VGND VNB VPB VPWR Y

  X0 A VGND VNB VPB VPWR Y sramgen_svt_inv_2

.ENDS sramgen_svt_inv_2_wrapper

.SUBCKT sramgen_svt_inv_4 A VGND VNB VPB VPWR Y

  X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740

  X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740

  X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740

  X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740


.ENDS sramgen_svt_inv_4

.SUBCKT sramgen_svt_inv_4_wrapper A VGND VNB VPB VPWR Y

  X0 A VGND VNB VPB VPWR Y sramgen_svt_inv_4

.ENDS sramgen_svt_inv_4_wrapper

.SUBCKT svt_inv_chain_30 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sramgen_svt_inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sramgen_svt_inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd x[2] sramgen_svt_inv_2_wrapper
  Xinv3 x[2] vss vss vdd vdd x[3] sramgen_svt_inv_2_wrapper
  Xinv4 x[3] vss vss vdd vdd x[4] sramgen_svt_inv_2_wrapper
  Xinv5 x[4] vss vss vdd vdd x[5] sramgen_svt_inv_2_wrapper
  Xinv6 x[5] vss vss vdd vdd x[6] sramgen_svt_inv_2_wrapper
  Xinv7 x[6] vss vss vdd vdd x[7] sramgen_svt_inv_2_wrapper
  Xinv8 x[7] vss vss vdd vdd x[8] sramgen_svt_inv_2_wrapper
  Xinv9 x[8] vss vss vdd vdd x[9] sramgen_svt_inv_2_wrapper
  Xinv10 x[9] vss vss vdd vdd x[10] sramgen_svt_inv_2_wrapper
  Xinv11 x[10] vss vss vdd vdd x[11] sramgen_svt_inv_2_wrapper
  Xinv12 x[11] vss vss vdd vdd x[12] sramgen_svt_inv_2_wrapper
  Xinv13 x[12] vss vss vdd vdd x[13] sramgen_svt_inv_2_wrapper
  Xinv14 x[13] vss vss vdd vdd x[14] sramgen_svt_inv_2_wrapper
  Xinv15 x[14] vss vss vdd vdd x[15] sramgen_svt_inv_2_wrapper
  Xinv16 x[15] vss vss vdd vdd x[16] sramgen_svt_inv_2_wrapper
  Xinv17 x[16] vss vss vdd vdd x[17] sramgen_svt_inv_2_wrapper
  Xinv18 x[17] vss vss vdd vdd x[18] sramgen_svt_inv_2_wrapper
  Xinv19 x[18] vss vss vdd vdd x[19] sramgen_svt_inv_2_wrapper
  Xinv20 x[19] vss vss vdd vdd x[20] sramgen_svt_inv_2_wrapper
  Xinv21 x[20] vss vss vdd vdd x[21] sramgen_svt_inv_2_wrapper
  Xinv22 x[21] vss vss vdd vdd x[22] sramgen_svt_inv_2_wrapper
  Xinv23 x[22] vss vss vdd vdd x[23] sramgen_svt_inv_2_wrapper
  Xinv24 x[23] vss vss vdd vdd x[24] sramgen_svt_inv_2_wrapper
  Xinv25 x[24] vss vss vdd vdd x[25] sramgen_svt_inv_2_wrapper
  Xinv26 x[25] vss vss vdd vdd x[26] sramgen_svt_inv_2_wrapper
  Xinv27 x[26] vss vss vdd vdd x[27] sramgen_svt_inv_2_wrapper
  Xinv28 x[27] vss vss vdd vdd x[28] sramgen_svt_inv_2_wrapper
  Xinv29 x[28] vss vss vdd vdd dout sramgen_svt_inv_4_wrapper

.ENDS svt_inv_chain_30

.SUBCKT inv_chain_14 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sky130_fd_sc_hs__inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd x[2] sky130_fd_sc_hs__inv_2_wrapper
  Xinv3 x[2] vss vss vdd vdd x[3] sky130_fd_sc_hs__inv_2_wrapper
  Xinv4 x[3] vss vss vdd vdd x[4] sky130_fd_sc_hs__inv_2_wrapper
  Xinv5 x[4] vss vss vdd vdd x[5] sky130_fd_sc_hs__inv_2_wrapper
  Xinv6 x[5] vss vss vdd vdd x[6] sky130_fd_sc_hs__inv_2_wrapper
  Xinv7 x[6] vss vss vdd vdd x[7] sky130_fd_sc_hs__inv_2_wrapper
  Xinv8 x[7] vss vss vdd vdd x[8] sky130_fd_sc_hs__inv_2_wrapper
  Xinv9 x[8] vss vss vdd vdd x[9] sky130_fd_sc_hs__inv_2_wrapper
  Xinv10 x[9] vss vss vdd vdd x[10] sky130_fd_sc_hs__inv_2_wrapper
  Xinv11 x[10] vss vss vdd vdd x[11] sky130_fd_sc_hs__inv_2_wrapper
  Xinv12 x[11] vss vss vdd vdd x[12] sky130_fd_sc_hs__inv_2_wrapper
  Xinv13 x[12] vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_14

.SUBCKT sky130_fd_sc_hs__nor2_4 A B VGND VNB VPB VPWR Y

  X0 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 a_27_368# B Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X3 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X4 Y B a_27_368# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X5 a_27_368# B Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X6 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X7 VPWR A a_27_368# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X8 VPWR A a_27_368# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X11 Y B a_27_368# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120


.ENDS sky130_fd_sc_hs__nor2_4

.SUBCKT sky130_fd_sc_hs__nor2_4_wrapper A B VGND VNB VPB VPWR Y

  X0 A B VGND VNB VPB VPWR Y sky130_fd_sc_hs__nor2_4

.ENDS sky130_fd_sc_hs__nor2_4_wrapper

.SUBCKT sky130_fd_sc_hs__nand2_4 A B VGND VNB VPB VPWR Y

  X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X2 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X3 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X4 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X5 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X6 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X8 Y B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X11 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__nand2_4

.SUBCKT sky130_fd_sc_hs__nand2_4_wrapper A B VGND VNB VPB VPWR Y

  X0 A B VGND VNB VPB VPWR Y sky130_fd_sc_hs__nand2_4

.ENDS sky130_fd_sc_hs__nand2_4_wrapper

.SUBCKT inv_chain_2 din dout vdd vss

  Xinv0 din vss vss vdd vdd x sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_2

.SUBCKT control_logic_replica_v2 clk ce we rstb rbl saen pc_b rwl wlen wrdrven vdd vss

  Xreset_inv rstb vss vss vdd vdd reset sky130_fd_sc_hs__inv_16_wrapper
  Xclk_delay clk clkd vdd vss inv_chain_12
  Xclk_gate clkd ce vss vss vdd vdd clk_buf sky130_fd_sc_hs__and2_2_wrapper
  Xclk_pulse clk_buf clkp0 vdd vss edge_detector
  Xclk_pulse_buf clkp0 vss vss vdd vdd clkp sky130_fd_sc_hs__buf_16_wrapper
  Xclk_pulse_inv clkp vss vss vdd vdd clkp_b sky130_fd_sc_hs__inv_16_wrapper
  Xclkp_delay clkp_b clkpd vdd vss inv_chain_3
  Xclkpd_inv clkpd vss vss vdd vdd clkpd_b sky130_fd_sc_hs__inv_2_wrapper
  Xclkpd_delay clkpd_b clkpdd vdd vss inv_chain_15
  Xmux_wlen_rst rbl_b clkpdd we vss vss vdd vdd decrepstart sky130_fd_sc_hs__mux2_4_wrapper
  Xdecoder_replica decrepstart decrepend vdd vss svt_inv_chain_30
  Xdecoder_replica_delay decrepend wlen_rst_decoderd vdd vss inv_chain_14
  Xinv_we we vss vss vdd vdd we_b sky130_fd_sc_hs__inv_2_wrapper
  Xinv_rbl rbl vss vss vdd vdd rbl_b sky130_fd_sc_hs__inv_2_wrapper
  Xwlen_grst decrepstart reset vss vss vdd vdd wlen_grst_b sky130_fd_sc_hs__nor2_4_wrapper
  Xpc_set wlen_rst_decoderd reset vss vss vdd vdd pc_set_b sky130_fd_sc_hs__nor2_4_wrapper
  Xwrdrven_grst decrepend reset vss vss vdd vdd wrdrven_grst_b sky130_fd_sc_hs__nor2_4_wrapper
  Xclkp_grst clkp reset vss vss vdd vdd clkp_grst_b sky130_fd_sc_hs__nor2_4_wrapper
  Xnand_sense_en we_b decrepend vss vss vdd vdd saen_set_b sky130_fd_sc_hs__nand2_4_wrapper
  Xnand_wlendb_web rbl_b we_b vss vss vdd vdd wlend sky130_fd_sc_hs__nand2_4_wrapper
  Xand_wlen wlen_q wlend vss vss vdd vdd wlen sky130_fd_sc_hs__and2_4_wrapper
  Xrwl_buf wlen_q vss vss vdd vdd rwl sky130_fd_sc_hs__buf_16_wrapper
  Xwl_ctl clkpd_b wlen_grst_b wlen_q wlen_b vdd vss sr_latch
  Xsaen_ctl saen_set_b clkp_grst_b saen saen_b vdd vss sr_latch
  Xpc_ctl pc_set_b clkp_b pc pc_b0 vdd vss sr_latch
  Xpc_b_buf pc_b0 vss vss vdd vdd pc_b sky130_fd_sc_hs__buf_16_wrapper
  Xwrdrven_set clkpd we vss vss vdd vdd wrdrven_set_b0 sky130_fd_sc_hs__nand2_4_wrapper
  Xwrdrven_set_delay wrdrven_set_b0 wrdrven_set_b vdd vss inv_chain_2
  Xwrdrven_ctl wrdrven_set_b wrdrven_grst_b wrdrven wrdrven_b vdd vss sr_latch

.ENDS control_logic_replica_v2

.SUBCKT decoder_stage_2 vdd vss y y_b predecode_0_0

  Xgate_0_0_0 vdd vss predecode_0_0 y_b folded_inv
  Xgate_1_0_0 vdd vss y_b y multi_finger_inv_3
  Xgate_1_0_1 vdd vss y_b y multi_finger_inv_3

.ENDS decoder_stage_2

.SUBCKT multi_finger_inv_4 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_4

.SUBCKT decoder_stage_3 vdd vss y y_b predecode_0_0

  Xgate_0_0_0 vdd vss predecode_0_0 y_b folded_inv
  Xgate_1_0_0 vdd vss y_b y multi_finger_inv_4
  Xgate_1_0_1 vdd vss y_b y multi_finger_inv_4

.ENDS decoder_stage_3

.SUBCKT sram_sp_cell BL BR VDD VSS WL VNB VPB

  X0 QB WL BR VNB sky130_fd_pr__special_nfet_pass l=0.150 nf=1 w=0.140

  X1 Q QB VSS VNB sky130_fd_pr__special_nfet_latch l=0.150 nf=1 w=0.210

  X2 BL WL Q VNB sky130_fd_pr__special_nfet_pass l=0.150 nf=1 w=0.140

  X3 Q WL Q VPB sky130_fd_pr__special_pfet_pass l=0.025 nf=1 w=0.140

  X4 QB WL QB VPB sky130_fd_pr__special_pfet_pass l=0.025 nf=1 w=0.140

  X5 VDD Q QB VPB sky130_fd_pr__special_pfet_pass l=0.150 nf=1 w=0.140

  X6 Q QB VDD VPB sky130_fd_pr__special_pfet_pass l=0.150 nf=1 w=0.140

  X7 VSS Q QB VNB sky130_fd_pr__special_nfet_latch l=0.150 nf=1 w=0.210


.ENDS sram_sp_cell

.SUBCKT sram_sp_cell_wrapper BL BR VDD VSS WL VNB VPB

  X0 BL BR VDD VSS WL VNB VPB sram_sp_cell

.ENDS sram_sp_cell_wrapper

.SUBCKT sram_sp_hstrap_wrapper BR VDD VSS BL VNB VPB

  X0 BR VDD VSS BL VNB VPB sram_sp_hstrap

.ENDS sram_sp_hstrap_wrapper

.SUBCKT sram_sp_horiz_wlstrap_p2 VSS VNB

  X0 VSS VSS VSS VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.420


.ENDS sram_sp_horiz_wlstrap_p2

.SUBCKT sram_sp_horiz_wlstrap_p2_wrapper VSS VNB

  X0 VSS VNB sram_sp_horiz_wlstrap_p2

.ENDS sram_sp_horiz_wlstrap_p2_wrapper

.SUBCKT sp_cell_array vdd vss dummy_bl dummy_br bl[0] bl[1] bl[2] bl[3] bl[4] bl[5] bl[6] bl[7] bl[8] bl[9] bl[10] bl[11] bl[12] bl[13] bl[14] bl[15] bl[16] bl[17] bl[18] bl[19] bl[20] bl[21] bl[22] bl[23] bl[24] bl[25] bl[26] bl[27] bl[28] bl[29] bl[30] bl[31] bl[32] bl[33] bl[34] bl[35] bl[36] bl[37] bl[38] bl[39] bl[40] bl[41] bl[42] bl[43] bl[44] bl[45] bl[46] bl[47] bl[48] bl[49] bl[50] bl[51] bl[52] bl[53] bl[54] bl[55] bl[56] bl[57] bl[58] bl[59] bl[60] bl[61] bl[62] bl[63] br[0] br[1] br[2] br[3] br[4] br[5] br[6] br[7] br[8] br[9] br[10] br[11] br[12] br[13] br[14] br[15] br[16] br[17] br[18] br[19] br[20] br[21] br[22] br[23] br[24] br[25] br[26] br[27] br[28] br[29] br[30] br[31] br[32] br[33] br[34] br[35] br[36] br[37] br[38] br[39] br[40] br[41] br[42] br[43] br[44] br[45] br[46] br[47] br[48] br[49] br[50] br[51] br[52] br[53] br[54] br[55] br[56] br[57] br[58] br[59] br[60] br[61] br[62] br[63] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127]

  Xcell_0_0 bl[0] br[0] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_1 bl[1] br[1] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_2 bl[2] br[2] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_3 bl[3] br[3] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_4 bl[4] br[4] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_5 bl[5] br[5] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_6 bl[6] br[6] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_7 bl[7] br[7] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_8 bl[8] br[8] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_9 bl[9] br[9] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_10 bl[10] br[10] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_11 bl[11] br[11] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_12 bl[12] br[12] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_13 bl[13] br[13] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_14 bl[14] br[14] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_15 bl[15] br[15] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_16 bl[16] br[16] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_17 bl[17] br[17] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_18 bl[18] br[18] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_19 bl[19] br[19] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_20 bl[20] br[20] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_21 bl[21] br[21] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_22 bl[22] br[22] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_23 bl[23] br[23] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_24 bl[24] br[24] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_25 bl[25] br[25] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_26 bl[26] br[26] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_27 bl[27] br[27] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_28 bl[28] br[28] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_29 bl[29] br[29] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_30 bl[30] br[30] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_31 bl[31] br[31] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_32 bl[32] br[32] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_33 bl[33] br[33] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_34 bl[34] br[34] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_35 bl[35] br[35] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_36 bl[36] br[36] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_37 bl[37] br[37] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_38 bl[38] br[38] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_39 bl[39] br[39] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_40 bl[40] br[40] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_41 bl[41] br[41] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_42 bl[42] br[42] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_43 bl[43] br[43] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_44 bl[44] br[44] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_45 bl[45] br[45] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_46 bl[46] br[46] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_47 bl[47] br[47] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_48 bl[48] br[48] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_49 bl[49] br[49] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_50 bl[50] br[50] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_51 bl[51] br[51] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_52 bl[52] br[52] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_53 bl[53] br[53] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_54 bl[54] br[54] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_55 bl[55] br[55] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_56 bl[56] br[56] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_57 bl[57] br[57] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_58 bl[58] br[58] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_59 bl[59] br[59] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_60 bl[60] br[60] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_61 bl[61] br[61] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_62 bl[62] br[62] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_63 bl[63] br[63] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_1_0 bl[0] br[0] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_1 bl[1] br[1] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_2 bl[2] br[2] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_3 bl[3] br[3] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_4 bl[4] br[4] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_5 bl[5] br[5] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_6 bl[6] br[6] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_7 bl[7] br[7] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_8 bl[8] br[8] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_9 bl[9] br[9] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_10 bl[10] br[10] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_11 bl[11] br[11] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_12 bl[12] br[12] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_13 bl[13] br[13] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_14 bl[14] br[14] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_15 bl[15] br[15] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_16 bl[16] br[16] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_17 bl[17] br[17] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_18 bl[18] br[18] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_19 bl[19] br[19] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_20 bl[20] br[20] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_21 bl[21] br[21] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_22 bl[22] br[22] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_23 bl[23] br[23] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_24 bl[24] br[24] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_25 bl[25] br[25] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_26 bl[26] br[26] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_27 bl[27] br[27] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_28 bl[28] br[28] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_29 bl[29] br[29] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_30 bl[30] br[30] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_31 bl[31] br[31] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_32 bl[32] br[32] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_33 bl[33] br[33] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_34 bl[34] br[34] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_35 bl[35] br[35] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_36 bl[36] br[36] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_37 bl[37] br[37] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_38 bl[38] br[38] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_39 bl[39] br[39] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_40 bl[40] br[40] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_41 bl[41] br[41] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_42 bl[42] br[42] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_43 bl[43] br[43] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_44 bl[44] br[44] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_45 bl[45] br[45] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_46 bl[46] br[46] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_47 bl[47] br[47] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_48 bl[48] br[48] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_49 bl[49] br[49] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_50 bl[50] br[50] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_51 bl[51] br[51] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_52 bl[52] br[52] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_53 bl[53] br[53] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_54 bl[54] br[54] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_55 bl[55] br[55] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_56 bl[56] br[56] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_57 bl[57] br[57] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_58 bl[58] br[58] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_59 bl[59] br[59] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_60 bl[60] br[60] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_61 bl[61] br[61] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_62 bl[62] br[62] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_63 bl[63] br[63] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_2_0 bl[0] br[0] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_1 bl[1] br[1] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_2 bl[2] br[2] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_3 bl[3] br[3] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_4 bl[4] br[4] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_5 bl[5] br[5] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_6 bl[6] br[6] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_7 bl[7] br[7] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_8 bl[8] br[8] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_9 bl[9] br[9] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_10 bl[10] br[10] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_11 bl[11] br[11] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_12 bl[12] br[12] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_13 bl[13] br[13] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_14 bl[14] br[14] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_15 bl[15] br[15] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_16 bl[16] br[16] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_17 bl[17] br[17] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_18 bl[18] br[18] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_19 bl[19] br[19] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_20 bl[20] br[20] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_21 bl[21] br[21] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_22 bl[22] br[22] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_23 bl[23] br[23] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_24 bl[24] br[24] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_25 bl[25] br[25] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_26 bl[26] br[26] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_27 bl[27] br[27] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_28 bl[28] br[28] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_29 bl[29] br[29] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_30 bl[30] br[30] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_31 bl[31] br[31] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_32 bl[32] br[32] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_33 bl[33] br[33] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_34 bl[34] br[34] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_35 bl[35] br[35] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_36 bl[36] br[36] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_37 bl[37] br[37] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_38 bl[38] br[38] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_39 bl[39] br[39] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_40 bl[40] br[40] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_41 bl[41] br[41] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_42 bl[42] br[42] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_43 bl[43] br[43] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_44 bl[44] br[44] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_45 bl[45] br[45] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_46 bl[46] br[46] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_47 bl[47] br[47] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_48 bl[48] br[48] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_49 bl[49] br[49] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_50 bl[50] br[50] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_51 bl[51] br[51] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_52 bl[52] br[52] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_53 bl[53] br[53] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_54 bl[54] br[54] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_55 bl[55] br[55] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_56 bl[56] br[56] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_57 bl[57] br[57] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_58 bl[58] br[58] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_59 bl[59] br[59] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_60 bl[60] br[60] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_61 bl[61] br[61] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_62 bl[62] br[62] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_63 bl[63] br[63] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_3_0 bl[0] br[0] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_1 bl[1] br[1] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_2 bl[2] br[2] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_3 bl[3] br[3] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_4 bl[4] br[4] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_5 bl[5] br[5] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_6 bl[6] br[6] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_7 bl[7] br[7] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_8 bl[8] br[8] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_9 bl[9] br[9] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_10 bl[10] br[10] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_11 bl[11] br[11] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_12 bl[12] br[12] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_13 bl[13] br[13] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_14 bl[14] br[14] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_15 bl[15] br[15] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_16 bl[16] br[16] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_17 bl[17] br[17] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_18 bl[18] br[18] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_19 bl[19] br[19] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_20 bl[20] br[20] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_21 bl[21] br[21] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_22 bl[22] br[22] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_23 bl[23] br[23] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_24 bl[24] br[24] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_25 bl[25] br[25] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_26 bl[26] br[26] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_27 bl[27] br[27] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_28 bl[28] br[28] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_29 bl[29] br[29] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_30 bl[30] br[30] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_31 bl[31] br[31] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_32 bl[32] br[32] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_33 bl[33] br[33] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_34 bl[34] br[34] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_35 bl[35] br[35] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_36 bl[36] br[36] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_37 bl[37] br[37] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_38 bl[38] br[38] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_39 bl[39] br[39] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_40 bl[40] br[40] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_41 bl[41] br[41] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_42 bl[42] br[42] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_43 bl[43] br[43] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_44 bl[44] br[44] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_45 bl[45] br[45] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_46 bl[46] br[46] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_47 bl[47] br[47] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_48 bl[48] br[48] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_49 bl[49] br[49] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_50 bl[50] br[50] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_51 bl[51] br[51] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_52 bl[52] br[52] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_53 bl[53] br[53] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_54 bl[54] br[54] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_55 bl[55] br[55] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_56 bl[56] br[56] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_57 bl[57] br[57] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_58 bl[58] br[58] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_59 bl[59] br[59] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_60 bl[60] br[60] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_61 bl[61] br[61] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_62 bl[62] br[62] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_63 bl[63] br[63] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_4_0 bl[0] br[0] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_1 bl[1] br[1] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_2 bl[2] br[2] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_3 bl[3] br[3] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_4 bl[4] br[4] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_5 bl[5] br[5] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_6 bl[6] br[6] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_7 bl[7] br[7] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_8 bl[8] br[8] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_9 bl[9] br[9] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_10 bl[10] br[10] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_11 bl[11] br[11] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_12 bl[12] br[12] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_13 bl[13] br[13] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_14 bl[14] br[14] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_15 bl[15] br[15] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_16 bl[16] br[16] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_17 bl[17] br[17] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_18 bl[18] br[18] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_19 bl[19] br[19] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_20 bl[20] br[20] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_21 bl[21] br[21] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_22 bl[22] br[22] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_23 bl[23] br[23] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_24 bl[24] br[24] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_25 bl[25] br[25] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_26 bl[26] br[26] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_27 bl[27] br[27] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_28 bl[28] br[28] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_29 bl[29] br[29] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_30 bl[30] br[30] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_31 bl[31] br[31] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_32 bl[32] br[32] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_33 bl[33] br[33] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_34 bl[34] br[34] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_35 bl[35] br[35] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_36 bl[36] br[36] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_37 bl[37] br[37] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_38 bl[38] br[38] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_39 bl[39] br[39] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_40 bl[40] br[40] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_41 bl[41] br[41] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_42 bl[42] br[42] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_43 bl[43] br[43] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_44 bl[44] br[44] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_45 bl[45] br[45] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_46 bl[46] br[46] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_47 bl[47] br[47] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_48 bl[48] br[48] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_49 bl[49] br[49] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_50 bl[50] br[50] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_51 bl[51] br[51] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_52 bl[52] br[52] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_53 bl[53] br[53] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_54 bl[54] br[54] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_55 bl[55] br[55] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_56 bl[56] br[56] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_57 bl[57] br[57] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_58 bl[58] br[58] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_59 bl[59] br[59] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_60 bl[60] br[60] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_61 bl[61] br[61] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_62 bl[62] br[62] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_63 bl[63] br[63] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_5_0 bl[0] br[0] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_1 bl[1] br[1] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_2 bl[2] br[2] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_3 bl[3] br[3] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_4 bl[4] br[4] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_5 bl[5] br[5] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_6 bl[6] br[6] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_7 bl[7] br[7] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_8 bl[8] br[8] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_9 bl[9] br[9] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_10 bl[10] br[10] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_11 bl[11] br[11] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_12 bl[12] br[12] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_13 bl[13] br[13] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_14 bl[14] br[14] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_15 bl[15] br[15] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_16 bl[16] br[16] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_17 bl[17] br[17] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_18 bl[18] br[18] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_19 bl[19] br[19] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_20 bl[20] br[20] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_21 bl[21] br[21] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_22 bl[22] br[22] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_23 bl[23] br[23] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_24 bl[24] br[24] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_25 bl[25] br[25] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_26 bl[26] br[26] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_27 bl[27] br[27] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_28 bl[28] br[28] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_29 bl[29] br[29] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_30 bl[30] br[30] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_31 bl[31] br[31] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_32 bl[32] br[32] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_33 bl[33] br[33] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_34 bl[34] br[34] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_35 bl[35] br[35] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_36 bl[36] br[36] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_37 bl[37] br[37] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_38 bl[38] br[38] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_39 bl[39] br[39] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_40 bl[40] br[40] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_41 bl[41] br[41] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_42 bl[42] br[42] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_43 bl[43] br[43] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_44 bl[44] br[44] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_45 bl[45] br[45] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_46 bl[46] br[46] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_47 bl[47] br[47] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_48 bl[48] br[48] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_49 bl[49] br[49] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_50 bl[50] br[50] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_51 bl[51] br[51] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_52 bl[52] br[52] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_53 bl[53] br[53] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_54 bl[54] br[54] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_55 bl[55] br[55] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_56 bl[56] br[56] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_57 bl[57] br[57] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_58 bl[58] br[58] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_59 bl[59] br[59] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_60 bl[60] br[60] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_61 bl[61] br[61] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_62 bl[62] br[62] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_63 bl[63] br[63] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_6_0 bl[0] br[0] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_1 bl[1] br[1] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_2 bl[2] br[2] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_3 bl[3] br[3] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_4 bl[4] br[4] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_5 bl[5] br[5] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_6 bl[6] br[6] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_7 bl[7] br[7] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_8 bl[8] br[8] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_9 bl[9] br[9] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_10 bl[10] br[10] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_11 bl[11] br[11] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_12 bl[12] br[12] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_13 bl[13] br[13] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_14 bl[14] br[14] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_15 bl[15] br[15] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_16 bl[16] br[16] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_17 bl[17] br[17] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_18 bl[18] br[18] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_19 bl[19] br[19] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_20 bl[20] br[20] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_21 bl[21] br[21] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_22 bl[22] br[22] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_23 bl[23] br[23] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_24 bl[24] br[24] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_25 bl[25] br[25] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_26 bl[26] br[26] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_27 bl[27] br[27] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_28 bl[28] br[28] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_29 bl[29] br[29] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_30 bl[30] br[30] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_31 bl[31] br[31] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_32 bl[32] br[32] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_33 bl[33] br[33] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_34 bl[34] br[34] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_35 bl[35] br[35] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_36 bl[36] br[36] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_37 bl[37] br[37] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_38 bl[38] br[38] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_39 bl[39] br[39] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_40 bl[40] br[40] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_41 bl[41] br[41] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_42 bl[42] br[42] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_43 bl[43] br[43] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_44 bl[44] br[44] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_45 bl[45] br[45] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_46 bl[46] br[46] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_47 bl[47] br[47] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_48 bl[48] br[48] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_49 bl[49] br[49] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_50 bl[50] br[50] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_51 bl[51] br[51] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_52 bl[52] br[52] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_53 bl[53] br[53] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_54 bl[54] br[54] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_55 bl[55] br[55] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_56 bl[56] br[56] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_57 bl[57] br[57] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_58 bl[58] br[58] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_59 bl[59] br[59] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_60 bl[60] br[60] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_61 bl[61] br[61] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_62 bl[62] br[62] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_63 bl[63] br[63] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_7_0 bl[0] br[0] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_1 bl[1] br[1] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_2 bl[2] br[2] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_3 bl[3] br[3] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_4 bl[4] br[4] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_5 bl[5] br[5] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_6 bl[6] br[6] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_7 bl[7] br[7] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_8 bl[8] br[8] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_9 bl[9] br[9] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_10 bl[10] br[10] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_11 bl[11] br[11] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_12 bl[12] br[12] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_13 bl[13] br[13] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_14 bl[14] br[14] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_15 bl[15] br[15] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_16 bl[16] br[16] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_17 bl[17] br[17] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_18 bl[18] br[18] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_19 bl[19] br[19] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_20 bl[20] br[20] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_21 bl[21] br[21] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_22 bl[22] br[22] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_23 bl[23] br[23] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_24 bl[24] br[24] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_25 bl[25] br[25] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_26 bl[26] br[26] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_27 bl[27] br[27] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_28 bl[28] br[28] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_29 bl[29] br[29] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_30 bl[30] br[30] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_31 bl[31] br[31] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_32 bl[32] br[32] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_33 bl[33] br[33] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_34 bl[34] br[34] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_35 bl[35] br[35] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_36 bl[36] br[36] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_37 bl[37] br[37] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_38 bl[38] br[38] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_39 bl[39] br[39] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_40 bl[40] br[40] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_41 bl[41] br[41] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_42 bl[42] br[42] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_43 bl[43] br[43] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_44 bl[44] br[44] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_45 bl[45] br[45] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_46 bl[46] br[46] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_47 bl[47] br[47] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_48 bl[48] br[48] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_49 bl[49] br[49] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_50 bl[50] br[50] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_51 bl[51] br[51] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_52 bl[52] br[52] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_53 bl[53] br[53] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_54 bl[54] br[54] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_55 bl[55] br[55] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_56 bl[56] br[56] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_57 bl[57] br[57] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_58 bl[58] br[58] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_59 bl[59] br[59] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_60 bl[60] br[60] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_61 bl[61] br[61] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_62 bl[62] br[62] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_63 bl[63] br[63] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_8_0 bl[0] br[0] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_1 bl[1] br[1] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_2 bl[2] br[2] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_3 bl[3] br[3] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_4 bl[4] br[4] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_5 bl[5] br[5] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_6 bl[6] br[6] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_7 bl[7] br[7] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_8 bl[8] br[8] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_9 bl[9] br[9] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_10 bl[10] br[10] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_11 bl[11] br[11] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_12 bl[12] br[12] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_13 bl[13] br[13] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_14 bl[14] br[14] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_15 bl[15] br[15] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_16 bl[16] br[16] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_17 bl[17] br[17] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_18 bl[18] br[18] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_19 bl[19] br[19] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_20 bl[20] br[20] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_21 bl[21] br[21] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_22 bl[22] br[22] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_23 bl[23] br[23] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_24 bl[24] br[24] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_25 bl[25] br[25] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_26 bl[26] br[26] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_27 bl[27] br[27] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_28 bl[28] br[28] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_29 bl[29] br[29] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_30 bl[30] br[30] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_31 bl[31] br[31] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_32 bl[32] br[32] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_33 bl[33] br[33] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_34 bl[34] br[34] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_35 bl[35] br[35] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_36 bl[36] br[36] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_37 bl[37] br[37] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_38 bl[38] br[38] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_39 bl[39] br[39] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_40 bl[40] br[40] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_41 bl[41] br[41] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_42 bl[42] br[42] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_43 bl[43] br[43] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_44 bl[44] br[44] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_45 bl[45] br[45] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_46 bl[46] br[46] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_47 bl[47] br[47] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_48 bl[48] br[48] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_49 bl[49] br[49] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_50 bl[50] br[50] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_51 bl[51] br[51] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_52 bl[52] br[52] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_53 bl[53] br[53] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_54 bl[54] br[54] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_55 bl[55] br[55] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_56 bl[56] br[56] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_57 bl[57] br[57] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_58 bl[58] br[58] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_59 bl[59] br[59] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_60 bl[60] br[60] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_61 bl[61] br[61] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_62 bl[62] br[62] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_63 bl[63] br[63] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_9_0 bl[0] br[0] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_1 bl[1] br[1] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_2 bl[2] br[2] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_3 bl[3] br[3] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_4 bl[4] br[4] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_5 bl[5] br[5] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_6 bl[6] br[6] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_7 bl[7] br[7] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_8 bl[8] br[8] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_9 bl[9] br[9] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_10 bl[10] br[10] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_11 bl[11] br[11] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_12 bl[12] br[12] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_13 bl[13] br[13] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_14 bl[14] br[14] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_15 bl[15] br[15] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_16 bl[16] br[16] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_17 bl[17] br[17] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_18 bl[18] br[18] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_19 bl[19] br[19] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_20 bl[20] br[20] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_21 bl[21] br[21] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_22 bl[22] br[22] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_23 bl[23] br[23] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_24 bl[24] br[24] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_25 bl[25] br[25] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_26 bl[26] br[26] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_27 bl[27] br[27] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_28 bl[28] br[28] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_29 bl[29] br[29] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_30 bl[30] br[30] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_31 bl[31] br[31] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_32 bl[32] br[32] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_33 bl[33] br[33] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_34 bl[34] br[34] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_35 bl[35] br[35] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_36 bl[36] br[36] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_37 bl[37] br[37] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_38 bl[38] br[38] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_39 bl[39] br[39] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_40 bl[40] br[40] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_41 bl[41] br[41] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_42 bl[42] br[42] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_43 bl[43] br[43] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_44 bl[44] br[44] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_45 bl[45] br[45] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_46 bl[46] br[46] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_47 bl[47] br[47] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_48 bl[48] br[48] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_49 bl[49] br[49] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_50 bl[50] br[50] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_51 bl[51] br[51] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_52 bl[52] br[52] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_53 bl[53] br[53] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_54 bl[54] br[54] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_55 bl[55] br[55] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_56 bl[56] br[56] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_57 bl[57] br[57] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_58 bl[58] br[58] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_59 bl[59] br[59] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_60 bl[60] br[60] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_61 bl[61] br[61] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_62 bl[62] br[62] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_63 bl[63] br[63] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_10_0 bl[0] br[0] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_1 bl[1] br[1] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_2 bl[2] br[2] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_3 bl[3] br[3] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_4 bl[4] br[4] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_5 bl[5] br[5] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_6 bl[6] br[6] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_7 bl[7] br[7] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_8 bl[8] br[8] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_9 bl[9] br[9] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_10 bl[10] br[10] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_11 bl[11] br[11] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_12 bl[12] br[12] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_13 bl[13] br[13] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_14 bl[14] br[14] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_15 bl[15] br[15] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_16 bl[16] br[16] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_17 bl[17] br[17] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_18 bl[18] br[18] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_19 bl[19] br[19] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_20 bl[20] br[20] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_21 bl[21] br[21] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_22 bl[22] br[22] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_23 bl[23] br[23] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_24 bl[24] br[24] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_25 bl[25] br[25] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_26 bl[26] br[26] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_27 bl[27] br[27] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_28 bl[28] br[28] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_29 bl[29] br[29] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_30 bl[30] br[30] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_31 bl[31] br[31] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_32 bl[32] br[32] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_33 bl[33] br[33] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_34 bl[34] br[34] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_35 bl[35] br[35] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_36 bl[36] br[36] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_37 bl[37] br[37] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_38 bl[38] br[38] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_39 bl[39] br[39] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_40 bl[40] br[40] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_41 bl[41] br[41] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_42 bl[42] br[42] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_43 bl[43] br[43] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_44 bl[44] br[44] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_45 bl[45] br[45] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_46 bl[46] br[46] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_47 bl[47] br[47] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_48 bl[48] br[48] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_49 bl[49] br[49] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_50 bl[50] br[50] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_51 bl[51] br[51] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_52 bl[52] br[52] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_53 bl[53] br[53] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_54 bl[54] br[54] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_55 bl[55] br[55] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_56 bl[56] br[56] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_57 bl[57] br[57] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_58 bl[58] br[58] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_59 bl[59] br[59] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_60 bl[60] br[60] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_61 bl[61] br[61] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_62 bl[62] br[62] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_63 bl[63] br[63] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_11_0 bl[0] br[0] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_1 bl[1] br[1] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_2 bl[2] br[2] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_3 bl[3] br[3] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_4 bl[4] br[4] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_5 bl[5] br[5] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_6 bl[6] br[6] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_7 bl[7] br[7] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_8 bl[8] br[8] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_9 bl[9] br[9] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_10 bl[10] br[10] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_11 bl[11] br[11] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_12 bl[12] br[12] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_13 bl[13] br[13] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_14 bl[14] br[14] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_15 bl[15] br[15] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_16 bl[16] br[16] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_17 bl[17] br[17] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_18 bl[18] br[18] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_19 bl[19] br[19] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_20 bl[20] br[20] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_21 bl[21] br[21] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_22 bl[22] br[22] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_23 bl[23] br[23] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_24 bl[24] br[24] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_25 bl[25] br[25] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_26 bl[26] br[26] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_27 bl[27] br[27] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_28 bl[28] br[28] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_29 bl[29] br[29] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_30 bl[30] br[30] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_31 bl[31] br[31] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_32 bl[32] br[32] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_33 bl[33] br[33] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_34 bl[34] br[34] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_35 bl[35] br[35] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_36 bl[36] br[36] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_37 bl[37] br[37] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_38 bl[38] br[38] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_39 bl[39] br[39] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_40 bl[40] br[40] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_41 bl[41] br[41] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_42 bl[42] br[42] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_43 bl[43] br[43] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_44 bl[44] br[44] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_45 bl[45] br[45] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_46 bl[46] br[46] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_47 bl[47] br[47] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_48 bl[48] br[48] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_49 bl[49] br[49] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_50 bl[50] br[50] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_51 bl[51] br[51] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_52 bl[52] br[52] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_53 bl[53] br[53] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_54 bl[54] br[54] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_55 bl[55] br[55] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_56 bl[56] br[56] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_57 bl[57] br[57] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_58 bl[58] br[58] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_59 bl[59] br[59] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_60 bl[60] br[60] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_61 bl[61] br[61] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_62 bl[62] br[62] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_63 bl[63] br[63] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_12_0 bl[0] br[0] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_1 bl[1] br[1] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_2 bl[2] br[2] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_3 bl[3] br[3] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_4 bl[4] br[4] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_5 bl[5] br[5] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_6 bl[6] br[6] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_7 bl[7] br[7] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_8 bl[8] br[8] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_9 bl[9] br[9] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_10 bl[10] br[10] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_11 bl[11] br[11] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_12 bl[12] br[12] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_13 bl[13] br[13] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_14 bl[14] br[14] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_15 bl[15] br[15] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_16 bl[16] br[16] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_17 bl[17] br[17] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_18 bl[18] br[18] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_19 bl[19] br[19] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_20 bl[20] br[20] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_21 bl[21] br[21] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_22 bl[22] br[22] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_23 bl[23] br[23] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_24 bl[24] br[24] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_25 bl[25] br[25] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_26 bl[26] br[26] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_27 bl[27] br[27] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_28 bl[28] br[28] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_29 bl[29] br[29] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_30 bl[30] br[30] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_31 bl[31] br[31] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_32 bl[32] br[32] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_33 bl[33] br[33] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_34 bl[34] br[34] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_35 bl[35] br[35] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_36 bl[36] br[36] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_37 bl[37] br[37] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_38 bl[38] br[38] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_39 bl[39] br[39] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_40 bl[40] br[40] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_41 bl[41] br[41] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_42 bl[42] br[42] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_43 bl[43] br[43] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_44 bl[44] br[44] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_45 bl[45] br[45] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_46 bl[46] br[46] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_47 bl[47] br[47] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_48 bl[48] br[48] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_49 bl[49] br[49] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_50 bl[50] br[50] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_51 bl[51] br[51] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_52 bl[52] br[52] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_53 bl[53] br[53] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_54 bl[54] br[54] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_55 bl[55] br[55] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_56 bl[56] br[56] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_57 bl[57] br[57] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_58 bl[58] br[58] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_59 bl[59] br[59] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_60 bl[60] br[60] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_61 bl[61] br[61] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_62 bl[62] br[62] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_63 bl[63] br[63] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_13_0 bl[0] br[0] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_1 bl[1] br[1] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_2 bl[2] br[2] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_3 bl[3] br[3] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_4 bl[4] br[4] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_5 bl[5] br[5] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_6 bl[6] br[6] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_7 bl[7] br[7] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_8 bl[8] br[8] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_9 bl[9] br[9] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_10 bl[10] br[10] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_11 bl[11] br[11] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_12 bl[12] br[12] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_13 bl[13] br[13] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_14 bl[14] br[14] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_15 bl[15] br[15] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_16 bl[16] br[16] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_17 bl[17] br[17] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_18 bl[18] br[18] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_19 bl[19] br[19] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_20 bl[20] br[20] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_21 bl[21] br[21] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_22 bl[22] br[22] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_23 bl[23] br[23] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_24 bl[24] br[24] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_25 bl[25] br[25] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_26 bl[26] br[26] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_27 bl[27] br[27] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_28 bl[28] br[28] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_29 bl[29] br[29] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_30 bl[30] br[30] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_31 bl[31] br[31] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_32 bl[32] br[32] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_33 bl[33] br[33] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_34 bl[34] br[34] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_35 bl[35] br[35] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_36 bl[36] br[36] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_37 bl[37] br[37] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_38 bl[38] br[38] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_39 bl[39] br[39] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_40 bl[40] br[40] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_41 bl[41] br[41] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_42 bl[42] br[42] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_43 bl[43] br[43] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_44 bl[44] br[44] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_45 bl[45] br[45] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_46 bl[46] br[46] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_47 bl[47] br[47] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_48 bl[48] br[48] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_49 bl[49] br[49] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_50 bl[50] br[50] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_51 bl[51] br[51] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_52 bl[52] br[52] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_53 bl[53] br[53] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_54 bl[54] br[54] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_55 bl[55] br[55] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_56 bl[56] br[56] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_57 bl[57] br[57] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_58 bl[58] br[58] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_59 bl[59] br[59] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_60 bl[60] br[60] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_61 bl[61] br[61] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_62 bl[62] br[62] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_63 bl[63] br[63] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_14_0 bl[0] br[0] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_1 bl[1] br[1] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_2 bl[2] br[2] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_3 bl[3] br[3] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_4 bl[4] br[4] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_5 bl[5] br[5] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_6 bl[6] br[6] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_7 bl[7] br[7] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_8 bl[8] br[8] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_9 bl[9] br[9] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_10 bl[10] br[10] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_11 bl[11] br[11] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_12 bl[12] br[12] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_13 bl[13] br[13] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_14 bl[14] br[14] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_15 bl[15] br[15] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_16 bl[16] br[16] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_17 bl[17] br[17] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_18 bl[18] br[18] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_19 bl[19] br[19] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_20 bl[20] br[20] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_21 bl[21] br[21] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_22 bl[22] br[22] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_23 bl[23] br[23] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_24 bl[24] br[24] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_25 bl[25] br[25] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_26 bl[26] br[26] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_27 bl[27] br[27] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_28 bl[28] br[28] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_29 bl[29] br[29] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_30 bl[30] br[30] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_31 bl[31] br[31] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_32 bl[32] br[32] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_33 bl[33] br[33] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_34 bl[34] br[34] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_35 bl[35] br[35] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_36 bl[36] br[36] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_37 bl[37] br[37] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_38 bl[38] br[38] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_39 bl[39] br[39] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_40 bl[40] br[40] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_41 bl[41] br[41] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_42 bl[42] br[42] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_43 bl[43] br[43] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_44 bl[44] br[44] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_45 bl[45] br[45] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_46 bl[46] br[46] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_47 bl[47] br[47] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_48 bl[48] br[48] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_49 bl[49] br[49] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_50 bl[50] br[50] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_51 bl[51] br[51] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_52 bl[52] br[52] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_53 bl[53] br[53] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_54 bl[54] br[54] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_55 bl[55] br[55] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_56 bl[56] br[56] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_57 bl[57] br[57] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_58 bl[58] br[58] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_59 bl[59] br[59] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_60 bl[60] br[60] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_61 bl[61] br[61] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_62 bl[62] br[62] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_63 bl[63] br[63] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_15_0 bl[0] br[0] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_1 bl[1] br[1] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_2 bl[2] br[2] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_3 bl[3] br[3] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_4 bl[4] br[4] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_5 bl[5] br[5] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_6 bl[6] br[6] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_7 bl[7] br[7] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_8 bl[8] br[8] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_9 bl[9] br[9] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_10 bl[10] br[10] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_11 bl[11] br[11] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_12 bl[12] br[12] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_13 bl[13] br[13] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_14 bl[14] br[14] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_15 bl[15] br[15] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_16 bl[16] br[16] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_17 bl[17] br[17] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_18 bl[18] br[18] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_19 bl[19] br[19] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_20 bl[20] br[20] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_21 bl[21] br[21] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_22 bl[22] br[22] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_23 bl[23] br[23] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_24 bl[24] br[24] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_25 bl[25] br[25] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_26 bl[26] br[26] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_27 bl[27] br[27] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_28 bl[28] br[28] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_29 bl[29] br[29] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_30 bl[30] br[30] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_31 bl[31] br[31] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_32 bl[32] br[32] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_33 bl[33] br[33] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_34 bl[34] br[34] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_35 bl[35] br[35] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_36 bl[36] br[36] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_37 bl[37] br[37] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_38 bl[38] br[38] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_39 bl[39] br[39] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_40 bl[40] br[40] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_41 bl[41] br[41] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_42 bl[42] br[42] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_43 bl[43] br[43] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_44 bl[44] br[44] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_45 bl[45] br[45] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_46 bl[46] br[46] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_47 bl[47] br[47] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_48 bl[48] br[48] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_49 bl[49] br[49] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_50 bl[50] br[50] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_51 bl[51] br[51] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_52 bl[52] br[52] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_53 bl[53] br[53] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_54 bl[54] br[54] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_55 bl[55] br[55] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_56 bl[56] br[56] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_57 bl[57] br[57] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_58 bl[58] br[58] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_59 bl[59] br[59] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_60 bl[60] br[60] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_61 bl[61] br[61] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_62 bl[62] br[62] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_63 bl[63] br[63] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_16_0 bl[0] br[0] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_1 bl[1] br[1] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_2 bl[2] br[2] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_3 bl[3] br[3] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_4 bl[4] br[4] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_5 bl[5] br[5] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_6 bl[6] br[6] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_7 bl[7] br[7] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_8 bl[8] br[8] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_9 bl[9] br[9] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_10 bl[10] br[10] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_11 bl[11] br[11] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_12 bl[12] br[12] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_13 bl[13] br[13] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_14 bl[14] br[14] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_15 bl[15] br[15] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_16 bl[16] br[16] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_17 bl[17] br[17] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_18 bl[18] br[18] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_19 bl[19] br[19] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_20 bl[20] br[20] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_21 bl[21] br[21] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_22 bl[22] br[22] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_23 bl[23] br[23] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_24 bl[24] br[24] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_25 bl[25] br[25] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_26 bl[26] br[26] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_27 bl[27] br[27] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_28 bl[28] br[28] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_29 bl[29] br[29] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_30 bl[30] br[30] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_31 bl[31] br[31] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_32 bl[32] br[32] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_33 bl[33] br[33] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_34 bl[34] br[34] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_35 bl[35] br[35] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_36 bl[36] br[36] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_37 bl[37] br[37] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_38 bl[38] br[38] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_39 bl[39] br[39] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_40 bl[40] br[40] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_41 bl[41] br[41] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_42 bl[42] br[42] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_43 bl[43] br[43] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_44 bl[44] br[44] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_45 bl[45] br[45] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_46 bl[46] br[46] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_47 bl[47] br[47] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_48 bl[48] br[48] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_49 bl[49] br[49] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_50 bl[50] br[50] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_51 bl[51] br[51] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_52 bl[52] br[52] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_53 bl[53] br[53] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_54 bl[54] br[54] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_55 bl[55] br[55] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_56 bl[56] br[56] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_57 bl[57] br[57] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_58 bl[58] br[58] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_59 bl[59] br[59] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_60 bl[60] br[60] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_61 bl[61] br[61] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_62 bl[62] br[62] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_63 bl[63] br[63] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_17_0 bl[0] br[0] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_1 bl[1] br[1] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_2 bl[2] br[2] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_3 bl[3] br[3] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_4 bl[4] br[4] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_5 bl[5] br[5] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_6 bl[6] br[6] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_7 bl[7] br[7] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_8 bl[8] br[8] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_9 bl[9] br[9] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_10 bl[10] br[10] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_11 bl[11] br[11] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_12 bl[12] br[12] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_13 bl[13] br[13] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_14 bl[14] br[14] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_15 bl[15] br[15] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_16 bl[16] br[16] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_17 bl[17] br[17] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_18 bl[18] br[18] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_19 bl[19] br[19] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_20 bl[20] br[20] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_21 bl[21] br[21] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_22 bl[22] br[22] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_23 bl[23] br[23] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_24 bl[24] br[24] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_25 bl[25] br[25] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_26 bl[26] br[26] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_27 bl[27] br[27] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_28 bl[28] br[28] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_29 bl[29] br[29] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_30 bl[30] br[30] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_31 bl[31] br[31] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_32 bl[32] br[32] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_33 bl[33] br[33] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_34 bl[34] br[34] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_35 bl[35] br[35] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_36 bl[36] br[36] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_37 bl[37] br[37] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_38 bl[38] br[38] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_39 bl[39] br[39] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_40 bl[40] br[40] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_41 bl[41] br[41] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_42 bl[42] br[42] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_43 bl[43] br[43] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_44 bl[44] br[44] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_45 bl[45] br[45] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_46 bl[46] br[46] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_47 bl[47] br[47] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_48 bl[48] br[48] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_49 bl[49] br[49] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_50 bl[50] br[50] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_51 bl[51] br[51] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_52 bl[52] br[52] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_53 bl[53] br[53] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_54 bl[54] br[54] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_55 bl[55] br[55] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_56 bl[56] br[56] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_57 bl[57] br[57] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_58 bl[58] br[58] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_59 bl[59] br[59] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_60 bl[60] br[60] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_61 bl[61] br[61] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_62 bl[62] br[62] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_63 bl[63] br[63] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_18_0 bl[0] br[0] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_1 bl[1] br[1] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_2 bl[2] br[2] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_3 bl[3] br[3] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_4 bl[4] br[4] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_5 bl[5] br[5] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_6 bl[6] br[6] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_7 bl[7] br[7] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_8 bl[8] br[8] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_9 bl[9] br[9] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_10 bl[10] br[10] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_11 bl[11] br[11] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_12 bl[12] br[12] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_13 bl[13] br[13] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_14 bl[14] br[14] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_15 bl[15] br[15] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_16 bl[16] br[16] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_17 bl[17] br[17] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_18 bl[18] br[18] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_19 bl[19] br[19] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_20 bl[20] br[20] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_21 bl[21] br[21] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_22 bl[22] br[22] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_23 bl[23] br[23] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_24 bl[24] br[24] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_25 bl[25] br[25] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_26 bl[26] br[26] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_27 bl[27] br[27] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_28 bl[28] br[28] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_29 bl[29] br[29] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_30 bl[30] br[30] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_31 bl[31] br[31] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_32 bl[32] br[32] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_33 bl[33] br[33] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_34 bl[34] br[34] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_35 bl[35] br[35] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_36 bl[36] br[36] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_37 bl[37] br[37] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_38 bl[38] br[38] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_39 bl[39] br[39] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_40 bl[40] br[40] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_41 bl[41] br[41] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_42 bl[42] br[42] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_43 bl[43] br[43] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_44 bl[44] br[44] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_45 bl[45] br[45] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_46 bl[46] br[46] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_47 bl[47] br[47] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_48 bl[48] br[48] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_49 bl[49] br[49] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_50 bl[50] br[50] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_51 bl[51] br[51] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_52 bl[52] br[52] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_53 bl[53] br[53] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_54 bl[54] br[54] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_55 bl[55] br[55] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_56 bl[56] br[56] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_57 bl[57] br[57] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_58 bl[58] br[58] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_59 bl[59] br[59] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_60 bl[60] br[60] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_61 bl[61] br[61] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_62 bl[62] br[62] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_63 bl[63] br[63] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_19_0 bl[0] br[0] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_1 bl[1] br[1] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_2 bl[2] br[2] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_3 bl[3] br[3] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_4 bl[4] br[4] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_5 bl[5] br[5] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_6 bl[6] br[6] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_7 bl[7] br[7] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_8 bl[8] br[8] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_9 bl[9] br[9] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_10 bl[10] br[10] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_11 bl[11] br[11] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_12 bl[12] br[12] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_13 bl[13] br[13] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_14 bl[14] br[14] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_15 bl[15] br[15] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_16 bl[16] br[16] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_17 bl[17] br[17] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_18 bl[18] br[18] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_19 bl[19] br[19] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_20 bl[20] br[20] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_21 bl[21] br[21] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_22 bl[22] br[22] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_23 bl[23] br[23] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_24 bl[24] br[24] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_25 bl[25] br[25] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_26 bl[26] br[26] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_27 bl[27] br[27] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_28 bl[28] br[28] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_29 bl[29] br[29] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_30 bl[30] br[30] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_31 bl[31] br[31] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_32 bl[32] br[32] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_33 bl[33] br[33] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_34 bl[34] br[34] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_35 bl[35] br[35] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_36 bl[36] br[36] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_37 bl[37] br[37] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_38 bl[38] br[38] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_39 bl[39] br[39] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_40 bl[40] br[40] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_41 bl[41] br[41] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_42 bl[42] br[42] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_43 bl[43] br[43] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_44 bl[44] br[44] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_45 bl[45] br[45] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_46 bl[46] br[46] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_47 bl[47] br[47] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_48 bl[48] br[48] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_49 bl[49] br[49] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_50 bl[50] br[50] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_51 bl[51] br[51] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_52 bl[52] br[52] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_53 bl[53] br[53] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_54 bl[54] br[54] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_55 bl[55] br[55] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_56 bl[56] br[56] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_57 bl[57] br[57] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_58 bl[58] br[58] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_59 bl[59] br[59] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_60 bl[60] br[60] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_61 bl[61] br[61] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_62 bl[62] br[62] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_63 bl[63] br[63] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_20_0 bl[0] br[0] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_1 bl[1] br[1] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_2 bl[2] br[2] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_3 bl[3] br[3] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_4 bl[4] br[4] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_5 bl[5] br[5] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_6 bl[6] br[6] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_7 bl[7] br[7] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_8 bl[8] br[8] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_9 bl[9] br[9] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_10 bl[10] br[10] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_11 bl[11] br[11] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_12 bl[12] br[12] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_13 bl[13] br[13] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_14 bl[14] br[14] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_15 bl[15] br[15] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_16 bl[16] br[16] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_17 bl[17] br[17] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_18 bl[18] br[18] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_19 bl[19] br[19] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_20 bl[20] br[20] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_21 bl[21] br[21] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_22 bl[22] br[22] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_23 bl[23] br[23] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_24 bl[24] br[24] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_25 bl[25] br[25] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_26 bl[26] br[26] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_27 bl[27] br[27] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_28 bl[28] br[28] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_29 bl[29] br[29] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_30 bl[30] br[30] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_31 bl[31] br[31] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_32 bl[32] br[32] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_33 bl[33] br[33] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_34 bl[34] br[34] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_35 bl[35] br[35] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_36 bl[36] br[36] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_37 bl[37] br[37] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_38 bl[38] br[38] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_39 bl[39] br[39] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_40 bl[40] br[40] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_41 bl[41] br[41] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_42 bl[42] br[42] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_43 bl[43] br[43] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_44 bl[44] br[44] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_45 bl[45] br[45] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_46 bl[46] br[46] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_47 bl[47] br[47] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_48 bl[48] br[48] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_49 bl[49] br[49] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_50 bl[50] br[50] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_51 bl[51] br[51] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_52 bl[52] br[52] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_53 bl[53] br[53] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_54 bl[54] br[54] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_55 bl[55] br[55] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_56 bl[56] br[56] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_57 bl[57] br[57] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_58 bl[58] br[58] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_59 bl[59] br[59] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_60 bl[60] br[60] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_61 bl[61] br[61] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_62 bl[62] br[62] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_63 bl[63] br[63] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_21_0 bl[0] br[0] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_1 bl[1] br[1] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_2 bl[2] br[2] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_3 bl[3] br[3] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_4 bl[4] br[4] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_5 bl[5] br[5] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_6 bl[6] br[6] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_7 bl[7] br[7] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_8 bl[8] br[8] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_9 bl[9] br[9] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_10 bl[10] br[10] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_11 bl[11] br[11] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_12 bl[12] br[12] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_13 bl[13] br[13] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_14 bl[14] br[14] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_15 bl[15] br[15] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_16 bl[16] br[16] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_17 bl[17] br[17] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_18 bl[18] br[18] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_19 bl[19] br[19] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_20 bl[20] br[20] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_21 bl[21] br[21] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_22 bl[22] br[22] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_23 bl[23] br[23] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_24 bl[24] br[24] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_25 bl[25] br[25] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_26 bl[26] br[26] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_27 bl[27] br[27] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_28 bl[28] br[28] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_29 bl[29] br[29] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_30 bl[30] br[30] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_31 bl[31] br[31] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_32 bl[32] br[32] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_33 bl[33] br[33] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_34 bl[34] br[34] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_35 bl[35] br[35] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_36 bl[36] br[36] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_37 bl[37] br[37] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_38 bl[38] br[38] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_39 bl[39] br[39] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_40 bl[40] br[40] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_41 bl[41] br[41] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_42 bl[42] br[42] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_43 bl[43] br[43] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_44 bl[44] br[44] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_45 bl[45] br[45] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_46 bl[46] br[46] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_47 bl[47] br[47] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_48 bl[48] br[48] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_49 bl[49] br[49] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_50 bl[50] br[50] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_51 bl[51] br[51] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_52 bl[52] br[52] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_53 bl[53] br[53] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_54 bl[54] br[54] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_55 bl[55] br[55] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_56 bl[56] br[56] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_57 bl[57] br[57] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_58 bl[58] br[58] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_59 bl[59] br[59] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_60 bl[60] br[60] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_61 bl[61] br[61] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_62 bl[62] br[62] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_63 bl[63] br[63] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_22_0 bl[0] br[0] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_1 bl[1] br[1] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_2 bl[2] br[2] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_3 bl[3] br[3] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_4 bl[4] br[4] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_5 bl[5] br[5] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_6 bl[6] br[6] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_7 bl[7] br[7] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_8 bl[8] br[8] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_9 bl[9] br[9] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_10 bl[10] br[10] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_11 bl[11] br[11] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_12 bl[12] br[12] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_13 bl[13] br[13] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_14 bl[14] br[14] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_15 bl[15] br[15] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_16 bl[16] br[16] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_17 bl[17] br[17] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_18 bl[18] br[18] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_19 bl[19] br[19] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_20 bl[20] br[20] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_21 bl[21] br[21] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_22 bl[22] br[22] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_23 bl[23] br[23] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_24 bl[24] br[24] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_25 bl[25] br[25] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_26 bl[26] br[26] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_27 bl[27] br[27] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_28 bl[28] br[28] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_29 bl[29] br[29] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_30 bl[30] br[30] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_31 bl[31] br[31] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_32 bl[32] br[32] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_33 bl[33] br[33] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_34 bl[34] br[34] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_35 bl[35] br[35] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_36 bl[36] br[36] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_37 bl[37] br[37] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_38 bl[38] br[38] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_39 bl[39] br[39] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_40 bl[40] br[40] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_41 bl[41] br[41] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_42 bl[42] br[42] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_43 bl[43] br[43] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_44 bl[44] br[44] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_45 bl[45] br[45] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_46 bl[46] br[46] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_47 bl[47] br[47] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_48 bl[48] br[48] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_49 bl[49] br[49] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_50 bl[50] br[50] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_51 bl[51] br[51] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_52 bl[52] br[52] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_53 bl[53] br[53] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_54 bl[54] br[54] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_55 bl[55] br[55] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_56 bl[56] br[56] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_57 bl[57] br[57] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_58 bl[58] br[58] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_59 bl[59] br[59] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_60 bl[60] br[60] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_61 bl[61] br[61] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_62 bl[62] br[62] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_63 bl[63] br[63] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_23_0 bl[0] br[0] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_1 bl[1] br[1] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_2 bl[2] br[2] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_3 bl[3] br[3] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_4 bl[4] br[4] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_5 bl[5] br[5] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_6 bl[6] br[6] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_7 bl[7] br[7] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_8 bl[8] br[8] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_9 bl[9] br[9] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_10 bl[10] br[10] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_11 bl[11] br[11] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_12 bl[12] br[12] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_13 bl[13] br[13] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_14 bl[14] br[14] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_15 bl[15] br[15] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_16 bl[16] br[16] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_17 bl[17] br[17] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_18 bl[18] br[18] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_19 bl[19] br[19] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_20 bl[20] br[20] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_21 bl[21] br[21] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_22 bl[22] br[22] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_23 bl[23] br[23] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_24 bl[24] br[24] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_25 bl[25] br[25] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_26 bl[26] br[26] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_27 bl[27] br[27] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_28 bl[28] br[28] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_29 bl[29] br[29] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_30 bl[30] br[30] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_31 bl[31] br[31] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_32 bl[32] br[32] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_33 bl[33] br[33] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_34 bl[34] br[34] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_35 bl[35] br[35] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_36 bl[36] br[36] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_37 bl[37] br[37] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_38 bl[38] br[38] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_39 bl[39] br[39] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_40 bl[40] br[40] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_41 bl[41] br[41] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_42 bl[42] br[42] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_43 bl[43] br[43] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_44 bl[44] br[44] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_45 bl[45] br[45] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_46 bl[46] br[46] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_47 bl[47] br[47] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_48 bl[48] br[48] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_49 bl[49] br[49] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_50 bl[50] br[50] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_51 bl[51] br[51] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_52 bl[52] br[52] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_53 bl[53] br[53] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_54 bl[54] br[54] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_55 bl[55] br[55] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_56 bl[56] br[56] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_57 bl[57] br[57] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_58 bl[58] br[58] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_59 bl[59] br[59] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_60 bl[60] br[60] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_61 bl[61] br[61] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_62 bl[62] br[62] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_63 bl[63] br[63] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_24_0 bl[0] br[0] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_1 bl[1] br[1] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_2 bl[2] br[2] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_3 bl[3] br[3] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_4 bl[4] br[4] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_5 bl[5] br[5] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_6 bl[6] br[6] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_7 bl[7] br[7] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_8 bl[8] br[8] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_9 bl[9] br[9] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_10 bl[10] br[10] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_11 bl[11] br[11] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_12 bl[12] br[12] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_13 bl[13] br[13] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_14 bl[14] br[14] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_15 bl[15] br[15] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_16 bl[16] br[16] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_17 bl[17] br[17] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_18 bl[18] br[18] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_19 bl[19] br[19] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_20 bl[20] br[20] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_21 bl[21] br[21] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_22 bl[22] br[22] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_23 bl[23] br[23] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_24 bl[24] br[24] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_25 bl[25] br[25] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_26 bl[26] br[26] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_27 bl[27] br[27] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_28 bl[28] br[28] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_29 bl[29] br[29] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_30 bl[30] br[30] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_31 bl[31] br[31] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_32 bl[32] br[32] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_33 bl[33] br[33] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_34 bl[34] br[34] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_35 bl[35] br[35] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_36 bl[36] br[36] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_37 bl[37] br[37] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_38 bl[38] br[38] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_39 bl[39] br[39] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_40 bl[40] br[40] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_41 bl[41] br[41] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_42 bl[42] br[42] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_43 bl[43] br[43] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_44 bl[44] br[44] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_45 bl[45] br[45] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_46 bl[46] br[46] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_47 bl[47] br[47] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_48 bl[48] br[48] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_49 bl[49] br[49] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_50 bl[50] br[50] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_51 bl[51] br[51] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_52 bl[52] br[52] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_53 bl[53] br[53] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_54 bl[54] br[54] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_55 bl[55] br[55] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_56 bl[56] br[56] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_57 bl[57] br[57] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_58 bl[58] br[58] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_59 bl[59] br[59] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_60 bl[60] br[60] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_61 bl[61] br[61] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_62 bl[62] br[62] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_63 bl[63] br[63] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_25_0 bl[0] br[0] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_1 bl[1] br[1] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_2 bl[2] br[2] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_3 bl[3] br[3] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_4 bl[4] br[4] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_5 bl[5] br[5] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_6 bl[6] br[6] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_7 bl[7] br[7] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_8 bl[8] br[8] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_9 bl[9] br[9] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_10 bl[10] br[10] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_11 bl[11] br[11] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_12 bl[12] br[12] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_13 bl[13] br[13] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_14 bl[14] br[14] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_15 bl[15] br[15] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_16 bl[16] br[16] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_17 bl[17] br[17] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_18 bl[18] br[18] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_19 bl[19] br[19] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_20 bl[20] br[20] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_21 bl[21] br[21] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_22 bl[22] br[22] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_23 bl[23] br[23] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_24 bl[24] br[24] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_25 bl[25] br[25] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_26 bl[26] br[26] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_27 bl[27] br[27] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_28 bl[28] br[28] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_29 bl[29] br[29] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_30 bl[30] br[30] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_31 bl[31] br[31] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_32 bl[32] br[32] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_33 bl[33] br[33] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_34 bl[34] br[34] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_35 bl[35] br[35] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_36 bl[36] br[36] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_37 bl[37] br[37] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_38 bl[38] br[38] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_39 bl[39] br[39] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_40 bl[40] br[40] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_41 bl[41] br[41] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_42 bl[42] br[42] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_43 bl[43] br[43] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_44 bl[44] br[44] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_45 bl[45] br[45] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_46 bl[46] br[46] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_47 bl[47] br[47] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_48 bl[48] br[48] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_49 bl[49] br[49] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_50 bl[50] br[50] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_51 bl[51] br[51] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_52 bl[52] br[52] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_53 bl[53] br[53] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_54 bl[54] br[54] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_55 bl[55] br[55] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_56 bl[56] br[56] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_57 bl[57] br[57] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_58 bl[58] br[58] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_59 bl[59] br[59] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_60 bl[60] br[60] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_61 bl[61] br[61] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_62 bl[62] br[62] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_63 bl[63] br[63] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_26_0 bl[0] br[0] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_1 bl[1] br[1] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_2 bl[2] br[2] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_3 bl[3] br[3] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_4 bl[4] br[4] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_5 bl[5] br[5] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_6 bl[6] br[6] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_7 bl[7] br[7] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_8 bl[8] br[8] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_9 bl[9] br[9] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_10 bl[10] br[10] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_11 bl[11] br[11] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_12 bl[12] br[12] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_13 bl[13] br[13] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_14 bl[14] br[14] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_15 bl[15] br[15] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_16 bl[16] br[16] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_17 bl[17] br[17] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_18 bl[18] br[18] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_19 bl[19] br[19] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_20 bl[20] br[20] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_21 bl[21] br[21] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_22 bl[22] br[22] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_23 bl[23] br[23] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_24 bl[24] br[24] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_25 bl[25] br[25] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_26 bl[26] br[26] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_27 bl[27] br[27] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_28 bl[28] br[28] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_29 bl[29] br[29] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_30 bl[30] br[30] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_31 bl[31] br[31] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_32 bl[32] br[32] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_33 bl[33] br[33] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_34 bl[34] br[34] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_35 bl[35] br[35] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_36 bl[36] br[36] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_37 bl[37] br[37] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_38 bl[38] br[38] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_39 bl[39] br[39] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_40 bl[40] br[40] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_41 bl[41] br[41] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_42 bl[42] br[42] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_43 bl[43] br[43] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_44 bl[44] br[44] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_45 bl[45] br[45] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_46 bl[46] br[46] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_47 bl[47] br[47] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_48 bl[48] br[48] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_49 bl[49] br[49] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_50 bl[50] br[50] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_51 bl[51] br[51] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_52 bl[52] br[52] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_53 bl[53] br[53] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_54 bl[54] br[54] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_55 bl[55] br[55] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_56 bl[56] br[56] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_57 bl[57] br[57] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_58 bl[58] br[58] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_59 bl[59] br[59] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_60 bl[60] br[60] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_61 bl[61] br[61] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_62 bl[62] br[62] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_63 bl[63] br[63] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_27_0 bl[0] br[0] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_1 bl[1] br[1] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_2 bl[2] br[2] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_3 bl[3] br[3] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_4 bl[4] br[4] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_5 bl[5] br[5] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_6 bl[6] br[6] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_7 bl[7] br[7] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_8 bl[8] br[8] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_9 bl[9] br[9] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_10 bl[10] br[10] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_11 bl[11] br[11] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_12 bl[12] br[12] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_13 bl[13] br[13] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_14 bl[14] br[14] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_15 bl[15] br[15] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_16 bl[16] br[16] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_17 bl[17] br[17] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_18 bl[18] br[18] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_19 bl[19] br[19] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_20 bl[20] br[20] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_21 bl[21] br[21] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_22 bl[22] br[22] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_23 bl[23] br[23] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_24 bl[24] br[24] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_25 bl[25] br[25] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_26 bl[26] br[26] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_27 bl[27] br[27] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_28 bl[28] br[28] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_29 bl[29] br[29] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_30 bl[30] br[30] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_31 bl[31] br[31] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_32 bl[32] br[32] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_33 bl[33] br[33] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_34 bl[34] br[34] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_35 bl[35] br[35] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_36 bl[36] br[36] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_37 bl[37] br[37] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_38 bl[38] br[38] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_39 bl[39] br[39] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_40 bl[40] br[40] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_41 bl[41] br[41] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_42 bl[42] br[42] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_43 bl[43] br[43] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_44 bl[44] br[44] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_45 bl[45] br[45] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_46 bl[46] br[46] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_47 bl[47] br[47] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_48 bl[48] br[48] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_49 bl[49] br[49] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_50 bl[50] br[50] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_51 bl[51] br[51] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_52 bl[52] br[52] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_53 bl[53] br[53] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_54 bl[54] br[54] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_55 bl[55] br[55] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_56 bl[56] br[56] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_57 bl[57] br[57] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_58 bl[58] br[58] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_59 bl[59] br[59] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_60 bl[60] br[60] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_61 bl[61] br[61] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_62 bl[62] br[62] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_63 bl[63] br[63] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_28_0 bl[0] br[0] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_1 bl[1] br[1] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_2 bl[2] br[2] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_3 bl[3] br[3] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_4 bl[4] br[4] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_5 bl[5] br[5] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_6 bl[6] br[6] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_7 bl[7] br[7] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_8 bl[8] br[8] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_9 bl[9] br[9] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_10 bl[10] br[10] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_11 bl[11] br[11] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_12 bl[12] br[12] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_13 bl[13] br[13] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_14 bl[14] br[14] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_15 bl[15] br[15] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_16 bl[16] br[16] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_17 bl[17] br[17] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_18 bl[18] br[18] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_19 bl[19] br[19] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_20 bl[20] br[20] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_21 bl[21] br[21] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_22 bl[22] br[22] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_23 bl[23] br[23] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_24 bl[24] br[24] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_25 bl[25] br[25] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_26 bl[26] br[26] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_27 bl[27] br[27] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_28 bl[28] br[28] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_29 bl[29] br[29] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_30 bl[30] br[30] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_31 bl[31] br[31] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_32 bl[32] br[32] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_33 bl[33] br[33] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_34 bl[34] br[34] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_35 bl[35] br[35] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_36 bl[36] br[36] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_37 bl[37] br[37] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_38 bl[38] br[38] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_39 bl[39] br[39] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_40 bl[40] br[40] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_41 bl[41] br[41] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_42 bl[42] br[42] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_43 bl[43] br[43] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_44 bl[44] br[44] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_45 bl[45] br[45] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_46 bl[46] br[46] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_47 bl[47] br[47] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_48 bl[48] br[48] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_49 bl[49] br[49] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_50 bl[50] br[50] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_51 bl[51] br[51] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_52 bl[52] br[52] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_53 bl[53] br[53] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_54 bl[54] br[54] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_55 bl[55] br[55] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_56 bl[56] br[56] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_57 bl[57] br[57] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_58 bl[58] br[58] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_59 bl[59] br[59] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_60 bl[60] br[60] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_61 bl[61] br[61] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_62 bl[62] br[62] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_63 bl[63] br[63] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_29_0 bl[0] br[0] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_1 bl[1] br[1] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_2 bl[2] br[2] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_3 bl[3] br[3] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_4 bl[4] br[4] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_5 bl[5] br[5] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_6 bl[6] br[6] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_7 bl[7] br[7] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_8 bl[8] br[8] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_9 bl[9] br[9] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_10 bl[10] br[10] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_11 bl[11] br[11] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_12 bl[12] br[12] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_13 bl[13] br[13] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_14 bl[14] br[14] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_15 bl[15] br[15] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_16 bl[16] br[16] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_17 bl[17] br[17] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_18 bl[18] br[18] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_19 bl[19] br[19] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_20 bl[20] br[20] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_21 bl[21] br[21] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_22 bl[22] br[22] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_23 bl[23] br[23] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_24 bl[24] br[24] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_25 bl[25] br[25] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_26 bl[26] br[26] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_27 bl[27] br[27] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_28 bl[28] br[28] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_29 bl[29] br[29] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_30 bl[30] br[30] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_31 bl[31] br[31] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_32 bl[32] br[32] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_33 bl[33] br[33] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_34 bl[34] br[34] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_35 bl[35] br[35] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_36 bl[36] br[36] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_37 bl[37] br[37] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_38 bl[38] br[38] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_39 bl[39] br[39] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_40 bl[40] br[40] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_41 bl[41] br[41] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_42 bl[42] br[42] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_43 bl[43] br[43] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_44 bl[44] br[44] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_45 bl[45] br[45] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_46 bl[46] br[46] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_47 bl[47] br[47] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_48 bl[48] br[48] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_49 bl[49] br[49] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_50 bl[50] br[50] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_51 bl[51] br[51] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_52 bl[52] br[52] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_53 bl[53] br[53] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_54 bl[54] br[54] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_55 bl[55] br[55] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_56 bl[56] br[56] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_57 bl[57] br[57] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_58 bl[58] br[58] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_59 bl[59] br[59] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_60 bl[60] br[60] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_61 bl[61] br[61] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_62 bl[62] br[62] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_63 bl[63] br[63] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_30_0 bl[0] br[0] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_1 bl[1] br[1] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_2 bl[2] br[2] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_3 bl[3] br[3] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_4 bl[4] br[4] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_5 bl[5] br[5] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_6 bl[6] br[6] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_7 bl[7] br[7] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_8 bl[8] br[8] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_9 bl[9] br[9] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_10 bl[10] br[10] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_11 bl[11] br[11] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_12 bl[12] br[12] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_13 bl[13] br[13] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_14 bl[14] br[14] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_15 bl[15] br[15] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_16 bl[16] br[16] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_17 bl[17] br[17] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_18 bl[18] br[18] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_19 bl[19] br[19] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_20 bl[20] br[20] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_21 bl[21] br[21] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_22 bl[22] br[22] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_23 bl[23] br[23] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_24 bl[24] br[24] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_25 bl[25] br[25] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_26 bl[26] br[26] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_27 bl[27] br[27] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_28 bl[28] br[28] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_29 bl[29] br[29] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_30 bl[30] br[30] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_31 bl[31] br[31] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_32 bl[32] br[32] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_33 bl[33] br[33] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_34 bl[34] br[34] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_35 bl[35] br[35] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_36 bl[36] br[36] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_37 bl[37] br[37] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_38 bl[38] br[38] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_39 bl[39] br[39] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_40 bl[40] br[40] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_41 bl[41] br[41] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_42 bl[42] br[42] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_43 bl[43] br[43] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_44 bl[44] br[44] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_45 bl[45] br[45] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_46 bl[46] br[46] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_47 bl[47] br[47] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_48 bl[48] br[48] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_49 bl[49] br[49] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_50 bl[50] br[50] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_51 bl[51] br[51] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_52 bl[52] br[52] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_53 bl[53] br[53] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_54 bl[54] br[54] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_55 bl[55] br[55] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_56 bl[56] br[56] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_57 bl[57] br[57] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_58 bl[58] br[58] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_59 bl[59] br[59] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_60 bl[60] br[60] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_61 bl[61] br[61] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_62 bl[62] br[62] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_63 bl[63] br[63] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_31_0 bl[0] br[0] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_1 bl[1] br[1] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_2 bl[2] br[2] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_3 bl[3] br[3] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_4 bl[4] br[4] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_5 bl[5] br[5] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_6 bl[6] br[6] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_7 bl[7] br[7] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_8 bl[8] br[8] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_9 bl[9] br[9] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_10 bl[10] br[10] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_11 bl[11] br[11] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_12 bl[12] br[12] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_13 bl[13] br[13] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_14 bl[14] br[14] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_15 bl[15] br[15] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_16 bl[16] br[16] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_17 bl[17] br[17] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_18 bl[18] br[18] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_19 bl[19] br[19] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_20 bl[20] br[20] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_21 bl[21] br[21] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_22 bl[22] br[22] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_23 bl[23] br[23] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_24 bl[24] br[24] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_25 bl[25] br[25] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_26 bl[26] br[26] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_27 bl[27] br[27] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_28 bl[28] br[28] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_29 bl[29] br[29] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_30 bl[30] br[30] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_31 bl[31] br[31] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_32 bl[32] br[32] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_33 bl[33] br[33] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_34 bl[34] br[34] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_35 bl[35] br[35] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_36 bl[36] br[36] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_37 bl[37] br[37] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_38 bl[38] br[38] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_39 bl[39] br[39] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_40 bl[40] br[40] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_41 bl[41] br[41] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_42 bl[42] br[42] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_43 bl[43] br[43] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_44 bl[44] br[44] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_45 bl[45] br[45] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_46 bl[46] br[46] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_47 bl[47] br[47] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_48 bl[48] br[48] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_49 bl[49] br[49] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_50 bl[50] br[50] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_51 bl[51] br[51] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_52 bl[52] br[52] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_53 bl[53] br[53] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_54 bl[54] br[54] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_55 bl[55] br[55] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_56 bl[56] br[56] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_57 bl[57] br[57] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_58 bl[58] br[58] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_59 bl[59] br[59] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_60 bl[60] br[60] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_61 bl[61] br[61] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_62 bl[62] br[62] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_63 bl[63] br[63] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_32_0 bl[0] br[0] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_1 bl[1] br[1] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_2 bl[2] br[2] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_3 bl[3] br[3] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_4 bl[4] br[4] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_5 bl[5] br[5] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_6 bl[6] br[6] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_7 bl[7] br[7] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_8 bl[8] br[8] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_9 bl[9] br[9] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_10 bl[10] br[10] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_11 bl[11] br[11] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_12 bl[12] br[12] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_13 bl[13] br[13] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_14 bl[14] br[14] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_15 bl[15] br[15] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_16 bl[16] br[16] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_17 bl[17] br[17] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_18 bl[18] br[18] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_19 bl[19] br[19] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_20 bl[20] br[20] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_21 bl[21] br[21] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_22 bl[22] br[22] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_23 bl[23] br[23] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_24 bl[24] br[24] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_25 bl[25] br[25] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_26 bl[26] br[26] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_27 bl[27] br[27] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_28 bl[28] br[28] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_29 bl[29] br[29] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_30 bl[30] br[30] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_31 bl[31] br[31] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_32 bl[32] br[32] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_33 bl[33] br[33] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_34 bl[34] br[34] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_35 bl[35] br[35] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_36 bl[36] br[36] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_37 bl[37] br[37] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_38 bl[38] br[38] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_39 bl[39] br[39] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_40 bl[40] br[40] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_41 bl[41] br[41] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_42 bl[42] br[42] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_43 bl[43] br[43] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_44 bl[44] br[44] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_45 bl[45] br[45] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_46 bl[46] br[46] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_47 bl[47] br[47] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_48 bl[48] br[48] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_49 bl[49] br[49] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_50 bl[50] br[50] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_51 bl[51] br[51] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_52 bl[52] br[52] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_53 bl[53] br[53] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_54 bl[54] br[54] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_55 bl[55] br[55] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_56 bl[56] br[56] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_57 bl[57] br[57] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_58 bl[58] br[58] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_59 bl[59] br[59] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_60 bl[60] br[60] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_61 bl[61] br[61] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_62 bl[62] br[62] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_63 bl[63] br[63] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_33_0 bl[0] br[0] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_1 bl[1] br[1] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_2 bl[2] br[2] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_3 bl[3] br[3] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_4 bl[4] br[4] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_5 bl[5] br[5] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_6 bl[6] br[6] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_7 bl[7] br[7] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_8 bl[8] br[8] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_9 bl[9] br[9] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_10 bl[10] br[10] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_11 bl[11] br[11] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_12 bl[12] br[12] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_13 bl[13] br[13] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_14 bl[14] br[14] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_15 bl[15] br[15] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_16 bl[16] br[16] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_17 bl[17] br[17] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_18 bl[18] br[18] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_19 bl[19] br[19] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_20 bl[20] br[20] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_21 bl[21] br[21] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_22 bl[22] br[22] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_23 bl[23] br[23] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_24 bl[24] br[24] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_25 bl[25] br[25] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_26 bl[26] br[26] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_27 bl[27] br[27] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_28 bl[28] br[28] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_29 bl[29] br[29] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_30 bl[30] br[30] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_31 bl[31] br[31] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_32 bl[32] br[32] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_33 bl[33] br[33] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_34 bl[34] br[34] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_35 bl[35] br[35] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_36 bl[36] br[36] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_37 bl[37] br[37] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_38 bl[38] br[38] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_39 bl[39] br[39] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_40 bl[40] br[40] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_41 bl[41] br[41] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_42 bl[42] br[42] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_43 bl[43] br[43] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_44 bl[44] br[44] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_45 bl[45] br[45] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_46 bl[46] br[46] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_47 bl[47] br[47] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_48 bl[48] br[48] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_49 bl[49] br[49] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_50 bl[50] br[50] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_51 bl[51] br[51] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_52 bl[52] br[52] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_53 bl[53] br[53] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_54 bl[54] br[54] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_55 bl[55] br[55] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_56 bl[56] br[56] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_57 bl[57] br[57] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_58 bl[58] br[58] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_59 bl[59] br[59] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_60 bl[60] br[60] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_61 bl[61] br[61] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_62 bl[62] br[62] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_63 bl[63] br[63] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_34_0 bl[0] br[0] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_1 bl[1] br[1] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_2 bl[2] br[2] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_3 bl[3] br[3] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_4 bl[4] br[4] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_5 bl[5] br[5] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_6 bl[6] br[6] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_7 bl[7] br[7] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_8 bl[8] br[8] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_9 bl[9] br[9] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_10 bl[10] br[10] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_11 bl[11] br[11] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_12 bl[12] br[12] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_13 bl[13] br[13] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_14 bl[14] br[14] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_15 bl[15] br[15] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_16 bl[16] br[16] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_17 bl[17] br[17] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_18 bl[18] br[18] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_19 bl[19] br[19] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_20 bl[20] br[20] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_21 bl[21] br[21] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_22 bl[22] br[22] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_23 bl[23] br[23] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_24 bl[24] br[24] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_25 bl[25] br[25] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_26 bl[26] br[26] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_27 bl[27] br[27] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_28 bl[28] br[28] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_29 bl[29] br[29] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_30 bl[30] br[30] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_31 bl[31] br[31] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_32 bl[32] br[32] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_33 bl[33] br[33] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_34 bl[34] br[34] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_35 bl[35] br[35] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_36 bl[36] br[36] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_37 bl[37] br[37] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_38 bl[38] br[38] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_39 bl[39] br[39] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_40 bl[40] br[40] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_41 bl[41] br[41] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_42 bl[42] br[42] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_43 bl[43] br[43] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_44 bl[44] br[44] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_45 bl[45] br[45] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_46 bl[46] br[46] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_47 bl[47] br[47] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_48 bl[48] br[48] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_49 bl[49] br[49] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_50 bl[50] br[50] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_51 bl[51] br[51] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_52 bl[52] br[52] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_53 bl[53] br[53] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_54 bl[54] br[54] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_55 bl[55] br[55] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_56 bl[56] br[56] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_57 bl[57] br[57] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_58 bl[58] br[58] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_59 bl[59] br[59] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_60 bl[60] br[60] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_61 bl[61] br[61] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_62 bl[62] br[62] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_63 bl[63] br[63] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_35_0 bl[0] br[0] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_1 bl[1] br[1] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_2 bl[2] br[2] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_3 bl[3] br[3] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_4 bl[4] br[4] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_5 bl[5] br[5] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_6 bl[6] br[6] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_7 bl[7] br[7] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_8 bl[8] br[8] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_9 bl[9] br[9] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_10 bl[10] br[10] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_11 bl[11] br[11] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_12 bl[12] br[12] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_13 bl[13] br[13] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_14 bl[14] br[14] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_15 bl[15] br[15] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_16 bl[16] br[16] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_17 bl[17] br[17] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_18 bl[18] br[18] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_19 bl[19] br[19] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_20 bl[20] br[20] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_21 bl[21] br[21] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_22 bl[22] br[22] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_23 bl[23] br[23] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_24 bl[24] br[24] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_25 bl[25] br[25] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_26 bl[26] br[26] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_27 bl[27] br[27] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_28 bl[28] br[28] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_29 bl[29] br[29] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_30 bl[30] br[30] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_31 bl[31] br[31] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_32 bl[32] br[32] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_33 bl[33] br[33] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_34 bl[34] br[34] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_35 bl[35] br[35] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_36 bl[36] br[36] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_37 bl[37] br[37] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_38 bl[38] br[38] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_39 bl[39] br[39] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_40 bl[40] br[40] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_41 bl[41] br[41] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_42 bl[42] br[42] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_43 bl[43] br[43] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_44 bl[44] br[44] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_45 bl[45] br[45] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_46 bl[46] br[46] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_47 bl[47] br[47] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_48 bl[48] br[48] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_49 bl[49] br[49] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_50 bl[50] br[50] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_51 bl[51] br[51] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_52 bl[52] br[52] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_53 bl[53] br[53] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_54 bl[54] br[54] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_55 bl[55] br[55] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_56 bl[56] br[56] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_57 bl[57] br[57] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_58 bl[58] br[58] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_59 bl[59] br[59] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_60 bl[60] br[60] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_61 bl[61] br[61] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_62 bl[62] br[62] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_63 bl[63] br[63] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_36_0 bl[0] br[0] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_1 bl[1] br[1] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_2 bl[2] br[2] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_3 bl[3] br[3] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_4 bl[4] br[4] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_5 bl[5] br[5] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_6 bl[6] br[6] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_7 bl[7] br[7] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_8 bl[8] br[8] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_9 bl[9] br[9] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_10 bl[10] br[10] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_11 bl[11] br[11] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_12 bl[12] br[12] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_13 bl[13] br[13] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_14 bl[14] br[14] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_15 bl[15] br[15] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_16 bl[16] br[16] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_17 bl[17] br[17] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_18 bl[18] br[18] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_19 bl[19] br[19] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_20 bl[20] br[20] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_21 bl[21] br[21] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_22 bl[22] br[22] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_23 bl[23] br[23] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_24 bl[24] br[24] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_25 bl[25] br[25] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_26 bl[26] br[26] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_27 bl[27] br[27] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_28 bl[28] br[28] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_29 bl[29] br[29] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_30 bl[30] br[30] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_31 bl[31] br[31] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_32 bl[32] br[32] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_33 bl[33] br[33] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_34 bl[34] br[34] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_35 bl[35] br[35] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_36 bl[36] br[36] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_37 bl[37] br[37] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_38 bl[38] br[38] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_39 bl[39] br[39] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_40 bl[40] br[40] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_41 bl[41] br[41] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_42 bl[42] br[42] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_43 bl[43] br[43] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_44 bl[44] br[44] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_45 bl[45] br[45] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_46 bl[46] br[46] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_47 bl[47] br[47] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_48 bl[48] br[48] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_49 bl[49] br[49] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_50 bl[50] br[50] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_51 bl[51] br[51] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_52 bl[52] br[52] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_53 bl[53] br[53] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_54 bl[54] br[54] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_55 bl[55] br[55] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_56 bl[56] br[56] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_57 bl[57] br[57] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_58 bl[58] br[58] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_59 bl[59] br[59] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_60 bl[60] br[60] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_61 bl[61] br[61] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_62 bl[62] br[62] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_63 bl[63] br[63] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_37_0 bl[0] br[0] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_1 bl[1] br[1] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_2 bl[2] br[2] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_3 bl[3] br[3] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_4 bl[4] br[4] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_5 bl[5] br[5] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_6 bl[6] br[6] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_7 bl[7] br[7] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_8 bl[8] br[8] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_9 bl[9] br[9] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_10 bl[10] br[10] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_11 bl[11] br[11] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_12 bl[12] br[12] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_13 bl[13] br[13] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_14 bl[14] br[14] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_15 bl[15] br[15] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_16 bl[16] br[16] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_17 bl[17] br[17] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_18 bl[18] br[18] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_19 bl[19] br[19] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_20 bl[20] br[20] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_21 bl[21] br[21] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_22 bl[22] br[22] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_23 bl[23] br[23] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_24 bl[24] br[24] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_25 bl[25] br[25] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_26 bl[26] br[26] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_27 bl[27] br[27] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_28 bl[28] br[28] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_29 bl[29] br[29] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_30 bl[30] br[30] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_31 bl[31] br[31] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_32 bl[32] br[32] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_33 bl[33] br[33] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_34 bl[34] br[34] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_35 bl[35] br[35] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_36 bl[36] br[36] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_37 bl[37] br[37] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_38 bl[38] br[38] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_39 bl[39] br[39] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_40 bl[40] br[40] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_41 bl[41] br[41] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_42 bl[42] br[42] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_43 bl[43] br[43] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_44 bl[44] br[44] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_45 bl[45] br[45] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_46 bl[46] br[46] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_47 bl[47] br[47] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_48 bl[48] br[48] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_49 bl[49] br[49] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_50 bl[50] br[50] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_51 bl[51] br[51] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_52 bl[52] br[52] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_53 bl[53] br[53] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_54 bl[54] br[54] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_55 bl[55] br[55] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_56 bl[56] br[56] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_57 bl[57] br[57] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_58 bl[58] br[58] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_59 bl[59] br[59] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_60 bl[60] br[60] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_61 bl[61] br[61] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_62 bl[62] br[62] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_63 bl[63] br[63] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_38_0 bl[0] br[0] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_1 bl[1] br[1] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_2 bl[2] br[2] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_3 bl[3] br[3] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_4 bl[4] br[4] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_5 bl[5] br[5] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_6 bl[6] br[6] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_7 bl[7] br[7] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_8 bl[8] br[8] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_9 bl[9] br[9] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_10 bl[10] br[10] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_11 bl[11] br[11] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_12 bl[12] br[12] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_13 bl[13] br[13] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_14 bl[14] br[14] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_15 bl[15] br[15] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_16 bl[16] br[16] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_17 bl[17] br[17] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_18 bl[18] br[18] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_19 bl[19] br[19] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_20 bl[20] br[20] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_21 bl[21] br[21] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_22 bl[22] br[22] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_23 bl[23] br[23] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_24 bl[24] br[24] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_25 bl[25] br[25] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_26 bl[26] br[26] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_27 bl[27] br[27] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_28 bl[28] br[28] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_29 bl[29] br[29] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_30 bl[30] br[30] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_31 bl[31] br[31] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_32 bl[32] br[32] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_33 bl[33] br[33] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_34 bl[34] br[34] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_35 bl[35] br[35] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_36 bl[36] br[36] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_37 bl[37] br[37] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_38 bl[38] br[38] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_39 bl[39] br[39] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_40 bl[40] br[40] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_41 bl[41] br[41] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_42 bl[42] br[42] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_43 bl[43] br[43] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_44 bl[44] br[44] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_45 bl[45] br[45] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_46 bl[46] br[46] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_47 bl[47] br[47] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_48 bl[48] br[48] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_49 bl[49] br[49] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_50 bl[50] br[50] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_51 bl[51] br[51] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_52 bl[52] br[52] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_53 bl[53] br[53] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_54 bl[54] br[54] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_55 bl[55] br[55] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_56 bl[56] br[56] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_57 bl[57] br[57] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_58 bl[58] br[58] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_59 bl[59] br[59] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_60 bl[60] br[60] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_61 bl[61] br[61] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_62 bl[62] br[62] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_63 bl[63] br[63] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_39_0 bl[0] br[0] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_1 bl[1] br[1] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_2 bl[2] br[2] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_3 bl[3] br[3] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_4 bl[4] br[4] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_5 bl[5] br[5] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_6 bl[6] br[6] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_7 bl[7] br[7] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_8 bl[8] br[8] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_9 bl[9] br[9] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_10 bl[10] br[10] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_11 bl[11] br[11] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_12 bl[12] br[12] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_13 bl[13] br[13] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_14 bl[14] br[14] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_15 bl[15] br[15] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_16 bl[16] br[16] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_17 bl[17] br[17] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_18 bl[18] br[18] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_19 bl[19] br[19] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_20 bl[20] br[20] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_21 bl[21] br[21] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_22 bl[22] br[22] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_23 bl[23] br[23] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_24 bl[24] br[24] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_25 bl[25] br[25] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_26 bl[26] br[26] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_27 bl[27] br[27] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_28 bl[28] br[28] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_29 bl[29] br[29] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_30 bl[30] br[30] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_31 bl[31] br[31] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_32 bl[32] br[32] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_33 bl[33] br[33] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_34 bl[34] br[34] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_35 bl[35] br[35] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_36 bl[36] br[36] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_37 bl[37] br[37] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_38 bl[38] br[38] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_39 bl[39] br[39] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_40 bl[40] br[40] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_41 bl[41] br[41] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_42 bl[42] br[42] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_43 bl[43] br[43] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_44 bl[44] br[44] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_45 bl[45] br[45] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_46 bl[46] br[46] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_47 bl[47] br[47] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_48 bl[48] br[48] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_49 bl[49] br[49] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_50 bl[50] br[50] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_51 bl[51] br[51] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_52 bl[52] br[52] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_53 bl[53] br[53] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_54 bl[54] br[54] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_55 bl[55] br[55] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_56 bl[56] br[56] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_57 bl[57] br[57] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_58 bl[58] br[58] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_59 bl[59] br[59] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_60 bl[60] br[60] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_61 bl[61] br[61] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_62 bl[62] br[62] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_63 bl[63] br[63] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_40_0 bl[0] br[0] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_1 bl[1] br[1] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_2 bl[2] br[2] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_3 bl[3] br[3] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_4 bl[4] br[4] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_5 bl[5] br[5] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_6 bl[6] br[6] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_7 bl[7] br[7] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_8 bl[8] br[8] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_9 bl[9] br[9] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_10 bl[10] br[10] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_11 bl[11] br[11] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_12 bl[12] br[12] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_13 bl[13] br[13] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_14 bl[14] br[14] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_15 bl[15] br[15] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_16 bl[16] br[16] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_17 bl[17] br[17] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_18 bl[18] br[18] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_19 bl[19] br[19] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_20 bl[20] br[20] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_21 bl[21] br[21] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_22 bl[22] br[22] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_23 bl[23] br[23] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_24 bl[24] br[24] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_25 bl[25] br[25] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_26 bl[26] br[26] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_27 bl[27] br[27] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_28 bl[28] br[28] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_29 bl[29] br[29] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_30 bl[30] br[30] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_31 bl[31] br[31] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_32 bl[32] br[32] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_33 bl[33] br[33] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_34 bl[34] br[34] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_35 bl[35] br[35] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_36 bl[36] br[36] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_37 bl[37] br[37] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_38 bl[38] br[38] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_39 bl[39] br[39] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_40 bl[40] br[40] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_41 bl[41] br[41] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_42 bl[42] br[42] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_43 bl[43] br[43] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_44 bl[44] br[44] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_45 bl[45] br[45] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_46 bl[46] br[46] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_47 bl[47] br[47] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_48 bl[48] br[48] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_49 bl[49] br[49] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_50 bl[50] br[50] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_51 bl[51] br[51] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_52 bl[52] br[52] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_53 bl[53] br[53] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_54 bl[54] br[54] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_55 bl[55] br[55] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_56 bl[56] br[56] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_57 bl[57] br[57] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_58 bl[58] br[58] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_59 bl[59] br[59] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_60 bl[60] br[60] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_61 bl[61] br[61] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_62 bl[62] br[62] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_63 bl[63] br[63] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_41_0 bl[0] br[0] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_1 bl[1] br[1] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_2 bl[2] br[2] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_3 bl[3] br[3] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_4 bl[4] br[4] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_5 bl[5] br[5] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_6 bl[6] br[6] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_7 bl[7] br[7] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_8 bl[8] br[8] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_9 bl[9] br[9] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_10 bl[10] br[10] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_11 bl[11] br[11] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_12 bl[12] br[12] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_13 bl[13] br[13] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_14 bl[14] br[14] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_15 bl[15] br[15] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_16 bl[16] br[16] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_17 bl[17] br[17] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_18 bl[18] br[18] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_19 bl[19] br[19] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_20 bl[20] br[20] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_21 bl[21] br[21] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_22 bl[22] br[22] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_23 bl[23] br[23] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_24 bl[24] br[24] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_25 bl[25] br[25] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_26 bl[26] br[26] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_27 bl[27] br[27] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_28 bl[28] br[28] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_29 bl[29] br[29] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_30 bl[30] br[30] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_31 bl[31] br[31] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_32 bl[32] br[32] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_33 bl[33] br[33] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_34 bl[34] br[34] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_35 bl[35] br[35] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_36 bl[36] br[36] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_37 bl[37] br[37] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_38 bl[38] br[38] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_39 bl[39] br[39] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_40 bl[40] br[40] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_41 bl[41] br[41] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_42 bl[42] br[42] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_43 bl[43] br[43] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_44 bl[44] br[44] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_45 bl[45] br[45] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_46 bl[46] br[46] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_47 bl[47] br[47] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_48 bl[48] br[48] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_49 bl[49] br[49] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_50 bl[50] br[50] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_51 bl[51] br[51] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_52 bl[52] br[52] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_53 bl[53] br[53] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_54 bl[54] br[54] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_55 bl[55] br[55] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_56 bl[56] br[56] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_57 bl[57] br[57] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_58 bl[58] br[58] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_59 bl[59] br[59] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_60 bl[60] br[60] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_61 bl[61] br[61] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_62 bl[62] br[62] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_63 bl[63] br[63] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_42_0 bl[0] br[0] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_1 bl[1] br[1] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_2 bl[2] br[2] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_3 bl[3] br[3] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_4 bl[4] br[4] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_5 bl[5] br[5] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_6 bl[6] br[6] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_7 bl[7] br[7] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_8 bl[8] br[8] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_9 bl[9] br[9] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_10 bl[10] br[10] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_11 bl[11] br[11] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_12 bl[12] br[12] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_13 bl[13] br[13] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_14 bl[14] br[14] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_15 bl[15] br[15] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_16 bl[16] br[16] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_17 bl[17] br[17] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_18 bl[18] br[18] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_19 bl[19] br[19] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_20 bl[20] br[20] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_21 bl[21] br[21] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_22 bl[22] br[22] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_23 bl[23] br[23] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_24 bl[24] br[24] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_25 bl[25] br[25] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_26 bl[26] br[26] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_27 bl[27] br[27] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_28 bl[28] br[28] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_29 bl[29] br[29] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_30 bl[30] br[30] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_31 bl[31] br[31] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_32 bl[32] br[32] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_33 bl[33] br[33] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_34 bl[34] br[34] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_35 bl[35] br[35] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_36 bl[36] br[36] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_37 bl[37] br[37] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_38 bl[38] br[38] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_39 bl[39] br[39] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_40 bl[40] br[40] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_41 bl[41] br[41] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_42 bl[42] br[42] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_43 bl[43] br[43] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_44 bl[44] br[44] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_45 bl[45] br[45] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_46 bl[46] br[46] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_47 bl[47] br[47] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_48 bl[48] br[48] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_49 bl[49] br[49] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_50 bl[50] br[50] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_51 bl[51] br[51] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_52 bl[52] br[52] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_53 bl[53] br[53] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_54 bl[54] br[54] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_55 bl[55] br[55] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_56 bl[56] br[56] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_57 bl[57] br[57] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_58 bl[58] br[58] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_59 bl[59] br[59] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_60 bl[60] br[60] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_61 bl[61] br[61] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_62 bl[62] br[62] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_63 bl[63] br[63] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_43_0 bl[0] br[0] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_1 bl[1] br[1] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_2 bl[2] br[2] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_3 bl[3] br[3] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_4 bl[4] br[4] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_5 bl[5] br[5] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_6 bl[6] br[6] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_7 bl[7] br[7] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_8 bl[8] br[8] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_9 bl[9] br[9] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_10 bl[10] br[10] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_11 bl[11] br[11] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_12 bl[12] br[12] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_13 bl[13] br[13] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_14 bl[14] br[14] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_15 bl[15] br[15] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_16 bl[16] br[16] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_17 bl[17] br[17] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_18 bl[18] br[18] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_19 bl[19] br[19] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_20 bl[20] br[20] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_21 bl[21] br[21] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_22 bl[22] br[22] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_23 bl[23] br[23] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_24 bl[24] br[24] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_25 bl[25] br[25] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_26 bl[26] br[26] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_27 bl[27] br[27] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_28 bl[28] br[28] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_29 bl[29] br[29] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_30 bl[30] br[30] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_31 bl[31] br[31] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_32 bl[32] br[32] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_33 bl[33] br[33] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_34 bl[34] br[34] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_35 bl[35] br[35] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_36 bl[36] br[36] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_37 bl[37] br[37] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_38 bl[38] br[38] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_39 bl[39] br[39] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_40 bl[40] br[40] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_41 bl[41] br[41] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_42 bl[42] br[42] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_43 bl[43] br[43] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_44 bl[44] br[44] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_45 bl[45] br[45] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_46 bl[46] br[46] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_47 bl[47] br[47] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_48 bl[48] br[48] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_49 bl[49] br[49] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_50 bl[50] br[50] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_51 bl[51] br[51] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_52 bl[52] br[52] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_53 bl[53] br[53] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_54 bl[54] br[54] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_55 bl[55] br[55] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_56 bl[56] br[56] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_57 bl[57] br[57] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_58 bl[58] br[58] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_59 bl[59] br[59] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_60 bl[60] br[60] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_61 bl[61] br[61] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_62 bl[62] br[62] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_63 bl[63] br[63] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_44_0 bl[0] br[0] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_1 bl[1] br[1] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_2 bl[2] br[2] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_3 bl[3] br[3] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_4 bl[4] br[4] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_5 bl[5] br[5] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_6 bl[6] br[6] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_7 bl[7] br[7] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_8 bl[8] br[8] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_9 bl[9] br[9] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_10 bl[10] br[10] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_11 bl[11] br[11] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_12 bl[12] br[12] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_13 bl[13] br[13] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_14 bl[14] br[14] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_15 bl[15] br[15] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_16 bl[16] br[16] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_17 bl[17] br[17] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_18 bl[18] br[18] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_19 bl[19] br[19] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_20 bl[20] br[20] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_21 bl[21] br[21] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_22 bl[22] br[22] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_23 bl[23] br[23] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_24 bl[24] br[24] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_25 bl[25] br[25] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_26 bl[26] br[26] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_27 bl[27] br[27] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_28 bl[28] br[28] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_29 bl[29] br[29] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_30 bl[30] br[30] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_31 bl[31] br[31] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_32 bl[32] br[32] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_33 bl[33] br[33] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_34 bl[34] br[34] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_35 bl[35] br[35] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_36 bl[36] br[36] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_37 bl[37] br[37] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_38 bl[38] br[38] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_39 bl[39] br[39] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_40 bl[40] br[40] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_41 bl[41] br[41] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_42 bl[42] br[42] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_43 bl[43] br[43] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_44 bl[44] br[44] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_45 bl[45] br[45] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_46 bl[46] br[46] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_47 bl[47] br[47] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_48 bl[48] br[48] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_49 bl[49] br[49] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_50 bl[50] br[50] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_51 bl[51] br[51] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_52 bl[52] br[52] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_53 bl[53] br[53] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_54 bl[54] br[54] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_55 bl[55] br[55] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_56 bl[56] br[56] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_57 bl[57] br[57] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_58 bl[58] br[58] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_59 bl[59] br[59] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_60 bl[60] br[60] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_61 bl[61] br[61] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_62 bl[62] br[62] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_63 bl[63] br[63] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_45_0 bl[0] br[0] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_1 bl[1] br[1] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_2 bl[2] br[2] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_3 bl[3] br[3] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_4 bl[4] br[4] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_5 bl[5] br[5] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_6 bl[6] br[6] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_7 bl[7] br[7] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_8 bl[8] br[8] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_9 bl[9] br[9] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_10 bl[10] br[10] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_11 bl[11] br[11] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_12 bl[12] br[12] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_13 bl[13] br[13] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_14 bl[14] br[14] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_15 bl[15] br[15] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_16 bl[16] br[16] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_17 bl[17] br[17] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_18 bl[18] br[18] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_19 bl[19] br[19] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_20 bl[20] br[20] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_21 bl[21] br[21] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_22 bl[22] br[22] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_23 bl[23] br[23] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_24 bl[24] br[24] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_25 bl[25] br[25] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_26 bl[26] br[26] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_27 bl[27] br[27] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_28 bl[28] br[28] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_29 bl[29] br[29] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_30 bl[30] br[30] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_31 bl[31] br[31] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_32 bl[32] br[32] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_33 bl[33] br[33] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_34 bl[34] br[34] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_35 bl[35] br[35] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_36 bl[36] br[36] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_37 bl[37] br[37] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_38 bl[38] br[38] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_39 bl[39] br[39] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_40 bl[40] br[40] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_41 bl[41] br[41] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_42 bl[42] br[42] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_43 bl[43] br[43] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_44 bl[44] br[44] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_45 bl[45] br[45] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_46 bl[46] br[46] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_47 bl[47] br[47] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_48 bl[48] br[48] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_49 bl[49] br[49] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_50 bl[50] br[50] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_51 bl[51] br[51] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_52 bl[52] br[52] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_53 bl[53] br[53] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_54 bl[54] br[54] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_55 bl[55] br[55] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_56 bl[56] br[56] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_57 bl[57] br[57] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_58 bl[58] br[58] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_59 bl[59] br[59] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_60 bl[60] br[60] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_61 bl[61] br[61] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_62 bl[62] br[62] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_63 bl[63] br[63] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_46_0 bl[0] br[0] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_1 bl[1] br[1] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_2 bl[2] br[2] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_3 bl[3] br[3] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_4 bl[4] br[4] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_5 bl[5] br[5] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_6 bl[6] br[6] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_7 bl[7] br[7] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_8 bl[8] br[8] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_9 bl[9] br[9] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_10 bl[10] br[10] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_11 bl[11] br[11] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_12 bl[12] br[12] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_13 bl[13] br[13] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_14 bl[14] br[14] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_15 bl[15] br[15] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_16 bl[16] br[16] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_17 bl[17] br[17] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_18 bl[18] br[18] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_19 bl[19] br[19] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_20 bl[20] br[20] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_21 bl[21] br[21] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_22 bl[22] br[22] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_23 bl[23] br[23] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_24 bl[24] br[24] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_25 bl[25] br[25] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_26 bl[26] br[26] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_27 bl[27] br[27] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_28 bl[28] br[28] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_29 bl[29] br[29] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_30 bl[30] br[30] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_31 bl[31] br[31] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_32 bl[32] br[32] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_33 bl[33] br[33] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_34 bl[34] br[34] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_35 bl[35] br[35] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_36 bl[36] br[36] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_37 bl[37] br[37] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_38 bl[38] br[38] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_39 bl[39] br[39] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_40 bl[40] br[40] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_41 bl[41] br[41] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_42 bl[42] br[42] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_43 bl[43] br[43] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_44 bl[44] br[44] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_45 bl[45] br[45] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_46 bl[46] br[46] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_47 bl[47] br[47] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_48 bl[48] br[48] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_49 bl[49] br[49] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_50 bl[50] br[50] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_51 bl[51] br[51] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_52 bl[52] br[52] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_53 bl[53] br[53] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_54 bl[54] br[54] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_55 bl[55] br[55] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_56 bl[56] br[56] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_57 bl[57] br[57] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_58 bl[58] br[58] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_59 bl[59] br[59] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_60 bl[60] br[60] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_61 bl[61] br[61] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_62 bl[62] br[62] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_63 bl[63] br[63] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_47_0 bl[0] br[0] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_1 bl[1] br[1] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_2 bl[2] br[2] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_3 bl[3] br[3] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_4 bl[4] br[4] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_5 bl[5] br[5] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_6 bl[6] br[6] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_7 bl[7] br[7] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_8 bl[8] br[8] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_9 bl[9] br[9] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_10 bl[10] br[10] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_11 bl[11] br[11] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_12 bl[12] br[12] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_13 bl[13] br[13] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_14 bl[14] br[14] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_15 bl[15] br[15] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_16 bl[16] br[16] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_17 bl[17] br[17] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_18 bl[18] br[18] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_19 bl[19] br[19] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_20 bl[20] br[20] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_21 bl[21] br[21] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_22 bl[22] br[22] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_23 bl[23] br[23] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_24 bl[24] br[24] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_25 bl[25] br[25] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_26 bl[26] br[26] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_27 bl[27] br[27] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_28 bl[28] br[28] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_29 bl[29] br[29] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_30 bl[30] br[30] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_31 bl[31] br[31] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_32 bl[32] br[32] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_33 bl[33] br[33] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_34 bl[34] br[34] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_35 bl[35] br[35] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_36 bl[36] br[36] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_37 bl[37] br[37] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_38 bl[38] br[38] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_39 bl[39] br[39] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_40 bl[40] br[40] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_41 bl[41] br[41] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_42 bl[42] br[42] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_43 bl[43] br[43] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_44 bl[44] br[44] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_45 bl[45] br[45] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_46 bl[46] br[46] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_47 bl[47] br[47] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_48 bl[48] br[48] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_49 bl[49] br[49] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_50 bl[50] br[50] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_51 bl[51] br[51] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_52 bl[52] br[52] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_53 bl[53] br[53] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_54 bl[54] br[54] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_55 bl[55] br[55] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_56 bl[56] br[56] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_57 bl[57] br[57] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_58 bl[58] br[58] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_59 bl[59] br[59] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_60 bl[60] br[60] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_61 bl[61] br[61] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_62 bl[62] br[62] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_63 bl[63] br[63] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_48_0 bl[0] br[0] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_1 bl[1] br[1] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_2 bl[2] br[2] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_3 bl[3] br[3] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_4 bl[4] br[4] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_5 bl[5] br[5] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_6 bl[6] br[6] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_7 bl[7] br[7] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_8 bl[8] br[8] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_9 bl[9] br[9] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_10 bl[10] br[10] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_11 bl[11] br[11] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_12 bl[12] br[12] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_13 bl[13] br[13] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_14 bl[14] br[14] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_15 bl[15] br[15] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_16 bl[16] br[16] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_17 bl[17] br[17] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_18 bl[18] br[18] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_19 bl[19] br[19] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_20 bl[20] br[20] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_21 bl[21] br[21] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_22 bl[22] br[22] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_23 bl[23] br[23] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_24 bl[24] br[24] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_25 bl[25] br[25] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_26 bl[26] br[26] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_27 bl[27] br[27] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_28 bl[28] br[28] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_29 bl[29] br[29] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_30 bl[30] br[30] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_31 bl[31] br[31] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_32 bl[32] br[32] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_33 bl[33] br[33] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_34 bl[34] br[34] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_35 bl[35] br[35] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_36 bl[36] br[36] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_37 bl[37] br[37] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_38 bl[38] br[38] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_39 bl[39] br[39] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_40 bl[40] br[40] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_41 bl[41] br[41] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_42 bl[42] br[42] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_43 bl[43] br[43] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_44 bl[44] br[44] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_45 bl[45] br[45] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_46 bl[46] br[46] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_47 bl[47] br[47] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_48 bl[48] br[48] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_49 bl[49] br[49] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_50 bl[50] br[50] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_51 bl[51] br[51] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_52 bl[52] br[52] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_53 bl[53] br[53] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_54 bl[54] br[54] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_55 bl[55] br[55] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_56 bl[56] br[56] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_57 bl[57] br[57] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_58 bl[58] br[58] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_59 bl[59] br[59] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_60 bl[60] br[60] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_61 bl[61] br[61] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_62 bl[62] br[62] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_63 bl[63] br[63] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_49_0 bl[0] br[0] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_1 bl[1] br[1] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_2 bl[2] br[2] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_3 bl[3] br[3] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_4 bl[4] br[4] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_5 bl[5] br[5] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_6 bl[6] br[6] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_7 bl[7] br[7] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_8 bl[8] br[8] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_9 bl[9] br[9] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_10 bl[10] br[10] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_11 bl[11] br[11] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_12 bl[12] br[12] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_13 bl[13] br[13] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_14 bl[14] br[14] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_15 bl[15] br[15] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_16 bl[16] br[16] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_17 bl[17] br[17] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_18 bl[18] br[18] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_19 bl[19] br[19] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_20 bl[20] br[20] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_21 bl[21] br[21] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_22 bl[22] br[22] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_23 bl[23] br[23] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_24 bl[24] br[24] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_25 bl[25] br[25] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_26 bl[26] br[26] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_27 bl[27] br[27] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_28 bl[28] br[28] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_29 bl[29] br[29] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_30 bl[30] br[30] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_31 bl[31] br[31] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_32 bl[32] br[32] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_33 bl[33] br[33] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_34 bl[34] br[34] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_35 bl[35] br[35] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_36 bl[36] br[36] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_37 bl[37] br[37] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_38 bl[38] br[38] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_39 bl[39] br[39] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_40 bl[40] br[40] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_41 bl[41] br[41] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_42 bl[42] br[42] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_43 bl[43] br[43] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_44 bl[44] br[44] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_45 bl[45] br[45] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_46 bl[46] br[46] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_47 bl[47] br[47] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_48 bl[48] br[48] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_49 bl[49] br[49] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_50 bl[50] br[50] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_51 bl[51] br[51] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_52 bl[52] br[52] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_53 bl[53] br[53] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_54 bl[54] br[54] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_55 bl[55] br[55] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_56 bl[56] br[56] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_57 bl[57] br[57] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_58 bl[58] br[58] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_59 bl[59] br[59] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_60 bl[60] br[60] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_61 bl[61] br[61] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_62 bl[62] br[62] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_63 bl[63] br[63] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_50_0 bl[0] br[0] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_1 bl[1] br[1] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_2 bl[2] br[2] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_3 bl[3] br[3] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_4 bl[4] br[4] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_5 bl[5] br[5] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_6 bl[6] br[6] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_7 bl[7] br[7] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_8 bl[8] br[8] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_9 bl[9] br[9] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_10 bl[10] br[10] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_11 bl[11] br[11] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_12 bl[12] br[12] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_13 bl[13] br[13] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_14 bl[14] br[14] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_15 bl[15] br[15] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_16 bl[16] br[16] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_17 bl[17] br[17] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_18 bl[18] br[18] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_19 bl[19] br[19] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_20 bl[20] br[20] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_21 bl[21] br[21] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_22 bl[22] br[22] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_23 bl[23] br[23] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_24 bl[24] br[24] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_25 bl[25] br[25] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_26 bl[26] br[26] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_27 bl[27] br[27] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_28 bl[28] br[28] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_29 bl[29] br[29] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_30 bl[30] br[30] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_31 bl[31] br[31] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_32 bl[32] br[32] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_33 bl[33] br[33] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_34 bl[34] br[34] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_35 bl[35] br[35] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_36 bl[36] br[36] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_37 bl[37] br[37] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_38 bl[38] br[38] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_39 bl[39] br[39] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_40 bl[40] br[40] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_41 bl[41] br[41] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_42 bl[42] br[42] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_43 bl[43] br[43] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_44 bl[44] br[44] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_45 bl[45] br[45] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_46 bl[46] br[46] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_47 bl[47] br[47] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_48 bl[48] br[48] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_49 bl[49] br[49] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_50 bl[50] br[50] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_51 bl[51] br[51] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_52 bl[52] br[52] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_53 bl[53] br[53] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_54 bl[54] br[54] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_55 bl[55] br[55] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_56 bl[56] br[56] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_57 bl[57] br[57] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_58 bl[58] br[58] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_59 bl[59] br[59] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_60 bl[60] br[60] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_61 bl[61] br[61] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_62 bl[62] br[62] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_63 bl[63] br[63] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_51_0 bl[0] br[0] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_1 bl[1] br[1] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_2 bl[2] br[2] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_3 bl[3] br[3] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_4 bl[4] br[4] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_5 bl[5] br[5] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_6 bl[6] br[6] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_7 bl[7] br[7] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_8 bl[8] br[8] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_9 bl[9] br[9] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_10 bl[10] br[10] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_11 bl[11] br[11] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_12 bl[12] br[12] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_13 bl[13] br[13] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_14 bl[14] br[14] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_15 bl[15] br[15] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_16 bl[16] br[16] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_17 bl[17] br[17] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_18 bl[18] br[18] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_19 bl[19] br[19] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_20 bl[20] br[20] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_21 bl[21] br[21] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_22 bl[22] br[22] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_23 bl[23] br[23] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_24 bl[24] br[24] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_25 bl[25] br[25] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_26 bl[26] br[26] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_27 bl[27] br[27] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_28 bl[28] br[28] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_29 bl[29] br[29] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_30 bl[30] br[30] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_31 bl[31] br[31] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_32 bl[32] br[32] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_33 bl[33] br[33] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_34 bl[34] br[34] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_35 bl[35] br[35] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_36 bl[36] br[36] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_37 bl[37] br[37] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_38 bl[38] br[38] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_39 bl[39] br[39] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_40 bl[40] br[40] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_41 bl[41] br[41] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_42 bl[42] br[42] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_43 bl[43] br[43] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_44 bl[44] br[44] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_45 bl[45] br[45] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_46 bl[46] br[46] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_47 bl[47] br[47] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_48 bl[48] br[48] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_49 bl[49] br[49] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_50 bl[50] br[50] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_51 bl[51] br[51] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_52 bl[52] br[52] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_53 bl[53] br[53] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_54 bl[54] br[54] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_55 bl[55] br[55] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_56 bl[56] br[56] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_57 bl[57] br[57] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_58 bl[58] br[58] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_59 bl[59] br[59] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_60 bl[60] br[60] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_61 bl[61] br[61] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_62 bl[62] br[62] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_63 bl[63] br[63] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_52_0 bl[0] br[0] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_1 bl[1] br[1] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_2 bl[2] br[2] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_3 bl[3] br[3] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_4 bl[4] br[4] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_5 bl[5] br[5] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_6 bl[6] br[6] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_7 bl[7] br[7] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_8 bl[8] br[8] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_9 bl[9] br[9] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_10 bl[10] br[10] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_11 bl[11] br[11] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_12 bl[12] br[12] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_13 bl[13] br[13] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_14 bl[14] br[14] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_15 bl[15] br[15] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_16 bl[16] br[16] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_17 bl[17] br[17] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_18 bl[18] br[18] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_19 bl[19] br[19] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_20 bl[20] br[20] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_21 bl[21] br[21] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_22 bl[22] br[22] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_23 bl[23] br[23] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_24 bl[24] br[24] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_25 bl[25] br[25] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_26 bl[26] br[26] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_27 bl[27] br[27] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_28 bl[28] br[28] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_29 bl[29] br[29] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_30 bl[30] br[30] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_31 bl[31] br[31] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_32 bl[32] br[32] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_33 bl[33] br[33] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_34 bl[34] br[34] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_35 bl[35] br[35] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_36 bl[36] br[36] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_37 bl[37] br[37] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_38 bl[38] br[38] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_39 bl[39] br[39] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_40 bl[40] br[40] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_41 bl[41] br[41] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_42 bl[42] br[42] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_43 bl[43] br[43] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_44 bl[44] br[44] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_45 bl[45] br[45] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_46 bl[46] br[46] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_47 bl[47] br[47] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_48 bl[48] br[48] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_49 bl[49] br[49] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_50 bl[50] br[50] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_51 bl[51] br[51] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_52 bl[52] br[52] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_53 bl[53] br[53] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_54 bl[54] br[54] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_55 bl[55] br[55] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_56 bl[56] br[56] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_57 bl[57] br[57] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_58 bl[58] br[58] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_59 bl[59] br[59] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_60 bl[60] br[60] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_61 bl[61] br[61] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_62 bl[62] br[62] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_63 bl[63] br[63] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_53_0 bl[0] br[0] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_1 bl[1] br[1] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_2 bl[2] br[2] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_3 bl[3] br[3] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_4 bl[4] br[4] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_5 bl[5] br[5] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_6 bl[6] br[6] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_7 bl[7] br[7] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_8 bl[8] br[8] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_9 bl[9] br[9] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_10 bl[10] br[10] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_11 bl[11] br[11] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_12 bl[12] br[12] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_13 bl[13] br[13] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_14 bl[14] br[14] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_15 bl[15] br[15] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_16 bl[16] br[16] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_17 bl[17] br[17] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_18 bl[18] br[18] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_19 bl[19] br[19] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_20 bl[20] br[20] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_21 bl[21] br[21] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_22 bl[22] br[22] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_23 bl[23] br[23] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_24 bl[24] br[24] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_25 bl[25] br[25] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_26 bl[26] br[26] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_27 bl[27] br[27] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_28 bl[28] br[28] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_29 bl[29] br[29] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_30 bl[30] br[30] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_31 bl[31] br[31] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_32 bl[32] br[32] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_33 bl[33] br[33] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_34 bl[34] br[34] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_35 bl[35] br[35] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_36 bl[36] br[36] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_37 bl[37] br[37] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_38 bl[38] br[38] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_39 bl[39] br[39] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_40 bl[40] br[40] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_41 bl[41] br[41] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_42 bl[42] br[42] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_43 bl[43] br[43] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_44 bl[44] br[44] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_45 bl[45] br[45] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_46 bl[46] br[46] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_47 bl[47] br[47] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_48 bl[48] br[48] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_49 bl[49] br[49] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_50 bl[50] br[50] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_51 bl[51] br[51] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_52 bl[52] br[52] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_53 bl[53] br[53] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_54 bl[54] br[54] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_55 bl[55] br[55] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_56 bl[56] br[56] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_57 bl[57] br[57] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_58 bl[58] br[58] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_59 bl[59] br[59] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_60 bl[60] br[60] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_61 bl[61] br[61] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_62 bl[62] br[62] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_63 bl[63] br[63] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_54_0 bl[0] br[0] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_1 bl[1] br[1] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_2 bl[2] br[2] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_3 bl[3] br[3] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_4 bl[4] br[4] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_5 bl[5] br[5] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_6 bl[6] br[6] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_7 bl[7] br[7] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_8 bl[8] br[8] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_9 bl[9] br[9] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_10 bl[10] br[10] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_11 bl[11] br[11] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_12 bl[12] br[12] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_13 bl[13] br[13] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_14 bl[14] br[14] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_15 bl[15] br[15] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_16 bl[16] br[16] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_17 bl[17] br[17] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_18 bl[18] br[18] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_19 bl[19] br[19] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_20 bl[20] br[20] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_21 bl[21] br[21] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_22 bl[22] br[22] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_23 bl[23] br[23] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_24 bl[24] br[24] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_25 bl[25] br[25] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_26 bl[26] br[26] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_27 bl[27] br[27] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_28 bl[28] br[28] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_29 bl[29] br[29] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_30 bl[30] br[30] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_31 bl[31] br[31] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_32 bl[32] br[32] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_33 bl[33] br[33] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_34 bl[34] br[34] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_35 bl[35] br[35] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_36 bl[36] br[36] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_37 bl[37] br[37] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_38 bl[38] br[38] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_39 bl[39] br[39] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_40 bl[40] br[40] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_41 bl[41] br[41] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_42 bl[42] br[42] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_43 bl[43] br[43] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_44 bl[44] br[44] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_45 bl[45] br[45] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_46 bl[46] br[46] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_47 bl[47] br[47] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_48 bl[48] br[48] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_49 bl[49] br[49] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_50 bl[50] br[50] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_51 bl[51] br[51] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_52 bl[52] br[52] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_53 bl[53] br[53] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_54 bl[54] br[54] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_55 bl[55] br[55] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_56 bl[56] br[56] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_57 bl[57] br[57] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_58 bl[58] br[58] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_59 bl[59] br[59] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_60 bl[60] br[60] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_61 bl[61] br[61] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_62 bl[62] br[62] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_63 bl[63] br[63] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_55_0 bl[0] br[0] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_1 bl[1] br[1] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_2 bl[2] br[2] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_3 bl[3] br[3] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_4 bl[4] br[4] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_5 bl[5] br[5] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_6 bl[6] br[6] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_7 bl[7] br[7] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_8 bl[8] br[8] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_9 bl[9] br[9] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_10 bl[10] br[10] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_11 bl[11] br[11] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_12 bl[12] br[12] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_13 bl[13] br[13] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_14 bl[14] br[14] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_15 bl[15] br[15] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_16 bl[16] br[16] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_17 bl[17] br[17] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_18 bl[18] br[18] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_19 bl[19] br[19] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_20 bl[20] br[20] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_21 bl[21] br[21] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_22 bl[22] br[22] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_23 bl[23] br[23] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_24 bl[24] br[24] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_25 bl[25] br[25] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_26 bl[26] br[26] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_27 bl[27] br[27] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_28 bl[28] br[28] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_29 bl[29] br[29] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_30 bl[30] br[30] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_31 bl[31] br[31] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_32 bl[32] br[32] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_33 bl[33] br[33] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_34 bl[34] br[34] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_35 bl[35] br[35] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_36 bl[36] br[36] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_37 bl[37] br[37] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_38 bl[38] br[38] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_39 bl[39] br[39] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_40 bl[40] br[40] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_41 bl[41] br[41] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_42 bl[42] br[42] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_43 bl[43] br[43] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_44 bl[44] br[44] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_45 bl[45] br[45] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_46 bl[46] br[46] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_47 bl[47] br[47] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_48 bl[48] br[48] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_49 bl[49] br[49] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_50 bl[50] br[50] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_51 bl[51] br[51] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_52 bl[52] br[52] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_53 bl[53] br[53] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_54 bl[54] br[54] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_55 bl[55] br[55] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_56 bl[56] br[56] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_57 bl[57] br[57] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_58 bl[58] br[58] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_59 bl[59] br[59] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_60 bl[60] br[60] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_61 bl[61] br[61] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_62 bl[62] br[62] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_63 bl[63] br[63] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_56_0 bl[0] br[0] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_1 bl[1] br[1] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_2 bl[2] br[2] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_3 bl[3] br[3] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_4 bl[4] br[4] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_5 bl[5] br[5] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_6 bl[6] br[6] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_7 bl[7] br[7] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_8 bl[8] br[8] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_9 bl[9] br[9] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_10 bl[10] br[10] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_11 bl[11] br[11] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_12 bl[12] br[12] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_13 bl[13] br[13] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_14 bl[14] br[14] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_15 bl[15] br[15] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_16 bl[16] br[16] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_17 bl[17] br[17] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_18 bl[18] br[18] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_19 bl[19] br[19] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_20 bl[20] br[20] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_21 bl[21] br[21] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_22 bl[22] br[22] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_23 bl[23] br[23] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_24 bl[24] br[24] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_25 bl[25] br[25] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_26 bl[26] br[26] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_27 bl[27] br[27] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_28 bl[28] br[28] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_29 bl[29] br[29] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_30 bl[30] br[30] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_31 bl[31] br[31] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_32 bl[32] br[32] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_33 bl[33] br[33] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_34 bl[34] br[34] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_35 bl[35] br[35] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_36 bl[36] br[36] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_37 bl[37] br[37] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_38 bl[38] br[38] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_39 bl[39] br[39] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_40 bl[40] br[40] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_41 bl[41] br[41] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_42 bl[42] br[42] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_43 bl[43] br[43] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_44 bl[44] br[44] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_45 bl[45] br[45] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_46 bl[46] br[46] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_47 bl[47] br[47] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_48 bl[48] br[48] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_49 bl[49] br[49] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_50 bl[50] br[50] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_51 bl[51] br[51] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_52 bl[52] br[52] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_53 bl[53] br[53] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_54 bl[54] br[54] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_55 bl[55] br[55] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_56 bl[56] br[56] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_57 bl[57] br[57] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_58 bl[58] br[58] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_59 bl[59] br[59] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_60 bl[60] br[60] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_61 bl[61] br[61] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_62 bl[62] br[62] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_63 bl[63] br[63] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_57_0 bl[0] br[0] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_1 bl[1] br[1] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_2 bl[2] br[2] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_3 bl[3] br[3] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_4 bl[4] br[4] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_5 bl[5] br[5] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_6 bl[6] br[6] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_7 bl[7] br[7] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_8 bl[8] br[8] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_9 bl[9] br[9] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_10 bl[10] br[10] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_11 bl[11] br[11] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_12 bl[12] br[12] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_13 bl[13] br[13] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_14 bl[14] br[14] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_15 bl[15] br[15] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_16 bl[16] br[16] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_17 bl[17] br[17] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_18 bl[18] br[18] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_19 bl[19] br[19] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_20 bl[20] br[20] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_21 bl[21] br[21] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_22 bl[22] br[22] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_23 bl[23] br[23] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_24 bl[24] br[24] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_25 bl[25] br[25] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_26 bl[26] br[26] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_27 bl[27] br[27] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_28 bl[28] br[28] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_29 bl[29] br[29] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_30 bl[30] br[30] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_31 bl[31] br[31] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_32 bl[32] br[32] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_33 bl[33] br[33] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_34 bl[34] br[34] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_35 bl[35] br[35] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_36 bl[36] br[36] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_37 bl[37] br[37] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_38 bl[38] br[38] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_39 bl[39] br[39] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_40 bl[40] br[40] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_41 bl[41] br[41] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_42 bl[42] br[42] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_43 bl[43] br[43] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_44 bl[44] br[44] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_45 bl[45] br[45] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_46 bl[46] br[46] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_47 bl[47] br[47] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_48 bl[48] br[48] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_49 bl[49] br[49] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_50 bl[50] br[50] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_51 bl[51] br[51] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_52 bl[52] br[52] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_53 bl[53] br[53] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_54 bl[54] br[54] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_55 bl[55] br[55] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_56 bl[56] br[56] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_57 bl[57] br[57] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_58 bl[58] br[58] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_59 bl[59] br[59] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_60 bl[60] br[60] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_61 bl[61] br[61] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_62 bl[62] br[62] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_63 bl[63] br[63] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_58_0 bl[0] br[0] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_1 bl[1] br[1] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_2 bl[2] br[2] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_3 bl[3] br[3] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_4 bl[4] br[4] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_5 bl[5] br[5] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_6 bl[6] br[6] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_7 bl[7] br[7] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_8 bl[8] br[8] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_9 bl[9] br[9] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_10 bl[10] br[10] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_11 bl[11] br[11] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_12 bl[12] br[12] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_13 bl[13] br[13] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_14 bl[14] br[14] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_15 bl[15] br[15] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_16 bl[16] br[16] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_17 bl[17] br[17] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_18 bl[18] br[18] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_19 bl[19] br[19] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_20 bl[20] br[20] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_21 bl[21] br[21] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_22 bl[22] br[22] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_23 bl[23] br[23] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_24 bl[24] br[24] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_25 bl[25] br[25] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_26 bl[26] br[26] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_27 bl[27] br[27] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_28 bl[28] br[28] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_29 bl[29] br[29] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_30 bl[30] br[30] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_31 bl[31] br[31] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_32 bl[32] br[32] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_33 bl[33] br[33] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_34 bl[34] br[34] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_35 bl[35] br[35] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_36 bl[36] br[36] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_37 bl[37] br[37] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_38 bl[38] br[38] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_39 bl[39] br[39] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_40 bl[40] br[40] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_41 bl[41] br[41] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_42 bl[42] br[42] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_43 bl[43] br[43] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_44 bl[44] br[44] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_45 bl[45] br[45] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_46 bl[46] br[46] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_47 bl[47] br[47] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_48 bl[48] br[48] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_49 bl[49] br[49] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_50 bl[50] br[50] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_51 bl[51] br[51] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_52 bl[52] br[52] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_53 bl[53] br[53] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_54 bl[54] br[54] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_55 bl[55] br[55] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_56 bl[56] br[56] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_57 bl[57] br[57] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_58 bl[58] br[58] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_59 bl[59] br[59] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_60 bl[60] br[60] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_61 bl[61] br[61] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_62 bl[62] br[62] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_63 bl[63] br[63] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_59_0 bl[0] br[0] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_1 bl[1] br[1] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_2 bl[2] br[2] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_3 bl[3] br[3] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_4 bl[4] br[4] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_5 bl[5] br[5] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_6 bl[6] br[6] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_7 bl[7] br[7] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_8 bl[8] br[8] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_9 bl[9] br[9] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_10 bl[10] br[10] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_11 bl[11] br[11] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_12 bl[12] br[12] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_13 bl[13] br[13] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_14 bl[14] br[14] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_15 bl[15] br[15] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_16 bl[16] br[16] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_17 bl[17] br[17] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_18 bl[18] br[18] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_19 bl[19] br[19] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_20 bl[20] br[20] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_21 bl[21] br[21] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_22 bl[22] br[22] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_23 bl[23] br[23] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_24 bl[24] br[24] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_25 bl[25] br[25] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_26 bl[26] br[26] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_27 bl[27] br[27] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_28 bl[28] br[28] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_29 bl[29] br[29] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_30 bl[30] br[30] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_31 bl[31] br[31] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_32 bl[32] br[32] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_33 bl[33] br[33] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_34 bl[34] br[34] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_35 bl[35] br[35] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_36 bl[36] br[36] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_37 bl[37] br[37] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_38 bl[38] br[38] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_39 bl[39] br[39] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_40 bl[40] br[40] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_41 bl[41] br[41] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_42 bl[42] br[42] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_43 bl[43] br[43] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_44 bl[44] br[44] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_45 bl[45] br[45] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_46 bl[46] br[46] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_47 bl[47] br[47] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_48 bl[48] br[48] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_49 bl[49] br[49] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_50 bl[50] br[50] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_51 bl[51] br[51] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_52 bl[52] br[52] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_53 bl[53] br[53] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_54 bl[54] br[54] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_55 bl[55] br[55] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_56 bl[56] br[56] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_57 bl[57] br[57] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_58 bl[58] br[58] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_59 bl[59] br[59] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_60 bl[60] br[60] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_61 bl[61] br[61] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_62 bl[62] br[62] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_63 bl[63] br[63] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_60_0 bl[0] br[0] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_1 bl[1] br[1] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_2 bl[2] br[2] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_3 bl[3] br[3] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_4 bl[4] br[4] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_5 bl[5] br[5] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_6 bl[6] br[6] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_7 bl[7] br[7] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_8 bl[8] br[8] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_9 bl[9] br[9] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_10 bl[10] br[10] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_11 bl[11] br[11] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_12 bl[12] br[12] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_13 bl[13] br[13] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_14 bl[14] br[14] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_15 bl[15] br[15] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_16 bl[16] br[16] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_17 bl[17] br[17] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_18 bl[18] br[18] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_19 bl[19] br[19] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_20 bl[20] br[20] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_21 bl[21] br[21] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_22 bl[22] br[22] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_23 bl[23] br[23] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_24 bl[24] br[24] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_25 bl[25] br[25] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_26 bl[26] br[26] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_27 bl[27] br[27] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_28 bl[28] br[28] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_29 bl[29] br[29] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_30 bl[30] br[30] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_31 bl[31] br[31] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_32 bl[32] br[32] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_33 bl[33] br[33] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_34 bl[34] br[34] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_35 bl[35] br[35] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_36 bl[36] br[36] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_37 bl[37] br[37] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_38 bl[38] br[38] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_39 bl[39] br[39] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_40 bl[40] br[40] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_41 bl[41] br[41] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_42 bl[42] br[42] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_43 bl[43] br[43] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_44 bl[44] br[44] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_45 bl[45] br[45] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_46 bl[46] br[46] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_47 bl[47] br[47] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_48 bl[48] br[48] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_49 bl[49] br[49] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_50 bl[50] br[50] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_51 bl[51] br[51] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_52 bl[52] br[52] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_53 bl[53] br[53] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_54 bl[54] br[54] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_55 bl[55] br[55] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_56 bl[56] br[56] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_57 bl[57] br[57] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_58 bl[58] br[58] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_59 bl[59] br[59] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_60 bl[60] br[60] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_61 bl[61] br[61] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_62 bl[62] br[62] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_63 bl[63] br[63] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_61_0 bl[0] br[0] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_1 bl[1] br[1] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_2 bl[2] br[2] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_3 bl[3] br[3] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_4 bl[4] br[4] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_5 bl[5] br[5] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_6 bl[6] br[6] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_7 bl[7] br[7] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_8 bl[8] br[8] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_9 bl[9] br[9] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_10 bl[10] br[10] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_11 bl[11] br[11] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_12 bl[12] br[12] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_13 bl[13] br[13] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_14 bl[14] br[14] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_15 bl[15] br[15] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_16 bl[16] br[16] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_17 bl[17] br[17] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_18 bl[18] br[18] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_19 bl[19] br[19] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_20 bl[20] br[20] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_21 bl[21] br[21] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_22 bl[22] br[22] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_23 bl[23] br[23] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_24 bl[24] br[24] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_25 bl[25] br[25] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_26 bl[26] br[26] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_27 bl[27] br[27] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_28 bl[28] br[28] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_29 bl[29] br[29] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_30 bl[30] br[30] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_31 bl[31] br[31] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_32 bl[32] br[32] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_33 bl[33] br[33] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_34 bl[34] br[34] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_35 bl[35] br[35] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_36 bl[36] br[36] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_37 bl[37] br[37] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_38 bl[38] br[38] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_39 bl[39] br[39] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_40 bl[40] br[40] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_41 bl[41] br[41] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_42 bl[42] br[42] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_43 bl[43] br[43] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_44 bl[44] br[44] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_45 bl[45] br[45] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_46 bl[46] br[46] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_47 bl[47] br[47] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_48 bl[48] br[48] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_49 bl[49] br[49] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_50 bl[50] br[50] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_51 bl[51] br[51] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_52 bl[52] br[52] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_53 bl[53] br[53] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_54 bl[54] br[54] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_55 bl[55] br[55] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_56 bl[56] br[56] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_57 bl[57] br[57] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_58 bl[58] br[58] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_59 bl[59] br[59] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_60 bl[60] br[60] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_61 bl[61] br[61] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_62 bl[62] br[62] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_63 bl[63] br[63] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_62_0 bl[0] br[0] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_1 bl[1] br[1] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_2 bl[2] br[2] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_3 bl[3] br[3] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_4 bl[4] br[4] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_5 bl[5] br[5] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_6 bl[6] br[6] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_7 bl[7] br[7] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_8 bl[8] br[8] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_9 bl[9] br[9] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_10 bl[10] br[10] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_11 bl[11] br[11] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_12 bl[12] br[12] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_13 bl[13] br[13] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_14 bl[14] br[14] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_15 bl[15] br[15] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_16 bl[16] br[16] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_17 bl[17] br[17] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_18 bl[18] br[18] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_19 bl[19] br[19] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_20 bl[20] br[20] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_21 bl[21] br[21] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_22 bl[22] br[22] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_23 bl[23] br[23] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_24 bl[24] br[24] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_25 bl[25] br[25] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_26 bl[26] br[26] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_27 bl[27] br[27] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_28 bl[28] br[28] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_29 bl[29] br[29] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_30 bl[30] br[30] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_31 bl[31] br[31] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_32 bl[32] br[32] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_33 bl[33] br[33] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_34 bl[34] br[34] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_35 bl[35] br[35] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_36 bl[36] br[36] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_37 bl[37] br[37] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_38 bl[38] br[38] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_39 bl[39] br[39] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_40 bl[40] br[40] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_41 bl[41] br[41] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_42 bl[42] br[42] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_43 bl[43] br[43] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_44 bl[44] br[44] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_45 bl[45] br[45] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_46 bl[46] br[46] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_47 bl[47] br[47] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_48 bl[48] br[48] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_49 bl[49] br[49] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_50 bl[50] br[50] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_51 bl[51] br[51] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_52 bl[52] br[52] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_53 bl[53] br[53] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_54 bl[54] br[54] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_55 bl[55] br[55] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_56 bl[56] br[56] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_57 bl[57] br[57] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_58 bl[58] br[58] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_59 bl[59] br[59] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_60 bl[60] br[60] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_61 bl[61] br[61] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_62 bl[62] br[62] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_63 bl[63] br[63] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_63_0 bl[0] br[0] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_1 bl[1] br[1] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_2 bl[2] br[2] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_3 bl[3] br[3] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_4 bl[4] br[4] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_5 bl[5] br[5] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_6 bl[6] br[6] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_7 bl[7] br[7] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_8 bl[8] br[8] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_9 bl[9] br[9] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_10 bl[10] br[10] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_11 bl[11] br[11] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_12 bl[12] br[12] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_13 bl[13] br[13] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_14 bl[14] br[14] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_15 bl[15] br[15] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_16 bl[16] br[16] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_17 bl[17] br[17] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_18 bl[18] br[18] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_19 bl[19] br[19] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_20 bl[20] br[20] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_21 bl[21] br[21] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_22 bl[22] br[22] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_23 bl[23] br[23] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_24 bl[24] br[24] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_25 bl[25] br[25] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_26 bl[26] br[26] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_27 bl[27] br[27] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_28 bl[28] br[28] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_29 bl[29] br[29] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_30 bl[30] br[30] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_31 bl[31] br[31] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_32 bl[32] br[32] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_33 bl[33] br[33] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_34 bl[34] br[34] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_35 bl[35] br[35] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_36 bl[36] br[36] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_37 bl[37] br[37] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_38 bl[38] br[38] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_39 bl[39] br[39] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_40 bl[40] br[40] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_41 bl[41] br[41] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_42 bl[42] br[42] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_43 bl[43] br[43] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_44 bl[44] br[44] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_45 bl[45] br[45] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_46 bl[46] br[46] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_47 bl[47] br[47] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_48 bl[48] br[48] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_49 bl[49] br[49] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_50 bl[50] br[50] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_51 bl[51] br[51] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_52 bl[52] br[52] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_53 bl[53] br[53] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_54 bl[54] br[54] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_55 bl[55] br[55] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_56 bl[56] br[56] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_57 bl[57] br[57] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_58 bl[58] br[58] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_59 bl[59] br[59] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_60 bl[60] br[60] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_61 bl[61] br[61] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_62 bl[62] br[62] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_63 bl[63] br[63] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_64_0 bl[0] br[0] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_1 bl[1] br[1] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_2 bl[2] br[2] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_3 bl[3] br[3] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_4 bl[4] br[4] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_5 bl[5] br[5] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_6 bl[6] br[6] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_7 bl[7] br[7] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_8 bl[8] br[8] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_9 bl[9] br[9] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_10 bl[10] br[10] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_11 bl[11] br[11] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_12 bl[12] br[12] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_13 bl[13] br[13] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_14 bl[14] br[14] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_15 bl[15] br[15] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_16 bl[16] br[16] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_17 bl[17] br[17] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_18 bl[18] br[18] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_19 bl[19] br[19] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_20 bl[20] br[20] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_21 bl[21] br[21] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_22 bl[22] br[22] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_23 bl[23] br[23] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_24 bl[24] br[24] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_25 bl[25] br[25] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_26 bl[26] br[26] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_27 bl[27] br[27] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_28 bl[28] br[28] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_29 bl[29] br[29] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_30 bl[30] br[30] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_31 bl[31] br[31] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_32 bl[32] br[32] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_33 bl[33] br[33] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_34 bl[34] br[34] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_35 bl[35] br[35] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_36 bl[36] br[36] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_37 bl[37] br[37] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_38 bl[38] br[38] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_39 bl[39] br[39] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_40 bl[40] br[40] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_41 bl[41] br[41] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_42 bl[42] br[42] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_43 bl[43] br[43] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_44 bl[44] br[44] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_45 bl[45] br[45] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_46 bl[46] br[46] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_47 bl[47] br[47] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_48 bl[48] br[48] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_49 bl[49] br[49] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_50 bl[50] br[50] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_51 bl[51] br[51] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_52 bl[52] br[52] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_53 bl[53] br[53] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_54 bl[54] br[54] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_55 bl[55] br[55] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_56 bl[56] br[56] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_57 bl[57] br[57] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_58 bl[58] br[58] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_59 bl[59] br[59] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_60 bl[60] br[60] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_61 bl[61] br[61] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_62 bl[62] br[62] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_63 bl[63] br[63] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_65_0 bl[0] br[0] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_1 bl[1] br[1] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_2 bl[2] br[2] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_3 bl[3] br[3] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_4 bl[4] br[4] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_5 bl[5] br[5] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_6 bl[6] br[6] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_7 bl[7] br[7] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_8 bl[8] br[8] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_9 bl[9] br[9] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_10 bl[10] br[10] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_11 bl[11] br[11] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_12 bl[12] br[12] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_13 bl[13] br[13] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_14 bl[14] br[14] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_15 bl[15] br[15] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_16 bl[16] br[16] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_17 bl[17] br[17] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_18 bl[18] br[18] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_19 bl[19] br[19] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_20 bl[20] br[20] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_21 bl[21] br[21] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_22 bl[22] br[22] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_23 bl[23] br[23] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_24 bl[24] br[24] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_25 bl[25] br[25] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_26 bl[26] br[26] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_27 bl[27] br[27] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_28 bl[28] br[28] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_29 bl[29] br[29] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_30 bl[30] br[30] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_31 bl[31] br[31] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_32 bl[32] br[32] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_33 bl[33] br[33] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_34 bl[34] br[34] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_35 bl[35] br[35] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_36 bl[36] br[36] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_37 bl[37] br[37] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_38 bl[38] br[38] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_39 bl[39] br[39] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_40 bl[40] br[40] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_41 bl[41] br[41] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_42 bl[42] br[42] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_43 bl[43] br[43] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_44 bl[44] br[44] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_45 bl[45] br[45] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_46 bl[46] br[46] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_47 bl[47] br[47] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_48 bl[48] br[48] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_49 bl[49] br[49] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_50 bl[50] br[50] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_51 bl[51] br[51] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_52 bl[52] br[52] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_53 bl[53] br[53] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_54 bl[54] br[54] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_55 bl[55] br[55] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_56 bl[56] br[56] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_57 bl[57] br[57] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_58 bl[58] br[58] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_59 bl[59] br[59] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_60 bl[60] br[60] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_61 bl[61] br[61] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_62 bl[62] br[62] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_63 bl[63] br[63] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_66_0 bl[0] br[0] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_1 bl[1] br[1] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_2 bl[2] br[2] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_3 bl[3] br[3] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_4 bl[4] br[4] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_5 bl[5] br[5] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_6 bl[6] br[6] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_7 bl[7] br[7] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_8 bl[8] br[8] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_9 bl[9] br[9] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_10 bl[10] br[10] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_11 bl[11] br[11] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_12 bl[12] br[12] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_13 bl[13] br[13] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_14 bl[14] br[14] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_15 bl[15] br[15] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_16 bl[16] br[16] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_17 bl[17] br[17] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_18 bl[18] br[18] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_19 bl[19] br[19] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_20 bl[20] br[20] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_21 bl[21] br[21] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_22 bl[22] br[22] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_23 bl[23] br[23] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_24 bl[24] br[24] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_25 bl[25] br[25] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_26 bl[26] br[26] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_27 bl[27] br[27] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_28 bl[28] br[28] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_29 bl[29] br[29] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_30 bl[30] br[30] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_31 bl[31] br[31] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_32 bl[32] br[32] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_33 bl[33] br[33] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_34 bl[34] br[34] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_35 bl[35] br[35] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_36 bl[36] br[36] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_37 bl[37] br[37] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_38 bl[38] br[38] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_39 bl[39] br[39] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_40 bl[40] br[40] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_41 bl[41] br[41] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_42 bl[42] br[42] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_43 bl[43] br[43] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_44 bl[44] br[44] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_45 bl[45] br[45] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_46 bl[46] br[46] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_47 bl[47] br[47] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_48 bl[48] br[48] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_49 bl[49] br[49] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_50 bl[50] br[50] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_51 bl[51] br[51] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_52 bl[52] br[52] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_53 bl[53] br[53] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_54 bl[54] br[54] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_55 bl[55] br[55] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_56 bl[56] br[56] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_57 bl[57] br[57] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_58 bl[58] br[58] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_59 bl[59] br[59] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_60 bl[60] br[60] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_61 bl[61] br[61] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_62 bl[62] br[62] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_63 bl[63] br[63] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_67_0 bl[0] br[0] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_1 bl[1] br[1] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_2 bl[2] br[2] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_3 bl[3] br[3] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_4 bl[4] br[4] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_5 bl[5] br[5] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_6 bl[6] br[6] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_7 bl[7] br[7] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_8 bl[8] br[8] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_9 bl[9] br[9] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_10 bl[10] br[10] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_11 bl[11] br[11] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_12 bl[12] br[12] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_13 bl[13] br[13] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_14 bl[14] br[14] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_15 bl[15] br[15] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_16 bl[16] br[16] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_17 bl[17] br[17] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_18 bl[18] br[18] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_19 bl[19] br[19] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_20 bl[20] br[20] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_21 bl[21] br[21] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_22 bl[22] br[22] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_23 bl[23] br[23] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_24 bl[24] br[24] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_25 bl[25] br[25] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_26 bl[26] br[26] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_27 bl[27] br[27] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_28 bl[28] br[28] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_29 bl[29] br[29] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_30 bl[30] br[30] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_31 bl[31] br[31] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_32 bl[32] br[32] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_33 bl[33] br[33] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_34 bl[34] br[34] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_35 bl[35] br[35] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_36 bl[36] br[36] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_37 bl[37] br[37] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_38 bl[38] br[38] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_39 bl[39] br[39] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_40 bl[40] br[40] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_41 bl[41] br[41] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_42 bl[42] br[42] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_43 bl[43] br[43] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_44 bl[44] br[44] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_45 bl[45] br[45] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_46 bl[46] br[46] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_47 bl[47] br[47] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_48 bl[48] br[48] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_49 bl[49] br[49] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_50 bl[50] br[50] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_51 bl[51] br[51] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_52 bl[52] br[52] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_53 bl[53] br[53] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_54 bl[54] br[54] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_55 bl[55] br[55] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_56 bl[56] br[56] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_57 bl[57] br[57] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_58 bl[58] br[58] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_59 bl[59] br[59] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_60 bl[60] br[60] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_61 bl[61] br[61] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_62 bl[62] br[62] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_63 bl[63] br[63] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_68_0 bl[0] br[0] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_1 bl[1] br[1] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_2 bl[2] br[2] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_3 bl[3] br[3] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_4 bl[4] br[4] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_5 bl[5] br[5] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_6 bl[6] br[6] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_7 bl[7] br[7] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_8 bl[8] br[8] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_9 bl[9] br[9] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_10 bl[10] br[10] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_11 bl[11] br[11] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_12 bl[12] br[12] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_13 bl[13] br[13] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_14 bl[14] br[14] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_15 bl[15] br[15] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_16 bl[16] br[16] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_17 bl[17] br[17] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_18 bl[18] br[18] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_19 bl[19] br[19] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_20 bl[20] br[20] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_21 bl[21] br[21] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_22 bl[22] br[22] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_23 bl[23] br[23] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_24 bl[24] br[24] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_25 bl[25] br[25] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_26 bl[26] br[26] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_27 bl[27] br[27] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_28 bl[28] br[28] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_29 bl[29] br[29] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_30 bl[30] br[30] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_31 bl[31] br[31] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_32 bl[32] br[32] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_33 bl[33] br[33] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_34 bl[34] br[34] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_35 bl[35] br[35] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_36 bl[36] br[36] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_37 bl[37] br[37] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_38 bl[38] br[38] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_39 bl[39] br[39] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_40 bl[40] br[40] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_41 bl[41] br[41] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_42 bl[42] br[42] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_43 bl[43] br[43] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_44 bl[44] br[44] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_45 bl[45] br[45] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_46 bl[46] br[46] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_47 bl[47] br[47] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_48 bl[48] br[48] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_49 bl[49] br[49] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_50 bl[50] br[50] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_51 bl[51] br[51] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_52 bl[52] br[52] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_53 bl[53] br[53] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_54 bl[54] br[54] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_55 bl[55] br[55] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_56 bl[56] br[56] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_57 bl[57] br[57] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_58 bl[58] br[58] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_59 bl[59] br[59] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_60 bl[60] br[60] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_61 bl[61] br[61] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_62 bl[62] br[62] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_63 bl[63] br[63] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_69_0 bl[0] br[0] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_1 bl[1] br[1] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_2 bl[2] br[2] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_3 bl[3] br[3] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_4 bl[4] br[4] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_5 bl[5] br[5] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_6 bl[6] br[6] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_7 bl[7] br[7] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_8 bl[8] br[8] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_9 bl[9] br[9] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_10 bl[10] br[10] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_11 bl[11] br[11] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_12 bl[12] br[12] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_13 bl[13] br[13] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_14 bl[14] br[14] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_15 bl[15] br[15] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_16 bl[16] br[16] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_17 bl[17] br[17] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_18 bl[18] br[18] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_19 bl[19] br[19] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_20 bl[20] br[20] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_21 bl[21] br[21] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_22 bl[22] br[22] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_23 bl[23] br[23] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_24 bl[24] br[24] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_25 bl[25] br[25] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_26 bl[26] br[26] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_27 bl[27] br[27] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_28 bl[28] br[28] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_29 bl[29] br[29] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_30 bl[30] br[30] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_31 bl[31] br[31] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_32 bl[32] br[32] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_33 bl[33] br[33] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_34 bl[34] br[34] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_35 bl[35] br[35] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_36 bl[36] br[36] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_37 bl[37] br[37] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_38 bl[38] br[38] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_39 bl[39] br[39] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_40 bl[40] br[40] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_41 bl[41] br[41] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_42 bl[42] br[42] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_43 bl[43] br[43] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_44 bl[44] br[44] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_45 bl[45] br[45] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_46 bl[46] br[46] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_47 bl[47] br[47] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_48 bl[48] br[48] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_49 bl[49] br[49] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_50 bl[50] br[50] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_51 bl[51] br[51] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_52 bl[52] br[52] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_53 bl[53] br[53] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_54 bl[54] br[54] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_55 bl[55] br[55] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_56 bl[56] br[56] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_57 bl[57] br[57] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_58 bl[58] br[58] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_59 bl[59] br[59] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_60 bl[60] br[60] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_61 bl[61] br[61] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_62 bl[62] br[62] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_63 bl[63] br[63] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_70_0 bl[0] br[0] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_1 bl[1] br[1] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_2 bl[2] br[2] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_3 bl[3] br[3] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_4 bl[4] br[4] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_5 bl[5] br[5] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_6 bl[6] br[6] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_7 bl[7] br[7] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_8 bl[8] br[8] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_9 bl[9] br[9] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_10 bl[10] br[10] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_11 bl[11] br[11] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_12 bl[12] br[12] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_13 bl[13] br[13] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_14 bl[14] br[14] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_15 bl[15] br[15] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_16 bl[16] br[16] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_17 bl[17] br[17] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_18 bl[18] br[18] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_19 bl[19] br[19] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_20 bl[20] br[20] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_21 bl[21] br[21] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_22 bl[22] br[22] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_23 bl[23] br[23] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_24 bl[24] br[24] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_25 bl[25] br[25] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_26 bl[26] br[26] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_27 bl[27] br[27] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_28 bl[28] br[28] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_29 bl[29] br[29] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_30 bl[30] br[30] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_31 bl[31] br[31] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_32 bl[32] br[32] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_33 bl[33] br[33] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_34 bl[34] br[34] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_35 bl[35] br[35] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_36 bl[36] br[36] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_37 bl[37] br[37] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_38 bl[38] br[38] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_39 bl[39] br[39] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_40 bl[40] br[40] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_41 bl[41] br[41] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_42 bl[42] br[42] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_43 bl[43] br[43] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_44 bl[44] br[44] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_45 bl[45] br[45] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_46 bl[46] br[46] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_47 bl[47] br[47] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_48 bl[48] br[48] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_49 bl[49] br[49] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_50 bl[50] br[50] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_51 bl[51] br[51] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_52 bl[52] br[52] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_53 bl[53] br[53] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_54 bl[54] br[54] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_55 bl[55] br[55] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_56 bl[56] br[56] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_57 bl[57] br[57] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_58 bl[58] br[58] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_59 bl[59] br[59] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_60 bl[60] br[60] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_61 bl[61] br[61] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_62 bl[62] br[62] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_63 bl[63] br[63] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_71_0 bl[0] br[0] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_1 bl[1] br[1] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_2 bl[2] br[2] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_3 bl[3] br[3] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_4 bl[4] br[4] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_5 bl[5] br[5] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_6 bl[6] br[6] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_7 bl[7] br[7] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_8 bl[8] br[8] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_9 bl[9] br[9] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_10 bl[10] br[10] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_11 bl[11] br[11] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_12 bl[12] br[12] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_13 bl[13] br[13] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_14 bl[14] br[14] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_15 bl[15] br[15] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_16 bl[16] br[16] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_17 bl[17] br[17] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_18 bl[18] br[18] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_19 bl[19] br[19] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_20 bl[20] br[20] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_21 bl[21] br[21] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_22 bl[22] br[22] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_23 bl[23] br[23] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_24 bl[24] br[24] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_25 bl[25] br[25] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_26 bl[26] br[26] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_27 bl[27] br[27] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_28 bl[28] br[28] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_29 bl[29] br[29] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_30 bl[30] br[30] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_31 bl[31] br[31] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_32 bl[32] br[32] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_33 bl[33] br[33] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_34 bl[34] br[34] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_35 bl[35] br[35] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_36 bl[36] br[36] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_37 bl[37] br[37] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_38 bl[38] br[38] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_39 bl[39] br[39] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_40 bl[40] br[40] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_41 bl[41] br[41] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_42 bl[42] br[42] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_43 bl[43] br[43] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_44 bl[44] br[44] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_45 bl[45] br[45] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_46 bl[46] br[46] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_47 bl[47] br[47] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_48 bl[48] br[48] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_49 bl[49] br[49] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_50 bl[50] br[50] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_51 bl[51] br[51] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_52 bl[52] br[52] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_53 bl[53] br[53] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_54 bl[54] br[54] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_55 bl[55] br[55] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_56 bl[56] br[56] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_57 bl[57] br[57] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_58 bl[58] br[58] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_59 bl[59] br[59] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_60 bl[60] br[60] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_61 bl[61] br[61] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_62 bl[62] br[62] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_63 bl[63] br[63] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_72_0 bl[0] br[0] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_1 bl[1] br[1] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_2 bl[2] br[2] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_3 bl[3] br[3] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_4 bl[4] br[4] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_5 bl[5] br[5] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_6 bl[6] br[6] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_7 bl[7] br[7] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_8 bl[8] br[8] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_9 bl[9] br[9] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_10 bl[10] br[10] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_11 bl[11] br[11] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_12 bl[12] br[12] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_13 bl[13] br[13] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_14 bl[14] br[14] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_15 bl[15] br[15] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_16 bl[16] br[16] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_17 bl[17] br[17] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_18 bl[18] br[18] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_19 bl[19] br[19] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_20 bl[20] br[20] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_21 bl[21] br[21] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_22 bl[22] br[22] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_23 bl[23] br[23] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_24 bl[24] br[24] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_25 bl[25] br[25] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_26 bl[26] br[26] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_27 bl[27] br[27] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_28 bl[28] br[28] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_29 bl[29] br[29] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_30 bl[30] br[30] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_31 bl[31] br[31] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_32 bl[32] br[32] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_33 bl[33] br[33] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_34 bl[34] br[34] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_35 bl[35] br[35] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_36 bl[36] br[36] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_37 bl[37] br[37] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_38 bl[38] br[38] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_39 bl[39] br[39] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_40 bl[40] br[40] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_41 bl[41] br[41] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_42 bl[42] br[42] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_43 bl[43] br[43] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_44 bl[44] br[44] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_45 bl[45] br[45] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_46 bl[46] br[46] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_47 bl[47] br[47] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_48 bl[48] br[48] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_49 bl[49] br[49] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_50 bl[50] br[50] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_51 bl[51] br[51] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_52 bl[52] br[52] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_53 bl[53] br[53] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_54 bl[54] br[54] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_55 bl[55] br[55] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_56 bl[56] br[56] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_57 bl[57] br[57] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_58 bl[58] br[58] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_59 bl[59] br[59] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_60 bl[60] br[60] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_61 bl[61] br[61] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_62 bl[62] br[62] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_63 bl[63] br[63] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_73_0 bl[0] br[0] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_1 bl[1] br[1] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_2 bl[2] br[2] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_3 bl[3] br[3] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_4 bl[4] br[4] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_5 bl[5] br[5] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_6 bl[6] br[6] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_7 bl[7] br[7] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_8 bl[8] br[8] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_9 bl[9] br[9] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_10 bl[10] br[10] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_11 bl[11] br[11] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_12 bl[12] br[12] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_13 bl[13] br[13] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_14 bl[14] br[14] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_15 bl[15] br[15] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_16 bl[16] br[16] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_17 bl[17] br[17] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_18 bl[18] br[18] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_19 bl[19] br[19] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_20 bl[20] br[20] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_21 bl[21] br[21] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_22 bl[22] br[22] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_23 bl[23] br[23] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_24 bl[24] br[24] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_25 bl[25] br[25] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_26 bl[26] br[26] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_27 bl[27] br[27] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_28 bl[28] br[28] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_29 bl[29] br[29] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_30 bl[30] br[30] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_31 bl[31] br[31] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_32 bl[32] br[32] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_33 bl[33] br[33] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_34 bl[34] br[34] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_35 bl[35] br[35] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_36 bl[36] br[36] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_37 bl[37] br[37] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_38 bl[38] br[38] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_39 bl[39] br[39] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_40 bl[40] br[40] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_41 bl[41] br[41] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_42 bl[42] br[42] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_43 bl[43] br[43] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_44 bl[44] br[44] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_45 bl[45] br[45] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_46 bl[46] br[46] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_47 bl[47] br[47] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_48 bl[48] br[48] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_49 bl[49] br[49] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_50 bl[50] br[50] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_51 bl[51] br[51] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_52 bl[52] br[52] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_53 bl[53] br[53] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_54 bl[54] br[54] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_55 bl[55] br[55] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_56 bl[56] br[56] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_57 bl[57] br[57] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_58 bl[58] br[58] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_59 bl[59] br[59] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_60 bl[60] br[60] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_61 bl[61] br[61] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_62 bl[62] br[62] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_63 bl[63] br[63] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_74_0 bl[0] br[0] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_1 bl[1] br[1] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_2 bl[2] br[2] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_3 bl[3] br[3] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_4 bl[4] br[4] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_5 bl[5] br[5] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_6 bl[6] br[6] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_7 bl[7] br[7] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_8 bl[8] br[8] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_9 bl[9] br[9] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_10 bl[10] br[10] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_11 bl[11] br[11] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_12 bl[12] br[12] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_13 bl[13] br[13] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_14 bl[14] br[14] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_15 bl[15] br[15] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_16 bl[16] br[16] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_17 bl[17] br[17] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_18 bl[18] br[18] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_19 bl[19] br[19] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_20 bl[20] br[20] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_21 bl[21] br[21] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_22 bl[22] br[22] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_23 bl[23] br[23] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_24 bl[24] br[24] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_25 bl[25] br[25] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_26 bl[26] br[26] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_27 bl[27] br[27] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_28 bl[28] br[28] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_29 bl[29] br[29] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_30 bl[30] br[30] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_31 bl[31] br[31] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_32 bl[32] br[32] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_33 bl[33] br[33] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_34 bl[34] br[34] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_35 bl[35] br[35] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_36 bl[36] br[36] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_37 bl[37] br[37] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_38 bl[38] br[38] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_39 bl[39] br[39] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_40 bl[40] br[40] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_41 bl[41] br[41] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_42 bl[42] br[42] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_43 bl[43] br[43] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_44 bl[44] br[44] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_45 bl[45] br[45] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_46 bl[46] br[46] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_47 bl[47] br[47] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_48 bl[48] br[48] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_49 bl[49] br[49] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_50 bl[50] br[50] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_51 bl[51] br[51] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_52 bl[52] br[52] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_53 bl[53] br[53] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_54 bl[54] br[54] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_55 bl[55] br[55] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_56 bl[56] br[56] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_57 bl[57] br[57] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_58 bl[58] br[58] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_59 bl[59] br[59] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_60 bl[60] br[60] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_61 bl[61] br[61] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_62 bl[62] br[62] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_63 bl[63] br[63] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_75_0 bl[0] br[0] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_1 bl[1] br[1] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_2 bl[2] br[2] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_3 bl[3] br[3] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_4 bl[4] br[4] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_5 bl[5] br[5] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_6 bl[6] br[6] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_7 bl[7] br[7] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_8 bl[8] br[8] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_9 bl[9] br[9] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_10 bl[10] br[10] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_11 bl[11] br[11] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_12 bl[12] br[12] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_13 bl[13] br[13] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_14 bl[14] br[14] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_15 bl[15] br[15] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_16 bl[16] br[16] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_17 bl[17] br[17] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_18 bl[18] br[18] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_19 bl[19] br[19] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_20 bl[20] br[20] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_21 bl[21] br[21] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_22 bl[22] br[22] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_23 bl[23] br[23] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_24 bl[24] br[24] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_25 bl[25] br[25] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_26 bl[26] br[26] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_27 bl[27] br[27] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_28 bl[28] br[28] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_29 bl[29] br[29] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_30 bl[30] br[30] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_31 bl[31] br[31] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_32 bl[32] br[32] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_33 bl[33] br[33] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_34 bl[34] br[34] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_35 bl[35] br[35] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_36 bl[36] br[36] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_37 bl[37] br[37] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_38 bl[38] br[38] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_39 bl[39] br[39] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_40 bl[40] br[40] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_41 bl[41] br[41] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_42 bl[42] br[42] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_43 bl[43] br[43] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_44 bl[44] br[44] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_45 bl[45] br[45] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_46 bl[46] br[46] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_47 bl[47] br[47] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_48 bl[48] br[48] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_49 bl[49] br[49] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_50 bl[50] br[50] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_51 bl[51] br[51] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_52 bl[52] br[52] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_53 bl[53] br[53] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_54 bl[54] br[54] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_55 bl[55] br[55] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_56 bl[56] br[56] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_57 bl[57] br[57] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_58 bl[58] br[58] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_59 bl[59] br[59] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_60 bl[60] br[60] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_61 bl[61] br[61] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_62 bl[62] br[62] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_63 bl[63] br[63] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_76_0 bl[0] br[0] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_1 bl[1] br[1] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_2 bl[2] br[2] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_3 bl[3] br[3] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_4 bl[4] br[4] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_5 bl[5] br[5] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_6 bl[6] br[6] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_7 bl[7] br[7] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_8 bl[8] br[8] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_9 bl[9] br[9] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_10 bl[10] br[10] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_11 bl[11] br[11] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_12 bl[12] br[12] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_13 bl[13] br[13] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_14 bl[14] br[14] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_15 bl[15] br[15] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_16 bl[16] br[16] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_17 bl[17] br[17] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_18 bl[18] br[18] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_19 bl[19] br[19] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_20 bl[20] br[20] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_21 bl[21] br[21] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_22 bl[22] br[22] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_23 bl[23] br[23] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_24 bl[24] br[24] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_25 bl[25] br[25] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_26 bl[26] br[26] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_27 bl[27] br[27] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_28 bl[28] br[28] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_29 bl[29] br[29] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_30 bl[30] br[30] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_31 bl[31] br[31] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_32 bl[32] br[32] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_33 bl[33] br[33] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_34 bl[34] br[34] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_35 bl[35] br[35] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_36 bl[36] br[36] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_37 bl[37] br[37] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_38 bl[38] br[38] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_39 bl[39] br[39] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_40 bl[40] br[40] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_41 bl[41] br[41] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_42 bl[42] br[42] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_43 bl[43] br[43] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_44 bl[44] br[44] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_45 bl[45] br[45] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_46 bl[46] br[46] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_47 bl[47] br[47] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_48 bl[48] br[48] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_49 bl[49] br[49] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_50 bl[50] br[50] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_51 bl[51] br[51] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_52 bl[52] br[52] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_53 bl[53] br[53] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_54 bl[54] br[54] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_55 bl[55] br[55] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_56 bl[56] br[56] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_57 bl[57] br[57] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_58 bl[58] br[58] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_59 bl[59] br[59] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_60 bl[60] br[60] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_61 bl[61] br[61] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_62 bl[62] br[62] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_63 bl[63] br[63] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_77_0 bl[0] br[0] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_1 bl[1] br[1] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_2 bl[2] br[2] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_3 bl[3] br[3] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_4 bl[4] br[4] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_5 bl[5] br[5] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_6 bl[6] br[6] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_7 bl[7] br[7] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_8 bl[8] br[8] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_9 bl[9] br[9] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_10 bl[10] br[10] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_11 bl[11] br[11] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_12 bl[12] br[12] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_13 bl[13] br[13] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_14 bl[14] br[14] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_15 bl[15] br[15] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_16 bl[16] br[16] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_17 bl[17] br[17] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_18 bl[18] br[18] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_19 bl[19] br[19] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_20 bl[20] br[20] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_21 bl[21] br[21] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_22 bl[22] br[22] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_23 bl[23] br[23] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_24 bl[24] br[24] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_25 bl[25] br[25] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_26 bl[26] br[26] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_27 bl[27] br[27] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_28 bl[28] br[28] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_29 bl[29] br[29] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_30 bl[30] br[30] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_31 bl[31] br[31] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_32 bl[32] br[32] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_33 bl[33] br[33] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_34 bl[34] br[34] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_35 bl[35] br[35] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_36 bl[36] br[36] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_37 bl[37] br[37] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_38 bl[38] br[38] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_39 bl[39] br[39] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_40 bl[40] br[40] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_41 bl[41] br[41] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_42 bl[42] br[42] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_43 bl[43] br[43] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_44 bl[44] br[44] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_45 bl[45] br[45] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_46 bl[46] br[46] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_47 bl[47] br[47] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_48 bl[48] br[48] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_49 bl[49] br[49] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_50 bl[50] br[50] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_51 bl[51] br[51] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_52 bl[52] br[52] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_53 bl[53] br[53] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_54 bl[54] br[54] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_55 bl[55] br[55] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_56 bl[56] br[56] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_57 bl[57] br[57] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_58 bl[58] br[58] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_59 bl[59] br[59] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_60 bl[60] br[60] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_61 bl[61] br[61] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_62 bl[62] br[62] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_63 bl[63] br[63] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_78_0 bl[0] br[0] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_1 bl[1] br[1] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_2 bl[2] br[2] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_3 bl[3] br[3] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_4 bl[4] br[4] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_5 bl[5] br[5] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_6 bl[6] br[6] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_7 bl[7] br[7] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_8 bl[8] br[8] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_9 bl[9] br[9] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_10 bl[10] br[10] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_11 bl[11] br[11] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_12 bl[12] br[12] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_13 bl[13] br[13] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_14 bl[14] br[14] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_15 bl[15] br[15] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_16 bl[16] br[16] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_17 bl[17] br[17] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_18 bl[18] br[18] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_19 bl[19] br[19] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_20 bl[20] br[20] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_21 bl[21] br[21] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_22 bl[22] br[22] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_23 bl[23] br[23] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_24 bl[24] br[24] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_25 bl[25] br[25] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_26 bl[26] br[26] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_27 bl[27] br[27] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_28 bl[28] br[28] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_29 bl[29] br[29] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_30 bl[30] br[30] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_31 bl[31] br[31] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_32 bl[32] br[32] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_33 bl[33] br[33] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_34 bl[34] br[34] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_35 bl[35] br[35] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_36 bl[36] br[36] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_37 bl[37] br[37] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_38 bl[38] br[38] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_39 bl[39] br[39] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_40 bl[40] br[40] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_41 bl[41] br[41] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_42 bl[42] br[42] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_43 bl[43] br[43] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_44 bl[44] br[44] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_45 bl[45] br[45] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_46 bl[46] br[46] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_47 bl[47] br[47] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_48 bl[48] br[48] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_49 bl[49] br[49] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_50 bl[50] br[50] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_51 bl[51] br[51] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_52 bl[52] br[52] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_53 bl[53] br[53] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_54 bl[54] br[54] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_55 bl[55] br[55] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_56 bl[56] br[56] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_57 bl[57] br[57] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_58 bl[58] br[58] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_59 bl[59] br[59] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_60 bl[60] br[60] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_61 bl[61] br[61] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_62 bl[62] br[62] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_63 bl[63] br[63] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_79_0 bl[0] br[0] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_1 bl[1] br[1] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_2 bl[2] br[2] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_3 bl[3] br[3] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_4 bl[4] br[4] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_5 bl[5] br[5] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_6 bl[6] br[6] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_7 bl[7] br[7] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_8 bl[8] br[8] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_9 bl[9] br[9] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_10 bl[10] br[10] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_11 bl[11] br[11] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_12 bl[12] br[12] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_13 bl[13] br[13] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_14 bl[14] br[14] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_15 bl[15] br[15] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_16 bl[16] br[16] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_17 bl[17] br[17] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_18 bl[18] br[18] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_19 bl[19] br[19] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_20 bl[20] br[20] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_21 bl[21] br[21] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_22 bl[22] br[22] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_23 bl[23] br[23] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_24 bl[24] br[24] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_25 bl[25] br[25] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_26 bl[26] br[26] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_27 bl[27] br[27] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_28 bl[28] br[28] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_29 bl[29] br[29] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_30 bl[30] br[30] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_31 bl[31] br[31] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_32 bl[32] br[32] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_33 bl[33] br[33] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_34 bl[34] br[34] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_35 bl[35] br[35] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_36 bl[36] br[36] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_37 bl[37] br[37] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_38 bl[38] br[38] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_39 bl[39] br[39] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_40 bl[40] br[40] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_41 bl[41] br[41] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_42 bl[42] br[42] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_43 bl[43] br[43] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_44 bl[44] br[44] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_45 bl[45] br[45] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_46 bl[46] br[46] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_47 bl[47] br[47] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_48 bl[48] br[48] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_49 bl[49] br[49] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_50 bl[50] br[50] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_51 bl[51] br[51] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_52 bl[52] br[52] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_53 bl[53] br[53] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_54 bl[54] br[54] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_55 bl[55] br[55] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_56 bl[56] br[56] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_57 bl[57] br[57] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_58 bl[58] br[58] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_59 bl[59] br[59] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_60 bl[60] br[60] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_61 bl[61] br[61] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_62 bl[62] br[62] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_63 bl[63] br[63] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_80_0 bl[0] br[0] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_1 bl[1] br[1] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_2 bl[2] br[2] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_3 bl[3] br[3] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_4 bl[4] br[4] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_5 bl[5] br[5] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_6 bl[6] br[6] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_7 bl[7] br[7] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_8 bl[8] br[8] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_9 bl[9] br[9] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_10 bl[10] br[10] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_11 bl[11] br[11] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_12 bl[12] br[12] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_13 bl[13] br[13] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_14 bl[14] br[14] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_15 bl[15] br[15] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_16 bl[16] br[16] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_17 bl[17] br[17] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_18 bl[18] br[18] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_19 bl[19] br[19] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_20 bl[20] br[20] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_21 bl[21] br[21] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_22 bl[22] br[22] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_23 bl[23] br[23] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_24 bl[24] br[24] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_25 bl[25] br[25] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_26 bl[26] br[26] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_27 bl[27] br[27] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_28 bl[28] br[28] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_29 bl[29] br[29] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_30 bl[30] br[30] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_31 bl[31] br[31] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_32 bl[32] br[32] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_33 bl[33] br[33] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_34 bl[34] br[34] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_35 bl[35] br[35] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_36 bl[36] br[36] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_37 bl[37] br[37] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_38 bl[38] br[38] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_39 bl[39] br[39] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_40 bl[40] br[40] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_41 bl[41] br[41] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_42 bl[42] br[42] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_43 bl[43] br[43] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_44 bl[44] br[44] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_45 bl[45] br[45] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_46 bl[46] br[46] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_47 bl[47] br[47] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_48 bl[48] br[48] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_49 bl[49] br[49] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_50 bl[50] br[50] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_51 bl[51] br[51] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_52 bl[52] br[52] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_53 bl[53] br[53] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_54 bl[54] br[54] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_55 bl[55] br[55] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_56 bl[56] br[56] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_57 bl[57] br[57] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_58 bl[58] br[58] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_59 bl[59] br[59] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_60 bl[60] br[60] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_61 bl[61] br[61] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_62 bl[62] br[62] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_63 bl[63] br[63] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_81_0 bl[0] br[0] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_1 bl[1] br[1] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_2 bl[2] br[2] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_3 bl[3] br[3] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_4 bl[4] br[4] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_5 bl[5] br[5] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_6 bl[6] br[6] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_7 bl[7] br[7] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_8 bl[8] br[8] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_9 bl[9] br[9] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_10 bl[10] br[10] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_11 bl[11] br[11] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_12 bl[12] br[12] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_13 bl[13] br[13] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_14 bl[14] br[14] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_15 bl[15] br[15] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_16 bl[16] br[16] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_17 bl[17] br[17] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_18 bl[18] br[18] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_19 bl[19] br[19] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_20 bl[20] br[20] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_21 bl[21] br[21] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_22 bl[22] br[22] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_23 bl[23] br[23] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_24 bl[24] br[24] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_25 bl[25] br[25] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_26 bl[26] br[26] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_27 bl[27] br[27] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_28 bl[28] br[28] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_29 bl[29] br[29] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_30 bl[30] br[30] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_31 bl[31] br[31] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_32 bl[32] br[32] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_33 bl[33] br[33] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_34 bl[34] br[34] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_35 bl[35] br[35] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_36 bl[36] br[36] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_37 bl[37] br[37] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_38 bl[38] br[38] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_39 bl[39] br[39] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_40 bl[40] br[40] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_41 bl[41] br[41] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_42 bl[42] br[42] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_43 bl[43] br[43] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_44 bl[44] br[44] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_45 bl[45] br[45] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_46 bl[46] br[46] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_47 bl[47] br[47] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_48 bl[48] br[48] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_49 bl[49] br[49] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_50 bl[50] br[50] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_51 bl[51] br[51] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_52 bl[52] br[52] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_53 bl[53] br[53] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_54 bl[54] br[54] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_55 bl[55] br[55] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_56 bl[56] br[56] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_57 bl[57] br[57] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_58 bl[58] br[58] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_59 bl[59] br[59] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_60 bl[60] br[60] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_61 bl[61] br[61] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_62 bl[62] br[62] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_63 bl[63] br[63] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_82_0 bl[0] br[0] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_1 bl[1] br[1] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_2 bl[2] br[2] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_3 bl[3] br[3] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_4 bl[4] br[4] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_5 bl[5] br[5] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_6 bl[6] br[6] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_7 bl[7] br[7] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_8 bl[8] br[8] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_9 bl[9] br[9] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_10 bl[10] br[10] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_11 bl[11] br[11] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_12 bl[12] br[12] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_13 bl[13] br[13] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_14 bl[14] br[14] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_15 bl[15] br[15] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_16 bl[16] br[16] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_17 bl[17] br[17] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_18 bl[18] br[18] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_19 bl[19] br[19] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_20 bl[20] br[20] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_21 bl[21] br[21] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_22 bl[22] br[22] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_23 bl[23] br[23] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_24 bl[24] br[24] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_25 bl[25] br[25] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_26 bl[26] br[26] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_27 bl[27] br[27] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_28 bl[28] br[28] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_29 bl[29] br[29] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_30 bl[30] br[30] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_31 bl[31] br[31] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_32 bl[32] br[32] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_33 bl[33] br[33] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_34 bl[34] br[34] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_35 bl[35] br[35] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_36 bl[36] br[36] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_37 bl[37] br[37] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_38 bl[38] br[38] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_39 bl[39] br[39] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_40 bl[40] br[40] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_41 bl[41] br[41] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_42 bl[42] br[42] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_43 bl[43] br[43] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_44 bl[44] br[44] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_45 bl[45] br[45] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_46 bl[46] br[46] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_47 bl[47] br[47] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_48 bl[48] br[48] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_49 bl[49] br[49] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_50 bl[50] br[50] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_51 bl[51] br[51] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_52 bl[52] br[52] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_53 bl[53] br[53] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_54 bl[54] br[54] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_55 bl[55] br[55] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_56 bl[56] br[56] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_57 bl[57] br[57] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_58 bl[58] br[58] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_59 bl[59] br[59] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_60 bl[60] br[60] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_61 bl[61] br[61] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_62 bl[62] br[62] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_63 bl[63] br[63] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_83_0 bl[0] br[0] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_1 bl[1] br[1] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_2 bl[2] br[2] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_3 bl[3] br[3] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_4 bl[4] br[4] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_5 bl[5] br[5] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_6 bl[6] br[6] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_7 bl[7] br[7] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_8 bl[8] br[8] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_9 bl[9] br[9] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_10 bl[10] br[10] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_11 bl[11] br[11] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_12 bl[12] br[12] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_13 bl[13] br[13] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_14 bl[14] br[14] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_15 bl[15] br[15] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_16 bl[16] br[16] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_17 bl[17] br[17] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_18 bl[18] br[18] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_19 bl[19] br[19] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_20 bl[20] br[20] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_21 bl[21] br[21] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_22 bl[22] br[22] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_23 bl[23] br[23] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_24 bl[24] br[24] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_25 bl[25] br[25] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_26 bl[26] br[26] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_27 bl[27] br[27] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_28 bl[28] br[28] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_29 bl[29] br[29] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_30 bl[30] br[30] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_31 bl[31] br[31] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_32 bl[32] br[32] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_33 bl[33] br[33] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_34 bl[34] br[34] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_35 bl[35] br[35] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_36 bl[36] br[36] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_37 bl[37] br[37] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_38 bl[38] br[38] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_39 bl[39] br[39] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_40 bl[40] br[40] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_41 bl[41] br[41] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_42 bl[42] br[42] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_43 bl[43] br[43] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_44 bl[44] br[44] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_45 bl[45] br[45] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_46 bl[46] br[46] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_47 bl[47] br[47] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_48 bl[48] br[48] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_49 bl[49] br[49] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_50 bl[50] br[50] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_51 bl[51] br[51] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_52 bl[52] br[52] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_53 bl[53] br[53] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_54 bl[54] br[54] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_55 bl[55] br[55] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_56 bl[56] br[56] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_57 bl[57] br[57] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_58 bl[58] br[58] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_59 bl[59] br[59] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_60 bl[60] br[60] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_61 bl[61] br[61] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_62 bl[62] br[62] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_63 bl[63] br[63] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_84_0 bl[0] br[0] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_1 bl[1] br[1] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_2 bl[2] br[2] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_3 bl[3] br[3] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_4 bl[4] br[4] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_5 bl[5] br[5] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_6 bl[6] br[6] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_7 bl[7] br[7] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_8 bl[8] br[8] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_9 bl[9] br[9] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_10 bl[10] br[10] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_11 bl[11] br[11] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_12 bl[12] br[12] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_13 bl[13] br[13] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_14 bl[14] br[14] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_15 bl[15] br[15] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_16 bl[16] br[16] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_17 bl[17] br[17] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_18 bl[18] br[18] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_19 bl[19] br[19] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_20 bl[20] br[20] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_21 bl[21] br[21] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_22 bl[22] br[22] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_23 bl[23] br[23] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_24 bl[24] br[24] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_25 bl[25] br[25] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_26 bl[26] br[26] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_27 bl[27] br[27] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_28 bl[28] br[28] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_29 bl[29] br[29] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_30 bl[30] br[30] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_31 bl[31] br[31] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_32 bl[32] br[32] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_33 bl[33] br[33] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_34 bl[34] br[34] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_35 bl[35] br[35] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_36 bl[36] br[36] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_37 bl[37] br[37] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_38 bl[38] br[38] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_39 bl[39] br[39] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_40 bl[40] br[40] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_41 bl[41] br[41] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_42 bl[42] br[42] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_43 bl[43] br[43] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_44 bl[44] br[44] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_45 bl[45] br[45] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_46 bl[46] br[46] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_47 bl[47] br[47] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_48 bl[48] br[48] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_49 bl[49] br[49] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_50 bl[50] br[50] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_51 bl[51] br[51] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_52 bl[52] br[52] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_53 bl[53] br[53] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_54 bl[54] br[54] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_55 bl[55] br[55] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_56 bl[56] br[56] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_57 bl[57] br[57] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_58 bl[58] br[58] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_59 bl[59] br[59] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_60 bl[60] br[60] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_61 bl[61] br[61] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_62 bl[62] br[62] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_63 bl[63] br[63] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_85_0 bl[0] br[0] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_1 bl[1] br[1] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_2 bl[2] br[2] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_3 bl[3] br[3] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_4 bl[4] br[4] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_5 bl[5] br[5] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_6 bl[6] br[6] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_7 bl[7] br[7] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_8 bl[8] br[8] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_9 bl[9] br[9] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_10 bl[10] br[10] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_11 bl[11] br[11] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_12 bl[12] br[12] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_13 bl[13] br[13] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_14 bl[14] br[14] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_15 bl[15] br[15] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_16 bl[16] br[16] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_17 bl[17] br[17] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_18 bl[18] br[18] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_19 bl[19] br[19] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_20 bl[20] br[20] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_21 bl[21] br[21] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_22 bl[22] br[22] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_23 bl[23] br[23] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_24 bl[24] br[24] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_25 bl[25] br[25] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_26 bl[26] br[26] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_27 bl[27] br[27] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_28 bl[28] br[28] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_29 bl[29] br[29] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_30 bl[30] br[30] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_31 bl[31] br[31] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_32 bl[32] br[32] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_33 bl[33] br[33] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_34 bl[34] br[34] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_35 bl[35] br[35] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_36 bl[36] br[36] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_37 bl[37] br[37] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_38 bl[38] br[38] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_39 bl[39] br[39] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_40 bl[40] br[40] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_41 bl[41] br[41] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_42 bl[42] br[42] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_43 bl[43] br[43] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_44 bl[44] br[44] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_45 bl[45] br[45] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_46 bl[46] br[46] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_47 bl[47] br[47] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_48 bl[48] br[48] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_49 bl[49] br[49] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_50 bl[50] br[50] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_51 bl[51] br[51] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_52 bl[52] br[52] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_53 bl[53] br[53] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_54 bl[54] br[54] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_55 bl[55] br[55] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_56 bl[56] br[56] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_57 bl[57] br[57] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_58 bl[58] br[58] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_59 bl[59] br[59] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_60 bl[60] br[60] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_61 bl[61] br[61] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_62 bl[62] br[62] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_63 bl[63] br[63] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_86_0 bl[0] br[0] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_1 bl[1] br[1] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_2 bl[2] br[2] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_3 bl[3] br[3] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_4 bl[4] br[4] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_5 bl[5] br[5] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_6 bl[6] br[6] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_7 bl[7] br[7] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_8 bl[8] br[8] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_9 bl[9] br[9] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_10 bl[10] br[10] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_11 bl[11] br[11] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_12 bl[12] br[12] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_13 bl[13] br[13] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_14 bl[14] br[14] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_15 bl[15] br[15] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_16 bl[16] br[16] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_17 bl[17] br[17] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_18 bl[18] br[18] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_19 bl[19] br[19] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_20 bl[20] br[20] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_21 bl[21] br[21] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_22 bl[22] br[22] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_23 bl[23] br[23] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_24 bl[24] br[24] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_25 bl[25] br[25] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_26 bl[26] br[26] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_27 bl[27] br[27] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_28 bl[28] br[28] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_29 bl[29] br[29] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_30 bl[30] br[30] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_31 bl[31] br[31] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_32 bl[32] br[32] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_33 bl[33] br[33] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_34 bl[34] br[34] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_35 bl[35] br[35] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_36 bl[36] br[36] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_37 bl[37] br[37] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_38 bl[38] br[38] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_39 bl[39] br[39] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_40 bl[40] br[40] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_41 bl[41] br[41] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_42 bl[42] br[42] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_43 bl[43] br[43] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_44 bl[44] br[44] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_45 bl[45] br[45] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_46 bl[46] br[46] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_47 bl[47] br[47] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_48 bl[48] br[48] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_49 bl[49] br[49] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_50 bl[50] br[50] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_51 bl[51] br[51] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_52 bl[52] br[52] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_53 bl[53] br[53] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_54 bl[54] br[54] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_55 bl[55] br[55] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_56 bl[56] br[56] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_57 bl[57] br[57] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_58 bl[58] br[58] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_59 bl[59] br[59] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_60 bl[60] br[60] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_61 bl[61] br[61] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_62 bl[62] br[62] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_63 bl[63] br[63] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_87_0 bl[0] br[0] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_1 bl[1] br[1] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_2 bl[2] br[2] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_3 bl[3] br[3] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_4 bl[4] br[4] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_5 bl[5] br[5] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_6 bl[6] br[6] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_7 bl[7] br[7] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_8 bl[8] br[8] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_9 bl[9] br[9] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_10 bl[10] br[10] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_11 bl[11] br[11] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_12 bl[12] br[12] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_13 bl[13] br[13] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_14 bl[14] br[14] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_15 bl[15] br[15] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_16 bl[16] br[16] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_17 bl[17] br[17] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_18 bl[18] br[18] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_19 bl[19] br[19] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_20 bl[20] br[20] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_21 bl[21] br[21] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_22 bl[22] br[22] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_23 bl[23] br[23] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_24 bl[24] br[24] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_25 bl[25] br[25] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_26 bl[26] br[26] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_27 bl[27] br[27] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_28 bl[28] br[28] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_29 bl[29] br[29] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_30 bl[30] br[30] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_31 bl[31] br[31] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_32 bl[32] br[32] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_33 bl[33] br[33] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_34 bl[34] br[34] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_35 bl[35] br[35] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_36 bl[36] br[36] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_37 bl[37] br[37] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_38 bl[38] br[38] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_39 bl[39] br[39] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_40 bl[40] br[40] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_41 bl[41] br[41] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_42 bl[42] br[42] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_43 bl[43] br[43] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_44 bl[44] br[44] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_45 bl[45] br[45] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_46 bl[46] br[46] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_47 bl[47] br[47] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_48 bl[48] br[48] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_49 bl[49] br[49] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_50 bl[50] br[50] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_51 bl[51] br[51] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_52 bl[52] br[52] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_53 bl[53] br[53] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_54 bl[54] br[54] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_55 bl[55] br[55] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_56 bl[56] br[56] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_57 bl[57] br[57] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_58 bl[58] br[58] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_59 bl[59] br[59] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_60 bl[60] br[60] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_61 bl[61] br[61] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_62 bl[62] br[62] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_63 bl[63] br[63] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_88_0 bl[0] br[0] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_1 bl[1] br[1] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_2 bl[2] br[2] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_3 bl[3] br[3] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_4 bl[4] br[4] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_5 bl[5] br[5] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_6 bl[6] br[6] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_7 bl[7] br[7] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_8 bl[8] br[8] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_9 bl[9] br[9] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_10 bl[10] br[10] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_11 bl[11] br[11] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_12 bl[12] br[12] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_13 bl[13] br[13] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_14 bl[14] br[14] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_15 bl[15] br[15] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_16 bl[16] br[16] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_17 bl[17] br[17] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_18 bl[18] br[18] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_19 bl[19] br[19] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_20 bl[20] br[20] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_21 bl[21] br[21] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_22 bl[22] br[22] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_23 bl[23] br[23] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_24 bl[24] br[24] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_25 bl[25] br[25] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_26 bl[26] br[26] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_27 bl[27] br[27] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_28 bl[28] br[28] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_29 bl[29] br[29] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_30 bl[30] br[30] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_31 bl[31] br[31] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_32 bl[32] br[32] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_33 bl[33] br[33] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_34 bl[34] br[34] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_35 bl[35] br[35] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_36 bl[36] br[36] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_37 bl[37] br[37] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_38 bl[38] br[38] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_39 bl[39] br[39] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_40 bl[40] br[40] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_41 bl[41] br[41] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_42 bl[42] br[42] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_43 bl[43] br[43] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_44 bl[44] br[44] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_45 bl[45] br[45] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_46 bl[46] br[46] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_47 bl[47] br[47] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_48 bl[48] br[48] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_49 bl[49] br[49] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_50 bl[50] br[50] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_51 bl[51] br[51] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_52 bl[52] br[52] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_53 bl[53] br[53] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_54 bl[54] br[54] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_55 bl[55] br[55] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_56 bl[56] br[56] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_57 bl[57] br[57] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_58 bl[58] br[58] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_59 bl[59] br[59] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_60 bl[60] br[60] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_61 bl[61] br[61] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_62 bl[62] br[62] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_63 bl[63] br[63] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_89_0 bl[0] br[0] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_1 bl[1] br[1] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_2 bl[2] br[2] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_3 bl[3] br[3] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_4 bl[4] br[4] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_5 bl[5] br[5] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_6 bl[6] br[6] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_7 bl[7] br[7] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_8 bl[8] br[8] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_9 bl[9] br[9] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_10 bl[10] br[10] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_11 bl[11] br[11] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_12 bl[12] br[12] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_13 bl[13] br[13] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_14 bl[14] br[14] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_15 bl[15] br[15] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_16 bl[16] br[16] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_17 bl[17] br[17] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_18 bl[18] br[18] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_19 bl[19] br[19] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_20 bl[20] br[20] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_21 bl[21] br[21] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_22 bl[22] br[22] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_23 bl[23] br[23] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_24 bl[24] br[24] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_25 bl[25] br[25] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_26 bl[26] br[26] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_27 bl[27] br[27] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_28 bl[28] br[28] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_29 bl[29] br[29] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_30 bl[30] br[30] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_31 bl[31] br[31] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_32 bl[32] br[32] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_33 bl[33] br[33] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_34 bl[34] br[34] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_35 bl[35] br[35] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_36 bl[36] br[36] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_37 bl[37] br[37] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_38 bl[38] br[38] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_39 bl[39] br[39] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_40 bl[40] br[40] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_41 bl[41] br[41] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_42 bl[42] br[42] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_43 bl[43] br[43] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_44 bl[44] br[44] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_45 bl[45] br[45] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_46 bl[46] br[46] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_47 bl[47] br[47] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_48 bl[48] br[48] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_49 bl[49] br[49] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_50 bl[50] br[50] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_51 bl[51] br[51] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_52 bl[52] br[52] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_53 bl[53] br[53] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_54 bl[54] br[54] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_55 bl[55] br[55] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_56 bl[56] br[56] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_57 bl[57] br[57] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_58 bl[58] br[58] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_59 bl[59] br[59] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_60 bl[60] br[60] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_61 bl[61] br[61] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_62 bl[62] br[62] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_63 bl[63] br[63] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_90_0 bl[0] br[0] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_1 bl[1] br[1] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_2 bl[2] br[2] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_3 bl[3] br[3] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_4 bl[4] br[4] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_5 bl[5] br[5] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_6 bl[6] br[6] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_7 bl[7] br[7] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_8 bl[8] br[8] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_9 bl[9] br[9] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_10 bl[10] br[10] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_11 bl[11] br[11] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_12 bl[12] br[12] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_13 bl[13] br[13] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_14 bl[14] br[14] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_15 bl[15] br[15] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_16 bl[16] br[16] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_17 bl[17] br[17] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_18 bl[18] br[18] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_19 bl[19] br[19] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_20 bl[20] br[20] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_21 bl[21] br[21] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_22 bl[22] br[22] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_23 bl[23] br[23] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_24 bl[24] br[24] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_25 bl[25] br[25] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_26 bl[26] br[26] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_27 bl[27] br[27] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_28 bl[28] br[28] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_29 bl[29] br[29] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_30 bl[30] br[30] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_31 bl[31] br[31] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_32 bl[32] br[32] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_33 bl[33] br[33] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_34 bl[34] br[34] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_35 bl[35] br[35] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_36 bl[36] br[36] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_37 bl[37] br[37] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_38 bl[38] br[38] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_39 bl[39] br[39] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_40 bl[40] br[40] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_41 bl[41] br[41] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_42 bl[42] br[42] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_43 bl[43] br[43] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_44 bl[44] br[44] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_45 bl[45] br[45] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_46 bl[46] br[46] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_47 bl[47] br[47] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_48 bl[48] br[48] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_49 bl[49] br[49] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_50 bl[50] br[50] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_51 bl[51] br[51] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_52 bl[52] br[52] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_53 bl[53] br[53] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_54 bl[54] br[54] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_55 bl[55] br[55] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_56 bl[56] br[56] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_57 bl[57] br[57] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_58 bl[58] br[58] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_59 bl[59] br[59] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_60 bl[60] br[60] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_61 bl[61] br[61] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_62 bl[62] br[62] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_63 bl[63] br[63] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_91_0 bl[0] br[0] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_1 bl[1] br[1] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_2 bl[2] br[2] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_3 bl[3] br[3] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_4 bl[4] br[4] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_5 bl[5] br[5] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_6 bl[6] br[6] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_7 bl[7] br[7] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_8 bl[8] br[8] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_9 bl[9] br[9] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_10 bl[10] br[10] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_11 bl[11] br[11] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_12 bl[12] br[12] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_13 bl[13] br[13] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_14 bl[14] br[14] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_15 bl[15] br[15] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_16 bl[16] br[16] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_17 bl[17] br[17] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_18 bl[18] br[18] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_19 bl[19] br[19] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_20 bl[20] br[20] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_21 bl[21] br[21] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_22 bl[22] br[22] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_23 bl[23] br[23] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_24 bl[24] br[24] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_25 bl[25] br[25] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_26 bl[26] br[26] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_27 bl[27] br[27] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_28 bl[28] br[28] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_29 bl[29] br[29] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_30 bl[30] br[30] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_31 bl[31] br[31] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_32 bl[32] br[32] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_33 bl[33] br[33] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_34 bl[34] br[34] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_35 bl[35] br[35] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_36 bl[36] br[36] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_37 bl[37] br[37] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_38 bl[38] br[38] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_39 bl[39] br[39] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_40 bl[40] br[40] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_41 bl[41] br[41] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_42 bl[42] br[42] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_43 bl[43] br[43] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_44 bl[44] br[44] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_45 bl[45] br[45] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_46 bl[46] br[46] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_47 bl[47] br[47] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_48 bl[48] br[48] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_49 bl[49] br[49] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_50 bl[50] br[50] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_51 bl[51] br[51] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_52 bl[52] br[52] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_53 bl[53] br[53] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_54 bl[54] br[54] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_55 bl[55] br[55] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_56 bl[56] br[56] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_57 bl[57] br[57] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_58 bl[58] br[58] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_59 bl[59] br[59] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_60 bl[60] br[60] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_61 bl[61] br[61] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_62 bl[62] br[62] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_63 bl[63] br[63] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_92_0 bl[0] br[0] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_1 bl[1] br[1] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_2 bl[2] br[2] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_3 bl[3] br[3] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_4 bl[4] br[4] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_5 bl[5] br[5] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_6 bl[6] br[6] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_7 bl[7] br[7] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_8 bl[8] br[8] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_9 bl[9] br[9] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_10 bl[10] br[10] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_11 bl[11] br[11] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_12 bl[12] br[12] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_13 bl[13] br[13] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_14 bl[14] br[14] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_15 bl[15] br[15] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_16 bl[16] br[16] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_17 bl[17] br[17] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_18 bl[18] br[18] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_19 bl[19] br[19] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_20 bl[20] br[20] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_21 bl[21] br[21] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_22 bl[22] br[22] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_23 bl[23] br[23] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_24 bl[24] br[24] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_25 bl[25] br[25] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_26 bl[26] br[26] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_27 bl[27] br[27] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_28 bl[28] br[28] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_29 bl[29] br[29] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_30 bl[30] br[30] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_31 bl[31] br[31] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_32 bl[32] br[32] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_33 bl[33] br[33] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_34 bl[34] br[34] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_35 bl[35] br[35] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_36 bl[36] br[36] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_37 bl[37] br[37] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_38 bl[38] br[38] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_39 bl[39] br[39] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_40 bl[40] br[40] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_41 bl[41] br[41] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_42 bl[42] br[42] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_43 bl[43] br[43] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_44 bl[44] br[44] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_45 bl[45] br[45] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_46 bl[46] br[46] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_47 bl[47] br[47] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_48 bl[48] br[48] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_49 bl[49] br[49] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_50 bl[50] br[50] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_51 bl[51] br[51] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_52 bl[52] br[52] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_53 bl[53] br[53] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_54 bl[54] br[54] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_55 bl[55] br[55] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_56 bl[56] br[56] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_57 bl[57] br[57] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_58 bl[58] br[58] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_59 bl[59] br[59] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_60 bl[60] br[60] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_61 bl[61] br[61] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_62 bl[62] br[62] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_63 bl[63] br[63] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_93_0 bl[0] br[0] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_1 bl[1] br[1] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_2 bl[2] br[2] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_3 bl[3] br[3] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_4 bl[4] br[4] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_5 bl[5] br[5] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_6 bl[6] br[6] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_7 bl[7] br[7] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_8 bl[8] br[8] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_9 bl[9] br[9] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_10 bl[10] br[10] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_11 bl[11] br[11] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_12 bl[12] br[12] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_13 bl[13] br[13] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_14 bl[14] br[14] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_15 bl[15] br[15] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_16 bl[16] br[16] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_17 bl[17] br[17] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_18 bl[18] br[18] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_19 bl[19] br[19] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_20 bl[20] br[20] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_21 bl[21] br[21] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_22 bl[22] br[22] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_23 bl[23] br[23] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_24 bl[24] br[24] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_25 bl[25] br[25] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_26 bl[26] br[26] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_27 bl[27] br[27] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_28 bl[28] br[28] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_29 bl[29] br[29] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_30 bl[30] br[30] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_31 bl[31] br[31] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_32 bl[32] br[32] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_33 bl[33] br[33] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_34 bl[34] br[34] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_35 bl[35] br[35] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_36 bl[36] br[36] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_37 bl[37] br[37] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_38 bl[38] br[38] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_39 bl[39] br[39] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_40 bl[40] br[40] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_41 bl[41] br[41] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_42 bl[42] br[42] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_43 bl[43] br[43] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_44 bl[44] br[44] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_45 bl[45] br[45] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_46 bl[46] br[46] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_47 bl[47] br[47] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_48 bl[48] br[48] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_49 bl[49] br[49] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_50 bl[50] br[50] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_51 bl[51] br[51] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_52 bl[52] br[52] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_53 bl[53] br[53] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_54 bl[54] br[54] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_55 bl[55] br[55] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_56 bl[56] br[56] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_57 bl[57] br[57] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_58 bl[58] br[58] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_59 bl[59] br[59] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_60 bl[60] br[60] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_61 bl[61] br[61] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_62 bl[62] br[62] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_63 bl[63] br[63] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_94_0 bl[0] br[0] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_1 bl[1] br[1] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_2 bl[2] br[2] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_3 bl[3] br[3] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_4 bl[4] br[4] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_5 bl[5] br[5] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_6 bl[6] br[6] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_7 bl[7] br[7] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_8 bl[8] br[8] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_9 bl[9] br[9] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_10 bl[10] br[10] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_11 bl[11] br[11] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_12 bl[12] br[12] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_13 bl[13] br[13] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_14 bl[14] br[14] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_15 bl[15] br[15] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_16 bl[16] br[16] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_17 bl[17] br[17] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_18 bl[18] br[18] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_19 bl[19] br[19] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_20 bl[20] br[20] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_21 bl[21] br[21] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_22 bl[22] br[22] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_23 bl[23] br[23] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_24 bl[24] br[24] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_25 bl[25] br[25] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_26 bl[26] br[26] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_27 bl[27] br[27] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_28 bl[28] br[28] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_29 bl[29] br[29] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_30 bl[30] br[30] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_31 bl[31] br[31] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_32 bl[32] br[32] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_33 bl[33] br[33] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_34 bl[34] br[34] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_35 bl[35] br[35] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_36 bl[36] br[36] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_37 bl[37] br[37] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_38 bl[38] br[38] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_39 bl[39] br[39] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_40 bl[40] br[40] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_41 bl[41] br[41] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_42 bl[42] br[42] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_43 bl[43] br[43] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_44 bl[44] br[44] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_45 bl[45] br[45] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_46 bl[46] br[46] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_47 bl[47] br[47] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_48 bl[48] br[48] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_49 bl[49] br[49] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_50 bl[50] br[50] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_51 bl[51] br[51] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_52 bl[52] br[52] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_53 bl[53] br[53] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_54 bl[54] br[54] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_55 bl[55] br[55] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_56 bl[56] br[56] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_57 bl[57] br[57] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_58 bl[58] br[58] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_59 bl[59] br[59] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_60 bl[60] br[60] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_61 bl[61] br[61] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_62 bl[62] br[62] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_63 bl[63] br[63] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_95_0 bl[0] br[0] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_1 bl[1] br[1] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_2 bl[2] br[2] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_3 bl[3] br[3] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_4 bl[4] br[4] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_5 bl[5] br[5] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_6 bl[6] br[6] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_7 bl[7] br[7] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_8 bl[8] br[8] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_9 bl[9] br[9] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_10 bl[10] br[10] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_11 bl[11] br[11] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_12 bl[12] br[12] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_13 bl[13] br[13] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_14 bl[14] br[14] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_15 bl[15] br[15] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_16 bl[16] br[16] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_17 bl[17] br[17] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_18 bl[18] br[18] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_19 bl[19] br[19] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_20 bl[20] br[20] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_21 bl[21] br[21] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_22 bl[22] br[22] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_23 bl[23] br[23] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_24 bl[24] br[24] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_25 bl[25] br[25] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_26 bl[26] br[26] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_27 bl[27] br[27] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_28 bl[28] br[28] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_29 bl[29] br[29] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_30 bl[30] br[30] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_31 bl[31] br[31] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_32 bl[32] br[32] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_33 bl[33] br[33] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_34 bl[34] br[34] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_35 bl[35] br[35] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_36 bl[36] br[36] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_37 bl[37] br[37] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_38 bl[38] br[38] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_39 bl[39] br[39] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_40 bl[40] br[40] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_41 bl[41] br[41] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_42 bl[42] br[42] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_43 bl[43] br[43] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_44 bl[44] br[44] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_45 bl[45] br[45] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_46 bl[46] br[46] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_47 bl[47] br[47] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_48 bl[48] br[48] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_49 bl[49] br[49] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_50 bl[50] br[50] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_51 bl[51] br[51] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_52 bl[52] br[52] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_53 bl[53] br[53] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_54 bl[54] br[54] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_55 bl[55] br[55] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_56 bl[56] br[56] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_57 bl[57] br[57] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_58 bl[58] br[58] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_59 bl[59] br[59] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_60 bl[60] br[60] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_61 bl[61] br[61] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_62 bl[62] br[62] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_63 bl[63] br[63] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_96_0 bl[0] br[0] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_1 bl[1] br[1] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_2 bl[2] br[2] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_3 bl[3] br[3] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_4 bl[4] br[4] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_5 bl[5] br[5] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_6 bl[6] br[6] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_7 bl[7] br[7] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_8 bl[8] br[8] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_9 bl[9] br[9] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_10 bl[10] br[10] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_11 bl[11] br[11] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_12 bl[12] br[12] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_13 bl[13] br[13] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_14 bl[14] br[14] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_15 bl[15] br[15] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_16 bl[16] br[16] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_17 bl[17] br[17] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_18 bl[18] br[18] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_19 bl[19] br[19] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_20 bl[20] br[20] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_21 bl[21] br[21] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_22 bl[22] br[22] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_23 bl[23] br[23] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_24 bl[24] br[24] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_25 bl[25] br[25] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_26 bl[26] br[26] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_27 bl[27] br[27] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_28 bl[28] br[28] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_29 bl[29] br[29] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_30 bl[30] br[30] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_31 bl[31] br[31] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_32 bl[32] br[32] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_33 bl[33] br[33] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_34 bl[34] br[34] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_35 bl[35] br[35] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_36 bl[36] br[36] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_37 bl[37] br[37] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_38 bl[38] br[38] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_39 bl[39] br[39] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_40 bl[40] br[40] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_41 bl[41] br[41] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_42 bl[42] br[42] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_43 bl[43] br[43] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_44 bl[44] br[44] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_45 bl[45] br[45] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_46 bl[46] br[46] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_47 bl[47] br[47] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_48 bl[48] br[48] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_49 bl[49] br[49] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_50 bl[50] br[50] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_51 bl[51] br[51] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_52 bl[52] br[52] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_53 bl[53] br[53] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_54 bl[54] br[54] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_55 bl[55] br[55] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_56 bl[56] br[56] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_57 bl[57] br[57] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_58 bl[58] br[58] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_59 bl[59] br[59] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_60 bl[60] br[60] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_61 bl[61] br[61] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_62 bl[62] br[62] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_63 bl[63] br[63] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_97_0 bl[0] br[0] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_1 bl[1] br[1] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_2 bl[2] br[2] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_3 bl[3] br[3] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_4 bl[4] br[4] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_5 bl[5] br[5] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_6 bl[6] br[6] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_7 bl[7] br[7] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_8 bl[8] br[8] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_9 bl[9] br[9] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_10 bl[10] br[10] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_11 bl[11] br[11] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_12 bl[12] br[12] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_13 bl[13] br[13] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_14 bl[14] br[14] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_15 bl[15] br[15] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_16 bl[16] br[16] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_17 bl[17] br[17] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_18 bl[18] br[18] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_19 bl[19] br[19] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_20 bl[20] br[20] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_21 bl[21] br[21] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_22 bl[22] br[22] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_23 bl[23] br[23] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_24 bl[24] br[24] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_25 bl[25] br[25] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_26 bl[26] br[26] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_27 bl[27] br[27] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_28 bl[28] br[28] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_29 bl[29] br[29] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_30 bl[30] br[30] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_31 bl[31] br[31] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_32 bl[32] br[32] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_33 bl[33] br[33] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_34 bl[34] br[34] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_35 bl[35] br[35] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_36 bl[36] br[36] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_37 bl[37] br[37] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_38 bl[38] br[38] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_39 bl[39] br[39] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_40 bl[40] br[40] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_41 bl[41] br[41] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_42 bl[42] br[42] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_43 bl[43] br[43] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_44 bl[44] br[44] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_45 bl[45] br[45] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_46 bl[46] br[46] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_47 bl[47] br[47] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_48 bl[48] br[48] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_49 bl[49] br[49] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_50 bl[50] br[50] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_51 bl[51] br[51] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_52 bl[52] br[52] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_53 bl[53] br[53] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_54 bl[54] br[54] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_55 bl[55] br[55] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_56 bl[56] br[56] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_57 bl[57] br[57] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_58 bl[58] br[58] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_59 bl[59] br[59] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_60 bl[60] br[60] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_61 bl[61] br[61] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_62 bl[62] br[62] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_63 bl[63] br[63] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_98_0 bl[0] br[0] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_1 bl[1] br[1] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_2 bl[2] br[2] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_3 bl[3] br[3] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_4 bl[4] br[4] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_5 bl[5] br[5] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_6 bl[6] br[6] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_7 bl[7] br[7] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_8 bl[8] br[8] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_9 bl[9] br[9] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_10 bl[10] br[10] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_11 bl[11] br[11] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_12 bl[12] br[12] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_13 bl[13] br[13] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_14 bl[14] br[14] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_15 bl[15] br[15] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_16 bl[16] br[16] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_17 bl[17] br[17] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_18 bl[18] br[18] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_19 bl[19] br[19] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_20 bl[20] br[20] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_21 bl[21] br[21] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_22 bl[22] br[22] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_23 bl[23] br[23] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_24 bl[24] br[24] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_25 bl[25] br[25] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_26 bl[26] br[26] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_27 bl[27] br[27] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_28 bl[28] br[28] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_29 bl[29] br[29] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_30 bl[30] br[30] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_31 bl[31] br[31] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_32 bl[32] br[32] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_33 bl[33] br[33] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_34 bl[34] br[34] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_35 bl[35] br[35] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_36 bl[36] br[36] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_37 bl[37] br[37] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_38 bl[38] br[38] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_39 bl[39] br[39] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_40 bl[40] br[40] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_41 bl[41] br[41] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_42 bl[42] br[42] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_43 bl[43] br[43] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_44 bl[44] br[44] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_45 bl[45] br[45] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_46 bl[46] br[46] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_47 bl[47] br[47] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_48 bl[48] br[48] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_49 bl[49] br[49] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_50 bl[50] br[50] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_51 bl[51] br[51] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_52 bl[52] br[52] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_53 bl[53] br[53] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_54 bl[54] br[54] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_55 bl[55] br[55] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_56 bl[56] br[56] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_57 bl[57] br[57] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_58 bl[58] br[58] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_59 bl[59] br[59] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_60 bl[60] br[60] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_61 bl[61] br[61] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_62 bl[62] br[62] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_63 bl[63] br[63] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_99_0 bl[0] br[0] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_1 bl[1] br[1] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_2 bl[2] br[2] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_3 bl[3] br[3] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_4 bl[4] br[4] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_5 bl[5] br[5] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_6 bl[6] br[6] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_7 bl[7] br[7] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_8 bl[8] br[8] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_9 bl[9] br[9] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_10 bl[10] br[10] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_11 bl[11] br[11] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_12 bl[12] br[12] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_13 bl[13] br[13] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_14 bl[14] br[14] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_15 bl[15] br[15] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_16 bl[16] br[16] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_17 bl[17] br[17] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_18 bl[18] br[18] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_19 bl[19] br[19] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_20 bl[20] br[20] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_21 bl[21] br[21] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_22 bl[22] br[22] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_23 bl[23] br[23] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_24 bl[24] br[24] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_25 bl[25] br[25] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_26 bl[26] br[26] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_27 bl[27] br[27] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_28 bl[28] br[28] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_29 bl[29] br[29] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_30 bl[30] br[30] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_31 bl[31] br[31] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_32 bl[32] br[32] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_33 bl[33] br[33] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_34 bl[34] br[34] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_35 bl[35] br[35] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_36 bl[36] br[36] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_37 bl[37] br[37] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_38 bl[38] br[38] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_39 bl[39] br[39] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_40 bl[40] br[40] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_41 bl[41] br[41] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_42 bl[42] br[42] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_43 bl[43] br[43] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_44 bl[44] br[44] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_45 bl[45] br[45] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_46 bl[46] br[46] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_47 bl[47] br[47] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_48 bl[48] br[48] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_49 bl[49] br[49] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_50 bl[50] br[50] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_51 bl[51] br[51] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_52 bl[52] br[52] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_53 bl[53] br[53] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_54 bl[54] br[54] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_55 bl[55] br[55] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_56 bl[56] br[56] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_57 bl[57] br[57] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_58 bl[58] br[58] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_59 bl[59] br[59] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_60 bl[60] br[60] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_61 bl[61] br[61] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_62 bl[62] br[62] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_63 bl[63] br[63] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_100_0 bl[0] br[0] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_1 bl[1] br[1] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_2 bl[2] br[2] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_3 bl[3] br[3] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_4 bl[4] br[4] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_5 bl[5] br[5] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_6 bl[6] br[6] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_7 bl[7] br[7] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_8 bl[8] br[8] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_9 bl[9] br[9] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_10 bl[10] br[10] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_11 bl[11] br[11] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_12 bl[12] br[12] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_13 bl[13] br[13] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_14 bl[14] br[14] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_15 bl[15] br[15] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_16 bl[16] br[16] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_17 bl[17] br[17] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_18 bl[18] br[18] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_19 bl[19] br[19] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_20 bl[20] br[20] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_21 bl[21] br[21] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_22 bl[22] br[22] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_23 bl[23] br[23] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_24 bl[24] br[24] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_25 bl[25] br[25] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_26 bl[26] br[26] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_27 bl[27] br[27] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_28 bl[28] br[28] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_29 bl[29] br[29] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_30 bl[30] br[30] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_31 bl[31] br[31] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_32 bl[32] br[32] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_33 bl[33] br[33] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_34 bl[34] br[34] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_35 bl[35] br[35] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_36 bl[36] br[36] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_37 bl[37] br[37] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_38 bl[38] br[38] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_39 bl[39] br[39] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_40 bl[40] br[40] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_41 bl[41] br[41] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_42 bl[42] br[42] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_43 bl[43] br[43] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_44 bl[44] br[44] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_45 bl[45] br[45] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_46 bl[46] br[46] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_47 bl[47] br[47] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_48 bl[48] br[48] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_49 bl[49] br[49] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_50 bl[50] br[50] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_51 bl[51] br[51] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_52 bl[52] br[52] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_53 bl[53] br[53] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_54 bl[54] br[54] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_55 bl[55] br[55] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_56 bl[56] br[56] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_57 bl[57] br[57] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_58 bl[58] br[58] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_59 bl[59] br[59] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_60 bl[60] br[60] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_61 bl[61] br[61] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_62 bl[62] br[62] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_63 bl[63] br[63] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_101_0 bl[0] br[0] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_1 bl[1] br[1] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_2 bl[2] br[2] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_3 bl[3] br[3] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_4 bl[4] br[4] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_5 bl[5] br[5] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_6 bl[6] br[6] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_7 bl[7] br[7] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_8 bl[8] br[8] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_9 bl[9] br[9] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_10 bl[10] br[10] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_11 bl[11] br[11] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_12 bl[12] br[12] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_13 bl[13] br[13] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_14 bl[14] br[14] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_15 bl[15] br[15] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_16 bl[16] br[16] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_17 bl[17] br[17] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_18 bl[18] br[18] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_19 bl[19] br[19] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_20 bl[20] br[20] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_21 bl[21] br[21] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_22 bl[22] br[22] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_23 bl[23] br[23] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_24 bl[24] br[24] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_25 bl[25] br[25] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_26 bl[26] br[26] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_27 bl[27] br[27] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_28 bl[28] br[28] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_29 bl[29] br[29] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_30 bl[30] br[30] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_31 bl[31] br[31] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_32 bl[32] br[32] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_33 bl[33] br[33] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_34 bl[34] br[34] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_35 bl[35] br[35] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_36 bl[36] br[36] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_37 bl[37] br[37] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_38 bl[38] br[38] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_39 bl[39] br[39] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_40 bl[40] br[40] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_41 bl[41] br[41] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_42 bl[42] br[42] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_43 bl[43] br[43] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_44 bl[44] br[44] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_45 bl[45] br[45] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_46 bl[46] br[46] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_47 bl[47] br[47] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_48 bl[48] br[48] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_49 bl[49] br[49] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_50 bl[50] br[50] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_51 bl[51] br[51] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_52 bl[52] br[52] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_53 bl[53] br[53] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_54 bl[54] br[54] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_55 bl[55] br[55] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_56 bl[56] br[56] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_57 bl[57] br[57] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_58 bl[58] br[58] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_59 bl[59] br[59] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_60 bl[60] br[60] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_61 bl[61] br[61] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_62 bl[62] br[62] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_63 bl[63] br[63] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_102_0 bl[0] br[0] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_1 bl[1] br[1] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_2 bl[2] br[2] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_3 bl[3] br[3] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_4 bl[4] br[4] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_5 bl[5] br[5] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_6 bl[6] br[6] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_7 bl[7] br[7] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_8 bl[8] br[8] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_9 bl[9] br[9] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_10 bl[10] br[10] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_11 bl[11] br[11] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_12 bl[12] br[12] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_13 bl[13] br[13] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_14 bl[14] br[14] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_15 bl[15] br[15] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_16 bl[16] br[16] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_17 bl[17] br[17] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_18 bl[18] br[18] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_19 bl[19] br[19] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_20 bl[20] br[20] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_21 bl[21] br[21] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_22 bl[22] br[22] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_23 bl[23] br[23] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_24 bl[24] br[24] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_25 bl[25] br[25] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_26 bl[26] br[26] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_27 bl[27] br[27] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_28 bl[28] br[28] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_29 bl[29] br[29] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_30 bl[30] br[30] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_31 bl[31] br[31] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_32 bl[32] br[32] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_33 bl[33] br[33] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_34 bl[34] br[34] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_35 bl[35] br[35] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_36 bl[36] br[36] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_37 bl[37] br[37] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_38 bl[38] br[38] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_39 bl[39] br[39] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_40 bl[40] br[40] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_41 bl[41] br[41] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_42 bl[42] br[42] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_43 bl[43] br[43] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_44 bl[44] br[44] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_45 bl[45] br[45] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_46 bl[46] br[46] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_47 bl[47] br[47] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_48 bl[48] br[48] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_49 bl[49] br[49] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_50 bl[50] br[50] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_51 bl[51] br[51] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_52 bl[52] br[52] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_53 bl[53] br[53] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_54 bl[54] br[54] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_55 bl[55] br[55] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_56 bl[56] br[56] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_57 bl[57] br[57] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_58 bl[58] br[58] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_59 bl[59] br[59] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_60 bl[60] br[60] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_61 bl[61] br[61] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_62 bl[62] br[62] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_63 bl[63] br[63] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_103_0 bl[0] br[0] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_1 bl[1] br[1] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_2 bl[2] br[2] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_3 bl[3] br[3] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_4 bl[4] br[4] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_5 bl[5] br[5] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_6 bl[6] br[6] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_7 bl[7] br[7] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_8 bl[8] br[8] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_9 bl[9] br[9] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_10 bl[10] br[10] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_11 bl[11] br[11] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_12 bl[12] br[12] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_13 bl[13] br[13] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_14 bl[14] br[14] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_15 bl[15] br[15] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_16 bl[16] br[16] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_17 bl[17] br[17] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_18 bl[18] br[18] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_19 bl[19] br[19] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_20 bl[20] br[20] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_21 bl[21] br[21] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_22 bl[22] br[22] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_23 bl[23] br[23] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_24 bl[24] br[24] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_25 bl[25] br[25] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_26 bl[26] br[26] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_27 bl[27] br[27] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_28 bl[28] br[28] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_29 bl[29] br[29] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_30 bl[30] br[30] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_31 bl[31] br[31] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_32 bl[32] br[32] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_33 bl[33] br[33] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_34 bl[34] br[34] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_35 bl[35] br[35] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_36 bl[36] br[36] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_37 bl[37] br[37] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_38 bl[38] br[38] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_39 bl[39] br[39] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_40 bl[40] br[40] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_41 bl[41] br[41] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_42 bl[42] br[42] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_43 bl[43] br[43] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_44 bl[44] br[44] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_45 bl[45] br[45] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_46 bl[46] br[46] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_47 bl[47] br[47] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_48 bl[48] br[48] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_49 bl[49] br[49] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_50 bl[50] br[50] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_51 bl[51] br[51] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_52 bl[52] br[52] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_53 bl[53] br[53] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_54 bl[54] br[54] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_55 bl[55] br[55] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_56 bl[56] br[56] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_57 bl[57] br[57] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_58 bl[58] br[58] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_59 bl[59] br[59] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_60 bl[60] br[60] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_61 bl[61] br[61] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_62 bl[62] br[62] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_63 bl[63] br[63] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_104_0 bl[0] br[0] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_1 bl[1] br[1] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_2 bl[2] br[2] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_3 bl[3] br[3] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_4 bl[4] br[4] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_5 bl[5] br[5] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_6 bl[6] br[6] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_7 bl[7] br[7] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_8 bl[8] br[8] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_9 bl[9] br[9] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_10 bl[10] br[10] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_11 bl[11] br[11] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_12 bl[12] br[12] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_13 bl[13] br[13] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_14 bl[14] br[14] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_15 bl[15] br[15] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_16 bl[16] br[16] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_17 bl[17] br[17] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_18 bl[18] br[18] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_19 bl[19] br[19] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_20 bl[20] br[20] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_21 bl[21] br[21] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_22 bl[22] br[22] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_23 bl[23] br[23] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_24 bl[24] br[24] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_25 bl[25] br[25] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_26 bl[26] br[26] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_27 bl[27] br[27] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_28 bl[28] br[28] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_29 bl[29] br[29] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_30 bl[30] br[30] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_31 bl[31] br[31] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_32 bl[32] br[32] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_33 bl[33] br[33] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_34 bl[34] br[34] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_35 bl[35] br[35] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_36 bl[36] br[36] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_37 bl[37] br[37] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_38 bl[38] br[38] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_39 bl[39] br[39] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_40 bl[40] br[40] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_41 bl[41] br[41] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_42 bl[42] br[42] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_43 bl[43] br[43] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_44 bl[44] br[44] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_45 bl[45] br[45] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_46 bl[46] br[46] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_47 bl[47] br[47] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_48 bl[48] br[48] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_49 bl[49] br[49] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_50 bl[50] br[50] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_51 bl[51] br[51] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_52 bl[52] br[52] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_53 bl[53] br[53] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_54 bl[54] br[54] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_55 bl[55] br[55] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_56 bl[56] br[56] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_57 bl[57] br[57] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_58 bl[58] br[58] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_59 bl[59] br[59] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_60 bl[60] br[60] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_61 bl[61] br[61] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_62 bl[62] br[62] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_63 bl[63] br[63] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_105_0 bl[0] br[0] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_1 bl[1] br[1] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_2 bl[2] br[2] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_3 bl[3] br[3] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_4 bl[4] br[4] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_5 bl[5] br[5] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_6 bl[6] br[6] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_7 bl[7] br[7] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_8 bl[8] br[8] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_9 bl[9] br[9] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_10 bl[10] br[10] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_11 bl[11] br[11] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_12 bl[12] br[12] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_13 bl[13] br[13] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_14 bl[14] br[14] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_15 bl[15] br[15] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_16 bl[16] br[16] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_17 bl[17] br[17] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_18 bl[18] br[18] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_19 bl[19] br[19] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_20 bl[20] br[20] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_21 bl[21] br[21] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_22 bl[22] br[22] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_23 bl[23] br[23] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_24 bl[24] br[24] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_25 bl[25] br[25] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_26 bl[26] br[26] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_27 bl[27] br[27] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_28 bl[28] br[28] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_29 bl[29] br[29] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_30 bl[30] br[30] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_31 bl[31] br[31] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_32 bl[32] br[32] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_33 bl[33] br[33] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_34 bl[34] br[34] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_35 bl[35] br[35] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_36 bl[36] br[36] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_37 bl[37] br[37] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_38 bl[38] br[38] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_39 bl[39] br[39] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_40 bl[40] br[40] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_41 bl[41] br[41] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_42 bl[42] br[42] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_43 bl[43] br[43] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_44 bl[44] br[44] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_45 bl[45] br[45] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_46 bl[46] br[46] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_47 bl[47] br[47] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_48 bl[48] br[48] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_49 bl[49] br[49] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_50 bl[50] br[50] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_51 bl[51] br[51] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_52 bl[52] br[52] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_53 bl[53] br[53] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_54 bl[54] br[54] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_55 bl[55] br[55] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_56 bl[56] br[56] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_57 bl[57] br[57] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_58 bl[58] br[58] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_59 bl[59] br[59] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_60 bl[60] br[60] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_61 bl[61] br[61] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_62 bl[62] br[62] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_63 bl[63] br[63] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_106_0 bl[0] br[0] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_1 bl[1] br[1] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_2 bl[2] br[2] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_3 bl[3] br[3] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_4 bl[4] br[4] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_5 bl[5] br[5] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_6 bl[6] br[6] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_7 bl[7] br[7] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_8 bl[8] br[8] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_9 bl[9] br[9] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_10 bl[10] br[10] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_11 bl[11] br[11] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_12 bl[12] br[12] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_13 bl[13] br[13] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_14 bl[14] br[14] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_15 bl[15] br[15] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_16 bl[16] br[16] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_17 bl[17] br[17] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_18 bl[18] br[18] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_19 bl[19] br[19] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_20 bl[20] br[20] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_21 bl[21] br[21] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_22 bl[22] br[22] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_23 bl[23] br[23] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_24 bl[24] br[24] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_25 bl[25] br[25] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_26 bl[26] br[26] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_27 bl[27] br[27] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_28 bl[28] br[28] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_29 bl[29] br[29] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_30 bl[30] br[30] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_31 bl[31] br[31] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_32 bl[32] br[32] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_33 bl[33] br[33] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_34 bl[34] br[34] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_35 bl[35] br[35] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_36 bl[36] br[36] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_37 bl[37] br[37] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_38 bl[38] br[38] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_39 bl[39] br[39] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_40 bl[40] br[40] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_41 bl[41] br[41] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_42 bl[42] br[42] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_43 bl[43] br[43] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_44 bl[44] br[44] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_45 bl[45] br[45] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_46 bl[46] br[46] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_47 bl[47] br[47] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_48 bl[48] br[48] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_49 bl[49] br[49] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_50 bl[50] br[50] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_51 bl[51] br[51] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_52 bl[52] br[52] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_53 bl[53] br[53] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_54 bl[54] br[54] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_55 bl[55] br[55] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_56 bl[56] br[56] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_57 bl[57] br[57] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_58 bl[58] br[58] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_59 bl[59] br[59] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_60 bl[60] br[60] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_61 bl[61] br[61] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_62 bl[62] br[62] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_63 bl[63] br[63] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_107_0 bl[0] br[0] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_1 bl[1] br[1] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_2 bl[2] br[2] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_3 bl[3] br[3] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_4 bl[4] br[4] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_5 bl[5] br[5] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_6 bl[6] br[6] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_7 bl[7] br[7] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_8 bl[8] br[8] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_9 bl[9] br[9] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_10 bl[10] br[10] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_11 bl[11] br[11] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_12 bl[12] br[12] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_13 bl[13] br[13] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_14 bl[14] br[14] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_15 bl[15] br[15] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_16 bl[16] br[16] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_17 bl[17] br[17] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_18 bl[18] br[18] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_19 bl[19] br[19] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_20 bl[20] br[20] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_21 bl[21] br[21] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_22 bl[22] br[22] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_23 bl[23] br[23] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_24 bl[24] br[24] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_25 bl[25] br[25] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_26 bl[26] br[26] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_27 bl[27] br[27] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_28 bl[28] br[28] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_29 bl[29] br[29] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_30 bl[30] br[30] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_31 bl[31] br[31] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_32 bl[32] br[32] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_33 bl[33] br[33] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_34 bl[34] br[34] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_35 bl[35] br[35] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_36 bl[36] br[36] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_37 bl[37] br[37] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_38 bl[38] br[38] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_39 bl[39] br[39] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_40 bl[40] br[40] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_41 bl[41] br[41] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_42 bl[42] br[42] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_43 bl[43] br[43] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_44 bl[44] br[44] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_45 bl[45] br[45] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_46 bl[46] br[46] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_47 bl[47] br[47] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_48 bl[48] br[48] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_49 bl[49] br[49] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_50 bl[50] br[50] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_51 bl[51] br[51] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_52 bl[52] br[52] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_53 bl[53] br[53] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_54 bl[54] br[54] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_55 bl[55] br[55] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_56 bl[56] br[56] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_57 bl[57] br[57] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_58 bl[58] br[58] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_59 bl[59] br[59] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_60 bl[60] br[60] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_61 bl[61] br[61] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_62 bl[62] br[62] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_63 bl[63] br[63] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_108_0 bl[0] br[0] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_1 bl[1] br[1] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_2 bl[2] br[2] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_3 bl[3] br[3] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_4 bl[4] br[4] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_5 bl[5] br[5] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_6 bl[6] br[6] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_7 bl[7] br[7] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_8 bl[8] br[8] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_9 bl[9] br[9] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_10 bl[10] br[10] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_11 bl[11] br[11] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_12 bl[12] br[12] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_13 bl[13] br[13] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_14 bl[14] br[14] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_15 bl[15] br[15] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_16 bl[16] br[16] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_17 bl[17] br[17] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_18 bl[18] br[18] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_19 bl[19] br[19] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_20 bl[20] br[20] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_21 bl[21] br[21] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_22 bl[22] br[22] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_23 bl[23] br[23] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_24 bl[24] br[24] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_25 bl[25] br[25] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_26 bl[26] br[26] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_27 bl[27] br[27] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_28 bl[28] br[28] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_29 bl[29] br[29] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_30 bl[30] br[30] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_31 bl[31] br[31] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_32 bl[32] br[32] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_33 bl[33] br[33] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_34 bl[34] br[34] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_35 bl[35] br[35] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_36 bl[36] br[36] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_37 bl[37] br[37] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_38 bl[38] br[38] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_39 bl[39] br[39] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_40 bl[40] br[40] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_41 bl[41] br[41] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_42 bl[42] br[42] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_43 bl[43] br[43] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_44 bl[44] br[44] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_45 bl[45] br[45] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_46 bl[46] br[46] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_47 bl[47] br[47] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_48 bl[48] br[48] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_49 bl[49] br[49] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_50 bl[50] br[50] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_51 bl[51] br[51] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_52 bl[52] br[52] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_53 bl[53] br[53] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_54 bl[54] br[54] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_55 bl[55] br[55] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_56 bl[56] br[56] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_57 bl[57] br[57] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_58 bl[58] br[58] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_59 bl[59] br[59] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_60 bl[60] br[60] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_61 bl[61] br[61] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_62 bl[62] br[62] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_63 bl[63] br[63] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_109_0 bl[0] br[0] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_1 bl[1] br[1] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_2 bl[2] br[2] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_3 bl[3] br[3] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_4 bl[4] br[4] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_5 bl[5] br[5] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_6 bl[6] br[6] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_7 bl[7] br[7] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_8 bl[8] br[8] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_9 bl[9] br[9] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_10 bl[10] br[10] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_11 bl[11] br[11] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_12 bl[12] br[12] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_13 bl[13] br[13] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_14 bl[14] br[14] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_15 bl[15] br[15] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_16 bl[16] br[16] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_17 bl[17] br[17] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_18 bl[18] br[18] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_19 bl[19] br[19] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_20 bl[20] br[20] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_21 bl[21] br[21] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_22 bl[22] br[22] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_23 bl[23] br[23] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_24 bl[24] br[24] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_25 bl[25] br[25] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_26 bl[26] br[26] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_27 bl[27] br[27] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_28 bl[28] br[28] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_29 bl[29] br[29] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_30 bl[30] br[30] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_31 bl[31] br[31] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_32 bl[32] br[32] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_33 bl[33] br[33] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_34 bl[34] br[34] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_35 bl[35] br[35] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_36 bl[36] br[36] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_37 bl[37] br[37] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_38 bl[38] br[38] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_39 bl[39] br[39] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_40 bl[40] br[40] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_41 bl[41] br[41] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_42 bl[42] br[42] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_43 bl[43] br[43] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_44 bl[44] br[44] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_45 bl[45] br[45] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_46 bl[46] br[46] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_47 bl[47] br[47] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_48 bl[48] br[48] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_49 bl[49] br[49] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_50 bl[50] br[50] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_51 bl[51] br[51] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_52 bl[52] br[52] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_53 bl[53] br[53] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_54 bl[54] br[54] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_55 bl[55] br[55] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_56 bl[56] br[56] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_57 bl[57] br[57] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_58 bl[58] br[58] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_59 bl[59] br[59] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_60 bl[60] br[60] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_61 bl[61] br[61] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_62 bl[62] br[62] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_63 bl[63] br[63] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_110_0 bl[0] br[0] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_1 bl[1] br[1] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_2 bl[2] br[2] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_3 bl[3] br[3] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_4 bl[4] br[4] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_5 bl[5] br[5] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_6 bl[6] br[6] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_7 bl[7] br[7] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_8 bl[8] br[8] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_9 bl[9] br[9] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_10 bl[10] br[10] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_11 bl[11] br[11] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_12 bl[12] br[12] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_13 bl[13] br[13] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_14 bl[14] br[14] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_15 bl[15] br[15] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_16 bl[16] br[16] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_17 bl[17] br[17] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_18 bl[18] br[18] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_19 bl[19] br[19] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_20 bl[20] br[20] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_21 bl[21] br[21] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_22 bl[22] br[22] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_23 bl[23] br[23] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_24 bl[24] br[24] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_25 bl[25] br[25] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_26 bl[26] br[26] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_27 bl[27] br[27] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_28 bl[28] br[28] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_29 bl[29] br[29] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_30 bl[30] br[30] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_31 bl[31] br[31] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_32 bl[32] br[32] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_33 bl[33] br[33] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_34 bl[34] br[34] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_35 bl[35] br[35] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_36 bl[36] br[36] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_37 bl[37] br[37] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_38 bl[38] br[38] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_39 bl[39] br[39] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_40 bl[40] br[40] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_41 bl[41] br[41] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_42 bl[42] br[42] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_43 bl[43] br[43] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_44 bl[44] br[44] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_45 bl[45] br[45] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_46 bl[46] br[46] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_47 bl[47] br[47] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_48 bl[48] br[48] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_49 bl[49] br[49] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_50 bl[50] br[50] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_51 bl[51] br[51] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_52 bl[52] br[52] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_53 bl[53] br[53] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_54 bl[54] br[54] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_55 bl[55] br[55] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_56 bl[56] br[56] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_57 bl[57] br[57] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_58 bl[58] br[58] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_59 bl[59] br[59] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_60 bl[60] br[60] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_61 bl[61] br[61] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_62 bl[62] br[62] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_63 bl[63] br[63] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_111_0 bl[0] br[0] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_1 bl[1] br[1] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_2 bl[2] br[2] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_3 bl[3] br[3] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_4 bl[4] br[4] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_5 bl[5] br[5] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_6 bl[6] br[6] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_7 bl[7] br[7] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_8 bl[8] br[8] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_9 bl[9] br[9] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_10 bl[10] br[10] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_11 bl[11] br[11] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_12 bl[12] br[12] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_13 bl[13] br[13] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_14 bl[14] br[14] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_15 bl[15] br[15] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_16 bl[16] br[16] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_17 bl[17] br[17] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_18 bl[18] br[18] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_19 bl[19] br[19] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_20 bl[20] br[20] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_21 bl[21] br[21] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_22 bl[22] br[22] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_23 bl[23] br[23] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_24 bl[24] br[24] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_25 bl[25] br[25] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_26 bl[26] br[26] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_27 bl[27] br[27] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_28 bl[28] br[28] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_29 bl[29] br[29] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_30 bl[30] br[30] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_31 bl[31] br[31] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_32 bl[32] br[32] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_33 bl[33] br[33] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_34 bl[34] br[34] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_35 bl[35] br[35] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_36 bl[36] br[36] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_37 bl[37] br[37] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_38 bl[38] br[38] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_39 bl[39] br[39] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_40 bl[40] br[40] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_41 bl[41] br[41] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_42 bl[42] br[42] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_43 bl[43] br[43] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_44 bl[44] br[44] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_45 bl[45] br[45] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_46 bl[46] br[46] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_47 bl[47] br[47] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_48 bl[48] br[48] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_49 bl[49] br[49] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_50 bl[50] br[50] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_51 bl[51] br[51] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_52 bl[52] br[52] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_53 bl[53] br[53] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_54 bl[54] br[54] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_55 bl[55] br[55] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_56 bl[56] br[56] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_57 bl[57] br[57] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_58 bl[58] br[58] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_59 bl[59] br[59] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_60 bl[60] br[60] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_61 bl[61] br[61] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_62 bl[62] br[62] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_63 bl[63] br[63] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_112_0 bl[0] br[0] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_1 bl[1] br[1] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_2 bl[2] br[2] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_3 bl[3] br[3] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_4 bl[4] br[4] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_5 bl[5] br[5] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_6 bl[6] br[6] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_7 bl[7] br[7] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_8 bl[8] br[8] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_9 bl[9] br[9] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_10 bl[10] br[10] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_11 bl[11] br[11] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_12 bl[12] br[12] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_13 bl[13] br[13] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_14 bl[14] br[14] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_15 bl[15] br[15] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_16 bl[16] br[16] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_17 bl[17] br[17] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_18 bl[18] br[18] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_19 bl[19] br[19] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_20 bl[20] br[20] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_21 bl[21] br[21] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_22 bl[22] br[22] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_23 bl[23] br[23] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_24 bl[24] br[24] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_25 bl[25] br[25] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_26 bl[26] br[26] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_27 bl[27] br[27] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_28 bl[28] br[28] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_29 bl[29] br[29] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_30 bl[30] br[30] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_31 bl[31] br[31] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_32 bl[32] br[32] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_33 bl[33] br[33] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_34 bl[34] br[34] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_35 bl[35] br[35] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_36 bl[36] br[36] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_37 bl[37] br[37] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_38 bl[38] br[38] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_39 bl[39] br[39] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_40 bl[40] br[40] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_41 bl[41] br[41] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_42 bl[42] br[42] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_43 bl[43] br[43] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_44 bl[44] br[44] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_45 bl[45] br[45] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_46 bl[46] br[46] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_47 bl[47] br[47] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_48 bl[48] br[48] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_49 bl[49] br[49] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_50 bl[50] br[50] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_51 bl[51] br[51] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_52 bl[52] br[52] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_53 bl[53] br[53] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_54 bl[54] br[54] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_55 bl[55] br[55] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_56 bl[56] br[56] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_57 bl[57] br[57] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_58 bl[58] br[58] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_59 bl[59] br[59] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_60 bl[60] br[60] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_61 bl[61] br[61] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_62 bl[62] br[62] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_63 bl[63] br[63] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_113_0 bl[0] br[0] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_1 bl[1] br[1] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_2 bl[2] br[2] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_3 bl[3] br[3] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_4 bl[4] br[4] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_5 bl[5] br[5] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_6 bl[6] br[6] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_7 bl[7] br[7] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_8 bl[8] br[8] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_9 bl[9] br[9] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_10 bl[10] br[10] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_11 bl[11] br[11] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_12 bl[12] br[12] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_13 bl[13] br[13] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_14 bl[14] br[14] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_15 bl[15] br[15] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_16 bl[16] br[16] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_17 bl[17] br[17] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_18 bl[18] br[18] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_19 bl[19] br[19] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_20 bl[20] br[20] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_21 bl[21] br[21] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_22 bl[22] br[22] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_23 bl[23] br[23] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_24 bl[24] br[24] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_25 bl[25] br[25] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_26 bl[26] br[26] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_27 bl[27] br[27] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_28 bl[28] br[28] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_29 bl[29] br[29] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_30 bl[30] br[30] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_31 bl[31] br[31] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_32 bl[32] br[32] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_33 bl[33] br[33] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_34 bl[34] br[34] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_35 bl[35] br[35] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_36 bl[36] br[36] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_37 bl[37] br[37] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_38 bl[38] br[38] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_39 bl[39] br[39] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_40 bl[40] br[40] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_41 bl[41] br[41] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_42 bl[42] br[42] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_43 bl[43] br[43] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_44 bl[44] br[44] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_45 bl[45] br[45] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_46 bl[46] br[46] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_47 bl[47] br[47] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_48 bl[48] br[48] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_49 bl[49] br[49] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_50 bl[50] br[50] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_51 bl[51] br[51] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_52 bl[52] br[52] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_53 bl[53] br[53] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_54 bl[54] br[54] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_55 bl[55] br[55] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_56 bl[56] br[56] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_57 bl[57] br[57] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_58 bl[58] br[58] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_59 bl[59] br[59] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_60 bl[60] br[60] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_61 bl[61] br[61] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_62 bl[62] br[62] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_63 bl[63] br[63] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_114_0 bl[0] br[0] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_1 bl[1] br[1] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_2 bl[2] br[2] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_3 bl[3] br[3] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_4 bl[4] br[4] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_5 bl[5] br[5] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_6 bl[6] br[6] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_7 bl[7] br[7] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_8 bl[8] br[8] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_9 bl[9] br[9] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_10 bl[10] br[10] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_11 bl[11] br[11] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_12 bl[12] br[12] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_13 bl[13] br[13] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_14 bl[14] br[14] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_15 bl[15] br[15] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_16 bl[16] br[16] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_17 bl[17] br[17] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_18 bl[18] br[18] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_19 bl[19] br[19] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_20 bl[20] br[20] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_21 bl[21] br[21] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_22 bl[22] br[22] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_23 bl[23] br[23] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_24 bl[24] br[24] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_25 bl[25] br[25] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_26 bl[26] br[26] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_27 bl[27] br[27] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_28 bl[28] br[28] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_29 bl[29] br[29] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_30 bl[30] br[30] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_31 bl[31] br[31] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_32 bl[32] br[32] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_33 bl[33] br[33] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_34 bl[34] br[34] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_35 bl[35] br[35] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_36 bl[36] br[36] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_37 bl[37] br[37] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_38 bl[38] br[38] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_39 bl[39] br[39] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_40 bl[40] br[40] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_41 bl[41] br[41] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_42 bl[42] br[42] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_43 bl[43] br[43] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_44 bl[44] br[44] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_45 bl[45] br[45] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_46 bl[46] br[46] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_47 bl[47] br[47] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_48 bl[48] br[48] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_49 bl[49] br[49] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_50 bl[50] br[50] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_51 bl[51] br[51] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_52 bl[52] br[52] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_53 bl[53] br[53] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_54 bl[54] br[54] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_55 bl[55] br[55] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_56 bl[56] br[56] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_57 bl[57] br[57] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_58 bl[58] br[58] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_59 bl[59] br[59] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_60 bl[60] br[60] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_61 bl[61] br[61] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_62 bl[62] br[62] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_63 bl[63] br[63] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_115_0 bl[0] br[0] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_1 bl[1] br[1] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_2 bl[2] br[2] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_3 bl[3] br[3] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_4 bl[4] br[4] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_5 bl[5] br[5] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_6 bl[6] br[6] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_7 bl[7] br[7] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_8 bl[8] br[8] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_9 bl[9] br[9] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_10 bl[10] br[10] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_11 bl[11] br[11] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_12 bl[12] br[12] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_13 bl[13] br[13] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_14 bl[14] br[14] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_15 bl[15] br[15] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_16 bl[16] br[16] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_17 bl[17] br[17] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_18 bl[18] br[18] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_19 bl[19] br[19] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_20 bl[20] br[20] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_21 bl[21] br[21] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_22 bl[22] br[22] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_23 bl[23] br[23] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_24 bl[24] br[24] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_25 bl[25] br[25] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_26 bl[26] br[26] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_27 bl[27] br[27] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_28 bl[28] br[28] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_29 bl[29] br[29] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_30 bl[30] br[30] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_31 bl[31] br[31] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_32 bl[32] br[32] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_33 bl[33] br[33] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_34 bl[34] br[34] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_35 bl[35] br[35] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_36 bl[36] br[36] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_37 bl[37] br[37] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_38 bl[38] br[38] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_39 bl[39] br[39] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_40 bl[40] br[40] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_41 bl[41] br[41] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_42 bl[42] br[42] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_43 bl[43] br[43] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_44 bl[44] br[44] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_45 bl[45] br[45] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_46 bl[46] br[46] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_47 bl[47] br[47] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_48 bl[48] br[48] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_49 bl[49] br[49] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_50 bl[50] br[50] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_51 bl[51] br[51] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_52 bl[52] br[52] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_53 bl[53] br[53] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_54 bl[54] br[54] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_55 bl[55] br[55] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_56 bl[56] br[56] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_57 bl[57] br[57] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_58 bl[58] br[58] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_59 bl[59] br[59] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_60 bl[60] br[60] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_61 bl[61] br[61] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_62 bl[62] br[62] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_63 bl[63] br[63] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_116_0 bl[0] br[0] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_1 bl[1] br[1] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_2 bl[2] br[2] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_3 bl[3] br[3] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_4 bl[4] br[4] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_5 bl[5] br[5] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_6 bl[6] br[6] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_7 bl[7] br[7] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_8 bl[8] br[8] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_9 bl[9] br[9] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_10 bl[10] br[10] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_11 bl[11] br[11] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_12 bl[12] br[12] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_13 bl[13] br[13] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_14 bl[14] br[14] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_15 bl[15] br[15] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_16 bl[16] br[16] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_17 bl[17] br[17] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_18 bl[18] br[18] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_19 bl[19] br[19] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_20 bl[20] br[20] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_21 bl[21] br[21] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_22 bl[22] br[22] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_23 bl[23] br[23] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_24 bl[24] br[24] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_25 bl[25] br[25] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_26 bl[26] br[26] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_27 bl[27] br[27] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_28 bl[28] br[28] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_29 bl[29] br[29] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_30 bl[30] br[30] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_31 bl[31] br[31] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_32 bl[32] br[32] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_33 bl[33] br[33] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_34 bl[34] br[34] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_35 bl[35] br[35] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_36 bl[36] br[36] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_37 bl[37] br[37] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_38 bl[38] br[38] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_39 bl[39] br[39] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_40 bl[40] br[40] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_41 bl[41] br[41] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_42 bl[42] br[42] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_43 bl[43] br[43] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_44 bl[44] br[44] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_45 bl[45] br[45] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_46 bl[46] br[46] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_47 bl[47] br[47] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_48 bl[48] br[48] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_49 bl[49] br[49] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_50 bl[50] br[50] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_51 bl[51] br[51] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_52 bl[52] br[52] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_53 bl[53] br[53] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_54 bl[54] br[54] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_55 bl[55] br[55] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_56 bl[56] br[56] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_57 bl[57] br[57] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_58 bl[58] br[58] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_59 bl[59] br[59] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_60 bl[60] br[60] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_61 bl[61] br[61] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_62 bl[62] br[62] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_63 bl[63] br[63] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_117_0 bl[0] br[0] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_1 bl[1] br[1] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_2 bl[2] br[2] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_3 bl[3] br[3] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_4 bl[4] br[4] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_5 bl[5] br[5] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_6 bl[6] br[6] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_7 bl[7] br[7] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_8 bl[8] br[8] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_9 bl[9] br[9] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_10 bl[10] br[10] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_11 bl[11] br[11] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_12 bl[12] br[12] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_13 bl[13] br[13] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_14 bl[14] br[14] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_15 bl[15] br[15] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_16 bl[16] br[16] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_17 bl[17] br[17] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_18 bl[18] br[18] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_19 bl[19] br[19] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_20 bl[20] br[20] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_21 bl[21] br[21] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_22 bl[22] br[22] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_23 bl[23] br[23] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_24 bl[24] br[24] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_25 bl[25] br[25] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_26 bl[26] br[26] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_27 bl[27] br[27] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_28 bl[28] br[28] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_29 bl[29] br[29] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_30 bl[30] br[30] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_31 bl[31] br[31] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_32 bl[32] br[32] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_33 bl[33] br[33] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_34 bl[34] br[34] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_35 bl[35] br[35] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_36 bl[36] br[36] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_37 bl[37] br[37] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_38 bl[38] br[38] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_39 bl[39] br[39] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_40 bl[40] br[40] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_41 bl[41] br[41] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_42 bl[42] br[42] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_43 bl[43] br[43] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_44 bl[44] br[44] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_45 bl[45] br[45] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_46 bl[46] br[46] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_47 bl[47] br[47] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_48 bl[48] br[48] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_49 bl[49] br[49] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_50 bl[50] br[50] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_51 bl[51] br[51] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_52 bl[52] br[52] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_53 bl[53] br[53] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_54 bl[54] br[54] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_55 bl[55] br[55] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_56 bl[56] br[56] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_57 bl[57] br[57] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_58 bl[58] br[58] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_59 bl[59] br[59] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_60 bl[60] br[60] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_61 bl[61] br[61] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_62 bl[62] br[62] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_63 bl[63] br[63] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_118_0 bl[0] br[0] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_1 bl[1] br[1] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_2 bl[2] br[2] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_3 bl[3] br[3] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_4 bl[4] br[4] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_5 bl[5] br[5] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_6 bl[6] br[6] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_7 bl[7] br[7] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_8 bl[8] br[8] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_9 bl[9] br[9] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_10 bl[10] br[10] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_11 bl[11] br[11] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_12 bl[12] br[12] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_13 bl[13] br[13] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_14 bl[14] br[14] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_15 bl[15] br[15] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_16 bl[16] br[16] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_17 bl[17] br[17] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_18 bl[18] br[18] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_19 bl[19] br[19] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_20 bl[20] br[20] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_21 bl[21] br[21] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_22 bl[22] br[22] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_23 bl[23] br[23] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_24 bl[24] br[24] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_25 bl[25] br[25] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_26 bl[26] br[26] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_27 bl[27] br[27] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_28 bl[28] br[28] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_29 bl[29] br[29] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_30 bl[30] br[30] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_31 bl[31] br[31] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_32 bl[32] br[32] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_33 bl[33] br[33] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_34 bl[34] br[34] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_35 bl[35] br[35] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_36 bl[36] br[36] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_37 bl[37] br[37] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_38 bl[38] br[38] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_39 bl[39] br[39] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_40 bl[40] br[40] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_41 bl[41] br[41] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_42 bl[42] br[42] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_43 bl[43] br[43] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_44 bl[44] br[44] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_45 bl[45] br[45] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_46 bl[46] br[46] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_47 bl[47] br[47] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_48 bl[48] br[48] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_49 bl[49] br[49] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_50 bl[50] br[50] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_51 bl[51] br[51] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_52 bl[52] br[52] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_53 bl[53] br[53] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_54 bl[54] br[54] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_55 bl[55] br[55] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_56 bl[56] br[56] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_57 bl[57] br[57] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_58 bl[58] br[58] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_59 bl[59] br[59] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_60 bl[60] br[60] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_61 bl[61] br[61] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_62 bl[62] br[62] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_63 bl[63] br[63] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_119_0 bl[0] br[0] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_1 bl[1] br[1] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_2 bl[2] br[2] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_3 bl[3] br[3] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_4 bl[4] br[4] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_5 bl[5] br[5] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_6 bl[6] br[6] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_7 bl[7] br[7] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_8 bl[8] br[8] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_9 bl[9] br[9] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_10 bl[10] br[10] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_11 bl[11] br[11] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_12 bl[12] br[12] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_13 bl[13] br[13] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_14 bl[14] br[14] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_15 bl[15] br[15] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_16 bl[16] br[16] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_17 bl[17] br[17] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_18 bl[18] br[18] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_19 bl[19] br[19] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_20 bl[20] br[20] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_21 bl[21] br[21] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_22 bl[22] br[22] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_23 bl[23] br[23] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_24 bl[24] br[24] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_25 bl[25] br[25] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_26 bl[26] br[26] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_27 bl[27] br[27] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_28 bl[28] br[28] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_29 bl[29] br[29] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_30 bl[30] br[30] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_31 bl[31] br[31] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_32 bl[32] br[32] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_33 bl[33] br[33] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_34 bl[34] br[34] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_35 bl[35] br[35] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_36 bl[36] br[36] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_37 bl[37] br[37] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_38 bl[38] br[38] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_39 bl[39] br[39] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_40 bl[40] br[40] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_41 bl[41] br[41] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_42 bl[42] br[42] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_43 bl[43] br[43] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_44 bl[44] br[44] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_45 bl[45] br[45] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_46 bl[46] br[46] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_47 bl[47] br[47] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_48 bl[48] br[48] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_49 bl[49] br[49] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_50 bl[50] br[50] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_51 bl[51] br[51] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_52 bl[52] br[52] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_53 bl[53] br[53] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_54 bl[54] br[54] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_55 bl[55] br[55] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_56 bl[56] br[56] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_57 bl[57] br[57] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_58 bl[58] br[58] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_59 bl[59] br[59] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_60 bl[60] br[60] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_61 bl[61] br[61] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_62 bl[62] br[62] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_63 bl[63] br[63] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_120_0 bl[0] br[0] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_1 bl[1] br[1] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_2 bl[2] br[2] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_3 bl[3] br[3] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_4 bl[4] br[4] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_5 bl[5] br[5] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_6 bl[6] br[6] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_7 bl[7] br[7] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_8 bl[8] br[8] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_9 bl[9] br[9] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_10 bl[10] br[10] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_11 bl[11] br[11] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_12 bl[12] br[12] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_13 bl[13] br[13] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_14 bl[14] br[14] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_15 bl[15] br[15] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_16 bl[16] br[16] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_17 bl[17] br[17] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_18 bl[18] br[18] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_19 bl[19] br[19] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_20 bl[20] br[20] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_21 bl[21] br[21] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_22 bl[22] br[22] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_23 bl[23] br[23] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_24 bl[24] br[24] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_25 bl[25] br[25] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_26 bl[26] br[26] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_27 bl[27] br[27] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_28 bl[28] br[28] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_29 bl[29] br[29] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_30 bl[30] br[30] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_31 bl[31] br[31] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_32 bl[32] br[32] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_33 bl[33] br[33] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_34 bl[34] br[34] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_35 bl[35] br[35] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_36 bl[36] br[36] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_37 bl[37] br[37] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_38 bl[38] br[38] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_39 bl[39] br[39] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_40 bl[40] br[40] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_41 bl[41] br[41] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_42 bl[42] br[42] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_43 bl[43] br[43] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_44 bl[44] br[44] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_45 bl[45] br[45] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_46 bl[46] br[46] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_47 bl[47] br[47] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_48 bl[48] br[48] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_49 bl[49] br[49] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_50 bl[50] br[50] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_51 bl[51] br[51] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_52 bl[52] br[52] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_53 bl[53] br[53] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_54 bl[54] br[54] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_55 bl[55] br[55] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_56 bl[56] br[56] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_57 bl[57] br[57] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_58 bl[58] br[58] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_59 bl[59] br[59] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_60 bl[60] br[60] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_61 bl[61] br[61] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_62 bl[62] br[62] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_63 bl[63] br[63] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_121_0 bl[0] br[0] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_1 bl[1] br[1] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_2 bl[2] br[2] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_3 bl[3] br[3] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_4 bl[4] br[4] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_5 bl[5] br[5] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_6 bl[6] br[6] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_7 bl[7] br[7] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_8 bl[8] br[8] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_9 bl[9] br[9] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_10 bl[10] br[10] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_11 bl[11] br[11] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_12 bl[12] br[12] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_13 bl[13] br[13] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_14 bl[14] br[14] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_15 bl[15] br[15] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_16 bl[16] br[16] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_17 bl[17] br[17] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_18 bl[18] br[18] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_19 bl[19] br[19] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_20 bl[20] br[20] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_21 bl[21] br[21] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_22 bl[22] br[22] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_23 bl[23] br[23] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_24 bl[24] br[24] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_25 bl[25] br[25] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_26 bl[26] br[26] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_27 bl[27] br[27] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_28 bl[28] br[28] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_29 bl[29] br[29] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_30 bl[30] br[30] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_31 bl[31] br[31] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_32 bl[32] br[32] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_33 bl[33] br[33] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_34 bl[34] br[34] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_35 bl[35] br[35] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_36 bl[36] br[36] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_37 bl[37] br[37] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_38 bl[38] br[38] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_39 bl[39] br[39] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_40 bl[40] br[40] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_41 bl[41] br[41] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_42 bl[42] br[42] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_43 bl[43] br[43] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_44 bl[44] br[44] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_45 bl[45] br[45] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_46 bl[46] br[46] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_47 bl[47] br[47] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_48 bl[48] br[48] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_49 bl[49] br[49] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_50 bl[50] br[50] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_51 bl[51] br[51] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_52 bl[52] br[52] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_53 bl[53] br[53] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_54 bl[54] br[54] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_55 bl[55] br[55] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_56 bl[56] br[56] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_57 bl[57] br[57] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_58 bl[58] br[58] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_59 bl[59] br[59] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_60 bl[60] br[60] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_61 bl[61] br[61] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_62 bl[62] br[62] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_63 bl[63] br[63] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_122_0 bl[0] br[0] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_1 bl[1] br[1] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_2 bl[2] br[2] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_3 bl[3] br[3] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_4 bl[4] br[4] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_5 bl[5] br[5] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_6 bl[6] br[6] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_7 bl[7] br[7] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_8 bl[8] br[8] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_9 bl[9] br[9] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_10 bl[10] br[10] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_11 bl[11] br[11] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_12 bl[12] br[12] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_13 bl[13] br[13] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_14 bl[14] br[14] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_15 bl[15] br[15] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_16 bl[16] br[16] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_17 bl[17] br[17] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_18 bl[18] br[18] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_19 bl[19] br[19] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_20 bl[20] br[20] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_21 bl[21] br[21] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_22 bl[22] br[22] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_23 bl[23] br[23] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_24 bl[24] br[24] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_25 bl[25] br[25] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_26 bl[26] br[26] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_27 bl[27] br[27] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_28 bl[28] br[28] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_29 bl[29] br[29] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_30 bl[30] br[30] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_31 bl[31] br[31] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_32 bl[32] br[32] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_33 bl[33] br[33] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_34 bl[34] br[34] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_35 bl[35] br[35] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_36 bl[36] br[36] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_37 bl[37] br[37] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_38 bl[38] br[38] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_39 bl[39] br[39] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_40 bl[40] br[40] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_41 bl[41] br[41] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_42 bl[42] br[42] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_43 bl[43] br[43] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_44 bl[44] br[44] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_45 bl[45] br[45] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_46 bl[46] br[46] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_47 bl[47] br[47] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_48 bl[48] br[48] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_49 bl[49] br[49] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_50 bl[50] br[50] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_51 bl[51] br[51] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_52 bl[52] br[52] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_53 bl[53] br[53] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_54 bl[54] br[54] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_55 bl[55] br[55] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_56 bl[56] br[56] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_57 bl[57] br[57] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_58 bl[58] br[58] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_59 bl[59] br[59] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_60 bl[60] br[60] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_61 bl[61] br[61] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_62 bl[62] br[62] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_63 bl[63] br[63] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_123_0 bl[0] br[0] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_1 bl[1] br[1] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_2 bl[2] br[2] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_3 bl[3] br[3] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_4 bl[4] br[4] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_5 bl[5] br[5] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_6 bl[6] br[6] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_7 bl[7] br[7] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_8 bl[8] br[8] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_9 bl[9] br[9] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_10 bl[10] br[10] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_11 bl[11] br[11] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_12 bl[12] br[12] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_13 bl[13] br[13] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_14 bl[14] br[14] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_15 bl[15] br[15] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_16 bl[16] br[16] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_17 bl[17] br[17] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_18 bl[18] br[18] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_19 bl[19] br[19] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_20 bl[20] br[20] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_21 bl[21] br[21] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_22 bl[22] br[22] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_23 bl[23] br[23] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_24 bl[24] br[24] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_25 bl[25] br[25] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_26 bl[26] br[26] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_27 bl[27] br[27] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_28 bl[28] br[28] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_29 bl[29] br[29] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_30 bl[30] br[30] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_31 bl[31] br[31] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_32 bl[32] br[32] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_33 bl[33] br[33] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_34 bl[34] br[34] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_35 bl[35] br[35] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_36 bl[36] br[36] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_37 bl[37] br[37] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_38 bl[38] br[38] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_39 bl[39] br[39] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_40 bl[40] br[40] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_41 bl[41] br[41] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_42 bl[42] br[42] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_43 bl[43] br[43] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_44 bl[44] br[44] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_45 bl[45] br[45] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_46 bl[46] br[46] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_47 bl[47] br[47] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_48 bl[48] br[48] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_49 bl[49] br[49] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_50 bl[50] br[50] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_51 bl[51] br[51] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_52 bl[52] br[52] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_53 bl[53] br[53] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_54 bl[54] br[54] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_55 bl[55] br[55] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_56 bl[56] br[56] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_57 bl[57] br[57] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_58 bl[58] br[58] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_59 bl[59] br[59] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_60 bl[60] br[60] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_61 bl[61] br[61] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_62 bl[62] br[62] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_63 bl[63] br[63] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_124_0 bl[0] br[0] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_1 bl[1] br[1] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_2 bl[2] br[2] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_3 bl[3] br[3] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_4 bl[4] br[4] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_5 bl[5] br[5] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_6 bl[6] br[6] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_7 bl[7] br[7] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_8 bl[8] br[8] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_9 bl[9] br[9] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_10 bl[10] br[10] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_11 bl[11] br[11] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_12 bl[12] br[12] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_13 bl[13] br[13] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_14 bl[14] br[14] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_15 bl[15] br[15] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_16 bl[16] br[16] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_17 bl[17] br[17] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_18 bl[18] br[18] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_19 bl[19] br[19] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_20 bl[20] br[20] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_21 bl[21] br[21] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_22 bl[22] br[22] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_23 bl[23] br[23] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_24 bl[24] br[24] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_25 bl[25] br[25] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_26 bl[26] br[26] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_27 bl[27] br[27] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_28 bl[28] br[28] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_29 bl[29] br[29] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_30 bl[30] br[30] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_31 bl[31] br[31] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_32 bl[32] br[32] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_33 bl[33] br[33] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_34 bl[34] br[34] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_35 bl[35] br[35] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_36 bl[36] br[36] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_37 bl[37] br[37] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_38 bl[38] br[38] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_39 bl[39] br[39] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_40 bl[40] br[40] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_41 bl[41] br[41] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_42 bl[42] br[42] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_43 bl[43] br[43] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_44 bl[44] br[44] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_45 bl[45] br[45] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_46 bl[46] br[46] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_47 bl[47] br[47] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_48 bl[48] br[48] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_49 bl[49] br[49] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_50 bl[50] br[50] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_51 bl[51] br[51] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_52 bl[52] br[52] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_53 bl[53] br[53] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_54 bl[54] br[54] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_55 bl[55] br[55] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_56 bl[56] br[56] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_57 bl[57] br[57] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_58 bl[58] br[58] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_59 bl[59] br[59] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_60 bl[60] br[60] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_61 bl[61] br[61] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_62 bl[62] br[62] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_63 bl[63] br[63] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_125_0 bl[0] br[0] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_1 bl[1] br[1] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_2 bl[2] br[2] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_3 bl[3] br[3] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_4 bl[4] br[4] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_5 bl[5] br[5] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_6 bl[6] br[6] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_7 bl[7] br[7] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_8 bl[8] br[8] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_9 bl[9] br[9] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_10 bl[10] br[10] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_11 bl[11] br[11] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_12 bl[12] br[12] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_13 bl[13] br[13] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_14 bl[14] br[14] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_15 bl[15] br[15] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_16 bl[16] br[16] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_17 bl[17] br[17] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_18 bl[18] br[18] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_19 bl[19] br[19] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_20 bl[20] br[20] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_21 bl[21] br[21] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_22 bl[22] br[22] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_23 bl[23] br[23] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_24 bl[24] br[24] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_25 bl[25] br[25] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_26 bl[26] br[26] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_27 bl[27] br[27] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_28 bl[28] br[28] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_29 bl[29] br[29] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_30 bl[30] br[30] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_31 bl[31] br[31] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_32 bl[32] br[32] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_33 bl[33] br[33] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_34 bl[34] br[34] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_35 bl[35] br[35] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_36 bl[36] br[36] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_37 bl[37] br[37] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_38 bl[38] br[38] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_39 bl[39] br[39] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_40 bl[40] br[40] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_41 bl[41] br[41] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_42 bl[42] br[42] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_43 bl[43] br[43] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_44 bl[44] br[44] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_45 bl[45] br[45] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_46 bl[46] br[46] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_47 bl[47] br[47] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_48 bl[48] br[48] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_49 bl[49] br[49] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_50 bl[50] br[50] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_51 bl[51] br[51] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_52 bl[52] br[52] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_53 bl[53] br[53] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_54 bl[54] br[54] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_55 bl[55] br[55] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_56 bl[56] br[56] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_57 bl[57] br[57] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_58 bl[58] br[58] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_59 bl[59] br[59] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_60 bl[60] br[60] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_61 bl[61] br[61] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_62 bl[62] br[62] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_63 bl[63] br[63] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_126_0 bl[0] br[0] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_1 bl[1] br[1] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_2 bl[2] br[2] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_3 bl[3] br[3] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_4 bl[4] br[4] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_5 bl[5] br[5] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_6 bl[6] br[6] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_7 bl[7] br[7] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_8 bl[8] br[8] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_9 bl[9] br[9] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_10 bl[10] br[10] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_11 bl[11] br[11] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_12 bl[12] br[12] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_13 bl[13] br[13] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_14 bl[14] br[14] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_15 bl[15] br[15] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_16 bl[16] br[16] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_17 bl[17] br[17] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_18 bl[18] br[18] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_19 bl[19] br[19] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_20 bl[20] br[20] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_21 bl[21] br[21] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_22 bl[22] br[22] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_23 bl[23] br[23] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_24 bl[24] br[24] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_25 bl[25] br[25] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_26 bl[26] br[26] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_27 bl[27] br[27] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_28 bl[28] br[28] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_29 bl[29] br[29] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_30 bl[30] br[30] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_31 bl[31] br[31] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_32 bl[32] br[32] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_33 bl[33] br[33] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_34 bl[34] br[34] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_35 bl[35] br[35] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_36 bl[36] br[36] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_37 bl[37] br[37] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_38 bl[38] br[38] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_39 bl[39] br[39] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_40 bl[40] br[40] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_41 bl[41] br[41] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_42 bl[42] br[42] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_43 bl[43] br[43] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_44 bl[44] br[44] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_45 bl[45] br[45] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_46 bl[46] br[46] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_47 bl[47] br[47] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_48 bl[48] br[48] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_49 bl[49] br[49] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_50 bl[50] br[50] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_51 bl[51] br[51] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_52 bl[52] br[52] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_53 bl[53] br[53] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_54 bl[54] br[54] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_55 bl[55] br[55] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_56 bl[56] br[56] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_57 bl[57] br[57] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_58 bl[58] br[58] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_59 bl[59] br[59] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_60 bl[60] br[60] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_61 bl[61] br[61] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_62 bl[62] br[62] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_63 bl[63] br[63] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_127_0 bl[0] br[0] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_1 bl[1] br[1] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_2 bl[2] br[2] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_3 bl[3] br[3] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_4 bl[4] br[4] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_5 bl[5] br[5] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_6 bl[6] br[6] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_7 bl[7] br[7] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_8 bl[8] br[8] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_9 bl[9] br[9] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_10 bl[10] br[10] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_11 bl[11] br[11] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_12 bl[12] br[12] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_13 bl[13] br[13] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_14 bl[14] br[14] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_15 bl[15] br[15] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_16 bl[16] br[16] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_17 bl[17] br[17] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_18 bl[18] br[18] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_19 bl[19] br[19] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_20 bl[20] br[20] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_21 bl[21] br[21] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_22 bl[22] br[22] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_23 bl[23] br[23] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_24 bl[24] br[24] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_25 bl[25] br[25] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_26 bl[26] br[26] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_27 bl[27] br[27] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_28 bl[28] br[28] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_29 bl[29] br[29] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_30 bl[30] br[30] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_31 bl[31] br[31] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_32 bl[32] br[32] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_33 bl[33] br[33] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_34 bl[34] br[34] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_35 bl[35] br[35] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_36 bl[36] br[36] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_37 bl[37] br[37] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_38 bl[38] br[38] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_39 bl[39] br[39] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_40 bl[40] br[40] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_41 bl[41] br[41] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_42 bl[42] br[42] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_43 bl[43] br[43] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_44 bl[44] br[44] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_45 bl[45] br[45] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_46 bl[46] br[46] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_47 bl[47] br[47] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_48 bl[48] br[48] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_49 bl[49] br[49] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_50 bl[50] br[50] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_51 bl[51] br[51] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_52 bl[52] br[52] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_53 bl[53] br[53] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_54 bl[54] br[54] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_55 bl[55] br[55] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_56 bl[56] br[56] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_57 bl[57] br[57] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_58 bl[58] br[58] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_59 bl[59] br[59] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_60 bl[60] br[60] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_61 bl[61] br[61] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_62 bl[62] br[62] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_63 bl[63] br[63] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_0 dummy_bl dummy_br vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_0 vdd vdd vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_1 dummy_bl dummy_br vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_1 vdd vdd vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_2 dummy_bl dummy_br vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_2 vdd vdd vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_3 dummy_bl dummy_br vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_3 vdd vdd vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_4 dummy_bl dummy_br vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_4 vdd vdd vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_5 dummy_bl dummy_br vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_5 vdd vdd vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_6 dummy_bl dummy_br vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_6 vdd vdd vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_7 dummy_bl dummy_br vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_7 vdd vdd vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_8 dummy_bl dummy_br vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_8 vdd vdd vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_9 dummy_bl dummy_br vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_9 vdd vdd vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_10 dummy_bl dummy_br vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_10 vdd vdd vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_11 dummy_bl dummy_br vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_11 vdd vdd vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_12 dummy_bl dummy_br vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_12 vdd vdd vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_13 dummy_bl dummy_br vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_13 vdd vdd vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_14 dummy_bl dummy_br vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_14 vdd vdd vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_15 dummy_bl dummy_br vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_15 vdd vdd vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_16 dummy_bl dummy_br vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_16 vdd vdd vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_17 dummy_bl dummy_br vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_17 vdd vdd vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_18 dummy_bl dummy_br vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_18 vdd vdd vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_19 dummy_bl dummy_br vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_19 vdd vdd vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_20 dummy_bl dummy_br vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_20 vdd vdd vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_21 dummy_bl dummy_br vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_21 vdd vdd vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_22 dummy_bl dummy_br vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_22 vdd vdd vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_23 dummy_bl dummy_br vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_23 vdd vdd vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_24 dummy_bl dummy_br vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_24 vdd vdd vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_25 dummy_bl dummy_br vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_25 vdd vdd vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_26 dummy_bl dummy_br vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_26 vdd vdd vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_27 dummy_bl dummy_br vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_27 vdd vdd vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_28 dummy_bl dummy_br vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_28 vdd vdd vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_29 dummy_bl dummy_br vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_29 vdd vdd vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_30 dummy_bl dummy_br vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_30 vdd vdd vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_31 dummy_bl dummy_br vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_31 vdd vdd vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_32 dummy_bl dummy_br vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_32 vdd vdd vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_33 dummy_bl dummy_br vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_33 vdd vdd vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_34 dummy_bl dummy_br vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_34 vdd vdd vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_35 dummy_bl dummy_br vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_35 vdd vdd vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_36 dummy_bl dummy_br vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_36 vdd vdd vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_37 dummy_bl dummy_br vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_37 vdd vdd vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_38 dummy_bl dummy_br vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_38 vdd vdd vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_39 dummy_bl dummy_br vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_39 vdd vdd vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_40 dummy_bl dummy_br vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_40 vdd vdd vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_41 dummy_bl dummy_br vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_41 vdd vdd vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_42 dummy_bl dummy_br vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_42 vdd vdd vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_43 dummy_bl dummy_br vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_43 vdd vdd vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_44 dummy_bl dummy_br vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_44 vdd vdd vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_45 dummy_bl dummy_br vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_45 vdd vdd vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_46 dummy_bl dummy_br vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_46 vdd vdd vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_47 dummy_bl dummy_br vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_47 vdd vdd vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_48 dummy_bl dummy_br vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_48 vdd vdd vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_49 dummy_bl dummy_br vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_49 vdd vdd vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_50 dummy_bl dummy_br vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_50 vdd vdd vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_51 dummy_bl dummy_br vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_51 vdd vdd vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_52 dummy_bl dummy_br vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_52 vdd vdd vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_53 dummy_bl dummy_br vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_53 vdd vdd vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_54 dummy_bl dummy_br vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_54 vdd vdd vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_55 dummy_bl dummy_br vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_55 vdd vdd vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_56 dummy_bl dummy_br vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_56 vdd vdd vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_57 dummy_bl dummy_br vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_57 vdd vdd vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_58 dummy_bl dummy_br vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_58 vdd vdd vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_59 dummy_bl dummy_br vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_59 vdd vdd vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_60 dummy_bl dummy_br vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_60 vdd vdd vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_61 dummy_bl dummy_br vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_61 vdd vdd vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_62 dummy_bl dummy_br vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_62 vdd vdd vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_63 dummy_bl dummy_br vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_63 vdd vdd vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_64 dummy_bl dummy_br vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_64 vdd vdd vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_65 dummy_bl dummy_br vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_65 vdd vdd vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_66 dummy_bl dummy_br vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_66 vdd vdd vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_67 dummy_bl dummy_br vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_67 vdd vdd vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_68 dummy_bl dummy_br vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_68 vdd vdd vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_69 dummy_bl dummy_br vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_69 vdd vdd vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_70 dummy_bl dummy_br vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_70 vdd vdd vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_71 dummy_bl dummy_br vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_71 vdd vdd vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_72 dummy_bl dummy_br vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_72 vdd vdd vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_73 dummy_bl dummy_br vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_73 vdd vdd vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_74 dummy_bl dummy_br vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_74 vdd vdd vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_75 dummy_bl dummy_br vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_75 vdd vdd vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_76 dummy_bl dummy_br vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_76 vdd vdd vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_77 dummy_bl dummy_br vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_77 vdd vdd vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_78 dummy_bl dummy_br vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_78 vdd vdd vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_79 dummy_bl dummy_br vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_79 vdd vdd vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_80 dummy_bl dummy_br vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_80 vdd vdd vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_81 dummy_bl dummy_br vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_81 vdd vdd vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_82 dummy_bl dummy_br vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_82 vdd vdd vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_83 dummy_bl dummy_br vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_83 vdd vdd vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_84 dummy_bl dummy_br vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_84 vdd vdd vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_85 dummy_bl dummy_br vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_85 vdd vdd vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_86 dummy_bl dummy_br vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_86 vdd vdd vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_87 dummy_bl dummy_br vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_87 vdd vdd vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_88 dummy_bl dummy_br vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_88 vdd vdd vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_89 dummy_bl dummy_br vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_89 vdd vdd vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_90 dummy_bl dummy_br vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_90 vdd vdd vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_91 dummy_bl dummy_br vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_91 vdd vdd vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_92 dummy_bl dummy_br vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_92 vdd vdd vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_93 dummy_bl dummy_br vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_93 vdd vdd vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_94 dummy_bl dummy_br vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_94 vdd vdd vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_95 dummy_bl dummy_br vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_95 vdd vdd vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_96 dummy_bl dummy_br vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_96 vdd vdd vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_97 dummy_bl dummy_br vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_97 vdd vdd vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_98 dummy_bl dummy_br vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_98 vdd vdd vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_99 dummy_bl dummy_br vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_99 vdd vdd vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_100 dummy_bl dummy_br vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_100 vdd vdd vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_101 dummy_bl dummy_br vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_101 vdd vdd vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_102 dummy_bl dummy_br vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_102 vdd vdd vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_103 dummy_bl dummy_br vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_103 vdd vdd vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_104 dummy_bl dummy_br vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_104 vdd vdd vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_105 dummy_bl dummy_br vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_105 vdd vdd vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_106 dummy_bl dummy_br vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_106 vdd vdd vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_107 dummy_bl dummy_br vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_107 vdd vdd vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_108 dummy_bl dummy_br vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_108 vdd vdd vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_109 dummy_bl dummy_br vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_109 vdd vdd vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_110 dummy_bl dummy_br vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_110 vdd vdd vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_111 dummy_bl dummy_br vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_111 vdd vdd vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_112 dummy_bl dummy_br vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_112 vdd vdd vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_113 dummy_bl dummy_br vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_113 vdd vdd vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_114 dummy_bl dummy_br vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_114 vdd vdd vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_115 dummy_bl dummy_br vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_115 vdd vdd vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_116 dummy_bl dummy_br vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_116 vdd vdd vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_117 dummy_bl dummy_br vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_117 vdd vdd vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_118 dummy_bl dummy_br vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_118 vdd vdd vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_119 dummy_bl dummy_br vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_119 vdd vdd vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_120 dummy_bl dummy_br vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_120 vdd vdd vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_121 dummy_bl dummy_br vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_121 vdd vdd vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_122 dummy_bl dummy_br vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_122 vdd vdd vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_123 dummy_bl dummy_br vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_123 vdd vdd vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_124 dummy_bl dummy_br vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_124 vdd vdd vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_125 dummy_bl dummy_br vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_125 vdd vdd vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_126 dummy_bl dummy_br vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_126 vdd vdd vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_127 dummy_bl dummy_br vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_127 vdd vdd vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_128 dummy_bl dummy_br vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_128 vdd vdd vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_129 dummy_bl dummy_br vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_129 vdd vdd vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_0 bl[0] br[0] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_0 bl[0] br[0] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_1 bl[1] br[1] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_1 bl[1] br[1] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_2 bl[2] br[2] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_2 bl[2] br[2] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_3 bl[3] br[3] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_3 bl[3] br[3] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_4 bl[4] br[4] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_4 bl[4] br[4] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_5 bl[5] br[5] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_5 bl[5] br[5] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_6 bl[6] br[6] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_6 bl[6] br[6] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_7 bl[7] br[7] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_7 bl[7] br[7] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_8 bl[8] br[8] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_8 bl[8] br[8] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_9 bl[9] br[9] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_9 bl[9] br[9] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_10 bl[10] br[10] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_10 bl[10] br[10] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_11 bl[11] br[11] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_11 bl[11] br[11] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_12 bl[12] br[12] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_12 bl[12] br[12] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_13 bl[13] br[13] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_13 bl[13] br[13] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_14 bl[14] br[14] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_14 bl[14] br[14] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_15 bl[15] br[15] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_15 bl[15] br[15] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_16 bl[16] br[16] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_16 bl[16] br[16] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_17 bl[17] br[17] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_17 bl[17] br[17] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_18 bl[18] br[18] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_18 bl[18] br[18] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_19 bl[19] br[19] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_19 bl[19] br[19] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_20 bl[20] br[20] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_20 bl[20] br[20] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_21 bl[21] br[21] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_21 bl[21] br[21] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_22 bl[22] br[22] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_22 bl[22] br[22] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_23 bl[23] br[23] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_23 bl[23] br[23] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_24 bl[24] br[24] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_24 bl[24] br[24] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_25 bl[25] br[25] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_25 bl[25] br[25] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_26 bl[26] br[26] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_26 bl[26] br[26] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_27 bl[27] br[27] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_27 bl[27] br[27] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_28 bl[28] br[28] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_28 bl[28] br[28] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_29 bl[29] br[29] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_29 bl[29] br[29] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_30 bl[30] br[30] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_30 bl[30] br[30] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_31 bl[31] br[31] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_31 bl[31] br[31] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_32 bl[32] br[32] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_32 bl[32] br[32] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_33 bl[33] br[33] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_33 bl[33] br[33] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_34 bl[34] br[34] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_34 bl[34] br[34] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_35 bl[35] br[35] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_35 bl[35] br[35] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_36 bl[36] br[36] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_36 bl[36] br[36] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_37 bl[37] br[37] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_37 bl[37] br[37] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_38 bl[38] br[38] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_38 bl[38] br[38] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_39 bl[39] br[39] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_39 bl[39] br[39] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_40 bl[40] br[40] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_40 bl[40] br[40] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_41 bl[41] br[41] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_41 bl[41] br[41] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_42 bl[42] br[42] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_42 bl[42] br[42] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_43 bl[43] br[43] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_43 bl[43] br[43] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_44 bl[44] br[44] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_44 bl[44] br[44] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_45 bl[45] br[45] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_45 bl[45] br[45] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_46 bl[46] br[46] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_46 bl[46] br[46] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_47 bl[47] br[47] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_47 bl[47] br[47] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_48 bl[48] br[48] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_48 bl[48] br[48] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_49 bl[49] br[49] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_49 bl[49] br[49] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_50 bl[50] br[50] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_50 bl[50] br[50] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_51 bl[51] br[51] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_51 bl[51] br[51] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_52 bl[52] br[52] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_52 bl[52] br[52] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_53 bl[53] br[53] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_53 bl[53] br[53] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_54 bl[54] br[54] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_54 bl[54] br[54] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_55 bl[55] br[55] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_55 bl[55] br[55] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_56 bl[56] br[56] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_56 bl[56] br[56] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_57 bl[57] br[57] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_57 bl[57] br[57] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_58 bl[58] br[58] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_58 bl[58] br[58] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_59 bl[59] br[59] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_59 bl[59] br[59] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_60 bl[60] br[60] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_60 bl[60] br[60] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_61 bl[61] br[61] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_61 bl[61] br[61] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_62 bl[62] br[62] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_62 bl[62] br[62] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_63 bl[63] br[63] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_63 bl[63] br[63] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xcolend_top_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_colend_wrapper
  Xcolend_bot_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_colend_wrapper
  Xhstrap_0_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_1 br[0] vdd vss bl[0] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_1 br[0] vdd vss bl[0] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_2 br[1] vdd vss bl[1] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_2 br[1] vdd vss bl[1] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_3 br[2] vdd vss bl[2] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_3 br[2] vdd vss bl[2] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_4 br[3] vdd vss bl[3] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_4 br[3] vdd vss bl[3] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_5 br[4] vdd vss bl[4] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_5 br[4] vdd vss bl[4] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_6 br[5] vdd vss bl[5] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_6 br[5] vdd vss bl[5] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_7 br[6] vdd vss bl[6] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_7 br[6] vdd vss bl[6] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_8 br[7] vdd vss bl[7] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_8 br[7] vdd vss bl[7] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_9 br[8] vdd vss bl[8] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_9 br[8] vdd vss bl[8] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_10 br[9] vdd vss bl[9] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_10 br[9] vdd vss bl[9] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_11 br[10] vdd vss bl[10] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_11 br[10] vdd vss bl[10] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_12 br[11] vdd vss bl[11] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_12 br[11] vdd vss bl[11] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_13 br[12] vdd vss bl[12] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_13 br[12] vdd vss bl[12] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_14 br[13] vdd vss bl[13] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_14 br[13] vdd vss bl[13] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_15 br[14] vdd vss bl[14] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_15 br[14] vdd vss bl[14] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_16 br[15] vdd vss bl[15] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_16 br[15] vdd vss bl[15] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_17 br[16] vdd vss bl[16] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_17 br[16] vdd vss bl[16] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_18 br[17] vdd vss bl[17] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_18 br[17] vdd vss bl[17] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_19 br[18] vdd vss bl[18] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_19 br[18] vdd vss bl[18] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_20 br[19] vdd vss bl[19] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_20 br[19] vdd vss bl[19] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_21 br[20] vdd vss bl[20] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_21 br[20] vdd vss bl[20] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_22 br[21] vdd vss bl[21] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_22 br[21] vdd vss bl[21] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_23 br[22] vdd vss bl[22] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_23 br[22] vdd vss bl[22] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_24 br[23] vdd vss bl[23] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_24 br[23] vdd vss bl[23] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_25 br[24] vdd vss bl[24] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_25 br[24] vdd vss bl[24] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_26 br[25] vdd vss bl[25] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_26 br[25] vdd vss bl[25] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_27 br[26] vdd vss bl[26] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_27 br[26] vdd vss bl[26] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_28 br[27] vdd vss bl[27] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_28 br[27] vdd vss bl[27] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_29 br[28] vdd vss bl[28] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_29 br[28] vdd vss bl[28] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_30 br[29] vdd vss bl[29] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_30 br[29] vdd vss bl[29] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_31 br[30] vdd vss bl[30] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_31 br[30] vdd vss bl[30] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_32 br[31] vdd vss bl[31] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_32 br[31] vdd vss bl[31] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_33 br[32] vdd vss bl[32] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_33 br[32] vdd vss bl[32] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_34 br[33] vdd vss bl[33] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_34 br[33] vdd vss bl[33] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_35 br[34] vdd vss bl[34] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_35 br[34] vdd vss bl[34] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_36 br[35] vdd vss bl[35] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_36 br[35] vdd vss bl[35] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_37 br[36] vdd vss bl[36] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_37 br[36] vdd vss bl[36] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_38 br[37] vdd vss bl[37] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_38 br[37] vdd vss bl[37] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_39 br[38] vdd vss bl[38] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_39 br[38] vdd vss bl[38] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_40 br[39] vdd vss bl[39] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_40 br[39] vdd vss bl[39] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_41 br[40] vdd vss bl[40] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_41 br[40] vdd vss bl[40] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_42 br[41] vdd vss bl[41] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_42 br[41] vdd vss bl[41] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_43 br[42] vdd vss bl[42] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_43 br[42] vdd vss bl[42] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_44 br[43] vdd vss bl[43] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_44 br[43] vdd vss bl[43] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_45 br[44] vdd vss bl[44] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_45 br[44] vdd vss bl[44] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_46 br[45] vdd vss bl[45] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_46 br[45] vdd vss bl[45] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_47 br[46] vdd vss bl[46] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_47 br[46] vdd vss bl[46] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_48 br[47] vdd vss bl[47] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_48 br[47] vdd vss bl[47] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_49 br[48] vdd vss bl[48] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_49 br[48] vdd vss bl[48] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_50 br[49] vdd vss bl[49] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_50 br[49] vdd vss bl[49] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_51 br[50] vdd vss bl[50] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_51 br[50] vdd vss bl[50] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_52 br[51] vdd vss bl[51] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_52 br[51] vdd vss bl[51] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_53 br[52] vdd vss bl[52] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_53 br[52] vdd vss bl[52] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_54 br[53] vdd vss bl[53] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_54 br[53] vdd vss bl[53] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_55 br[54] vdd vss bl[54] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_55 br[54] vdd vss bl[54] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_56 br[55] vdd vss bl[55] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_56 br[55] vdd vss bl[55] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_57 br[56] vdd vss bl[56] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_57 br[56] vdd vss bl[56] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_58 br[57] vdd vss bl[57] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_58 br[57] vdd vss bl[57] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_59 br[58] vdd vss bl[58] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_59 br[58] vdd vss bl[58] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_60 br[59] vdd vss bl[59] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_60 br[59] vdd vss bl[59] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_61 br[60] vdd vss bl[60] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_61 br[60] vdd vss bl[60] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_62 br[61] vdd vss bl[61] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_62 br[61] vdd vss bl[61] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_63 br[62] vdd vss bl[62] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_63 br[62] vdd vss bl[62] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_64 br[63] vdd vss bl[63] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_64 br[63] vdd vss bl[63] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_65 vdd vdd vss vdd vss vdd sram_sp_colend_wrapper
  Xcolend_bot_65 vdd vdd vss vdd vss vdd sram_sp_colend_wrapper
  Xhstrap_0_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhoriz_wlstrap_0_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper

.ENDS sp_cell_array

.SUBCKT sram_sp_rowtapend_replica VSS VNB

  X0 VSS VSS VSS VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.420


.ENDS sram_sp_rowtapend_replica

.SUBCKT sram_sp_rowtapend_replica_wrapper VSS VNB

  X0 VSS VNB sram_sp_rowtapend_replica

.ENDS sram_sp_rowtapend_replica_wrapper

.SUBCKT replica_cell_array vdd vss rbl rbr rwl

  Xcell_0_0 rbl rbr vss vdd vdd vss rwl sram_sp_cell_replica_wrapper
  Xcell_0_1 rbl rbr vss vdd vdd vss rwl sram_sp_cell_replica_wrapper
  Xcell_1_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_1_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_2_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_2_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_3_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_3_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_4_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_4_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_5_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_5_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_6_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_6_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_7_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_7_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_8_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_8_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_9_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_9_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_10_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_10_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_11_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_11_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_12_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_12_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_13_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_13_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_14_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_14_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_15_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_15_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_16_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_16_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_17_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_17_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_18_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_18_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_19_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_19_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_20_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_20_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_21_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_21_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_22_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_22_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_23_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_23_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_24_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_24_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_25_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_25_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcolend_0_0 rbr vdd vss rbl vss vdd sram_sp_colend_wrapper
  Xcolend_1_0 rbr vdd vss rbl vss vdd sram_sp_colend_wrapper
  Xcolend_0_1 rbr vdd vss rbl vss vdd sram_sp_colend_wrapper
  Xcolend_1_1 rbr vdd vss rbl vss vdd sram_sp_colend_wrapper
  Xrowtapend_0_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_0_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_0_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_0_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xrowtapend_1_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_1_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_1_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xrowtapend_2_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_2_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_2_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xrowtapend_3_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_3_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_3_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xrowtapend_4_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_4_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_4_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xrowtapend_5_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_5_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_5_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xrowtapend_6_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_6_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_6_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper

.ENDS replica_cell_array

.SUBCKT dff_array_8 vdd vss clk rb d[0] d[1] d[2] d[3] d[4] d[5] d[6] d[7] q[0] q[1] q[2] q[3] q[4] q[5] q[6] q[7] qn[0] qn[1] qn[2] qn[3] qn[4] qn[5] qn[6] qn[7]

  Xdff_0 clk d[0] rb vss vss vdd vdd q[0] qn[0] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_1 clk d[1] rb vss vss vdd vdd q[1] qn[1] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_2 clk d[2] rb vss vss vdd vdd q[2] qn[2] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_3 clk d[3] rb vss vss vdd vdd q[3] qn[3] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_4 clk d[4] rb vss vss vdd vdd q[4] qn[4] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_5 clk d[5] rb vss vss vdd vdd q[5] qn[5] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_6 clk d[6] rb vss vss vdd vdd q[6] qn[6] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_7 clk d[7] rb vss vss vdd vdd q[7] qn[7] sky130_fd_sc_hs__dfrbp_2_wrapper

.ENDS dff_array_8

.SUBCKT mos_w3350_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=3.350


.ENDS mos_w3350_l150_m1_nf1_id1

.SUBCKT mos_w1350_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.350


.ENDS mos_w1350_l150_m1_nf1_id0

.SUBCKT folded_inv_3 vdd vss a y

  XMP0 y a vdd vdd mos_w3350_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w1350_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w3350_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w1350_l150_m1_nf1_id0

.ENDS folded_inv_3

.SUBCKT decoder_stage_7 vdd vss y y_b predecode_0_0 predecode_1_0

  Xgate_0_0_0 vdd vss predecode_0_0 predecode_1_0 x_0 nand2_1
  Xgate_1_0_0 vdd vss x_0 x_1 folded_inv_2
  Xgate_2_0_0 vdd vss x_1 y_b folded_inv_3
  Xgate_3_0_0 vdd vss y_b y folded_inv_3

.ENDS decoder_stage_7

.SUBCKT mos_w5000_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=5.000


.ENDS mos_w5000_l150_m1_nf1_id0

.SUBCKT tristate_inv din en en_b din_b vdd vss

  Xmn_en din_b en nint vss mos_w5000_l150_m1_nf1_id0
  Xmn_pd nint din vss vss mos_w5000_l150_m1_nf1_id0
  Xmp_en din_b en_b pint vdd mos_w5000_l150_m1_nf1_id1
  Xmp_pu pint din vdd vdd mos_w5000_l150_m1_nf1_id1

.ENDS tristate_inv

.SUBCKT write_driver en en_b data data_b bl br vdd vss

  Xbldriver data_b en en_b bl vdd vss tristate_inv
  Xbrdriver data en en_b br vdd vss tristate_inv

.ENDS write_driver

.SUBCKT sramgen_sp_sense_amp clk inn inp outn outp VDD VSS

  XSWOP outp clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=1.000

  XSWON outn clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=1.000

  XSWMP midp clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=1.000

  XSWMN midn clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=1.000

  XPFBP outp outn VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=2.000

  XPFBN outn outp VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=2.000

  XTAIL tail clk VSS VSS sky130_fd_pr__nfet_01v8 l=0.150 nf=4 w=1.680

  XNFBP outp outn midp VSS sky130_fd_pr__nfet_01v8 l=0.150 nf=2 w=1.680

  XNFBN outn outp midn VSS sky130_fd_pr__nfet_01v8 l=0.150 nf=2 w=1.680

  XINP midn inp tail VSS sky130_fd_pr__nfet_01v8 l=0.150 nf=2 w=1.680

  XINN midp inn tail VSS sky130_fd_pr__nfet_01v8 l=0.150 nf=2 w=1.680


.ENDS sramgen_sp_sense_amp

.SUBCKT sramgen_sp_sense_amp_wrapper clk inn inp outn outp VDD VSS

  X0 clk inn inp outn outp VDD VSS sramgen_sp_sense_amp

.ENDS sramgen_sp_sense_amp_wrapper

.SUBCKT mos_w1000_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000


.ENDS mos_w1000_l150_m1_nf1_id1

.SUBCKT folded_inv_7 vdd vss a y

  XMP0 y a vdd vdd mos_w1000_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w600_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w1000_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w600_l150_m1_nf1_id0

.ENDS folded_inv_7

.SUBCKT mos_w1000_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.000


.ENDS mos_w1000_l150_m1_nf1_id0

.SUBCKT diff_latch vdd vss din1 din2 dout1 dout2

  Xinbuf_1 vdd vss din1 rst folded_inv_7
  Xinbuf_2 vdd vss din2 set folded_inv_7
  Xoutbuf_1 vdd vss q dout2 folded_inv_7
  Xoutbuf_2 vdd vss qb dout1 folded_inv_7
  Xinvq_1 vdd vss q qb folded_inv_7
  Xinvq_2 vdd vss qb q folded_inv_7
  XMN10 q rst vss vss mos_w1000_l150_m1_nf1_id0
  XMN11 q rst vss vss mos_w1000_l150_m1_nf1_id0
  XMN20 qb set vss vss mos_w1000_l150_m1_nf1_id0
  XMN21 qb set vss vss mos_w1000_l150_m1_nf1_id0

.ENDS diff_latch

.SUBCKT column clk rstb vdd vss bl[0] bl[1] bl[2] bl[3] bl[4] bl[5] bl[6] bl[7] br[0] br[1] br[2] br[3] br[4] br[5] br[6] br[7] pc_b sel[0] sel[1] sel[2] sel[3] sel[4] sel[5] sel[6] sel[7] sel_b[0] sel_b[1] sel_b[2] sel_b[3] sel_b[4] sel_b[5] sel_b[6] sel_b[7] we we_b din dout sense_en

  Xprecharge_0 vdd bl[0] br[0] pc_b precharge_1
  Xmux_0 sel_b[0] sel[0] bl[0] br[0] bl_out br_out vdd vss tgate_mux
  Xprecharge_1 vdd bl[1] br[1] pc_b precharge_1
  Xmux_1 sel_b[1] sel[1] bl[1] br[1] bl_out br_out vdd vss tgate_mux
  Xprecharge_2 vdd bl[2] br[2] pc_b precharge_1
  Xmux_2 sel_b[2] sel[2] bl[2] br[2] bl_out br_out vdd vss tgate_mux
  Xprecharge_3 vdd bl[3] br[3] pc_b precharge_1
  Xmux_3 sel_b[3] sel[3] bl[3] br[3] bl_out br_out vdd vss tgate_mux
  Xprecharge_4 vdd bl[4] br[4] pc_b precharge_1
  Xmux_4 sel_b[4] sel[4] bl[4] br[4] bl_out br_out vdd vss tgate_mux
  Xprecharge_5 vdd bl[5] br[5] pc_b precharge_1
  Xmux_5 sel_b[5] sel[5] bl[5] br[5] bl_out br_out vdd vss tgate_mux
  Xprecharge_6 vdd bl[6] br[6] pc_b precharge_1
  Xmux_6 sel_b[6] sel[6] bl[6] br[6] bl_out br_out vdd vss tgate_mux
  Xprecharge_7 vdd bl[7] br[7] pc_b precharge_1
  Xmux_7 sel_b[7] sel[7] bl[7] br[7] bl_out br_out vdd vss tgate_mux
  Xwrite_driver we we_b q q_b bl_out br_out vdd vss write_driver
  Xsense_amp sense_en br_out bl_out sa_outn sa_outp vdd vss sramgen_sp_sense_amp_wrapper
  Xlatch vdd vss sa_outp sa_outn dout diff_latch_outn diff_latch
  Xdff clk din rstb vss vss vdd vdd q q_b sky130_fd_sc_hs__dfrbp_2_wrapper

.ENDS column

.SUBCKT col_peripherals clk rstb vdd vss sense_en bl[0] bl[1] bl[2] bl[3] bl[4] bl[5] bl[6] bl[7] bl[8] bl[9] bl[10] bl[11] bl[12] bl[13] bl[14] bl[15] bl[16] bl[17] bl[18] bl[19] bl[20] bl[21] bl[22] bl[23] bl[24] bl[25] bl[26] bl[27] bl[28] bl[29] bl[30] bl[31] bl[32] bl[33] bl[34] bl[35] bl[36] bl[37] bl[38] bl[39] bl[40] bl[41] bl[42] bl[43] bl[44] bl[45] bl[46] bl[47] bl[48] bl[49] bl[50] bl[51] bl[52] bl[53] bl[54] bl[55] bl[56] bl[57] bl[58] bl[59] bl[60] bl[61] bl[62] bl[63] br[0] br[1] br[2] br[3] br[4] br[5] br[6] br[7] br[8] br[9] br[10] br[11] br[12] br[13] br[14] br[15] br[16] br[17] br[18] br[19] br[20] br[21] br[22] br[23] br[24] br[25] br[26] br[27] br[28] br[29] br[30] br[31] br[32] br[33] br[34] br[35] br[36] br[37] br[38] br[39] br[40] br[41] br[42] br[43] br[44] br[45] br[46] br[47] br[48] br[49] br[50] br[51] br[52] br[53] br[54] br[55] br[56] br[57] br[58] br[59] br[60] br[61] br[62] br[63] pc_b sel[0] sel[1] sel[2] sel[3] sel[4] sel[5] sel[6] sel[7] sel_b[0] sel_b[1] sel_b[2] sel_b[3] sel_b[4] sel_b[5] sel_b[6] sel_b[7] we wmask[0] wmask[1] wmask[2] wmask[3] wmask[4] wmask[5] wmask[6] wmask[7] din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] dout[0] dout[1] dout[2] dout[3] dout[4] dout[5] dout[6] dout[7]

  Xwmask_dffs vdd vss clk rstb wmask[0] wmask[1] wmask[2] wmask[3] wmask[4] wmask[5] wmask[6] wmask[7] wmask_in[0] wmask_in[1] wmask_in[2] wmask_in[3] wmask_in[4] wmask_in[5] wmask_in[6] wmask_in[7] wmask_in_b[0] wmask_in_b[1] wmask_in_b[2] wmask_in_b[3] wmask_in_b[4] wmask_in_b[5] wmask_in_b[6] wmask_in_b[7] dff_array_8
  Xwmask_and_0 vdd vss we_i[0] we_ib[0] we wmask_in[0] decoder_stage_7
  Xwmask_and_1 vdd vss we_i[1] we_ib[1] we wmask_in[1] decoder_stage_7
  Xwmask_and_2 vdd vss we_i[2] we_ib[2] we wmask_in[2] decoder_stage_7
  Xwmask_and_3 vdd vss we_i[3] we_ib[3] we wmask_in[3] decoder_stage_7
  Xwmask_and_4 vdd vss we_i[4] we_ib[4] we wmask_in[4] decoder_stage_7
  Xwmask_and_5 vdd vss we_i[5] we_ib[5] we wmask_in[5] decoder_stage_7
  Xwmask_and_6 vdd vss we_i[6] we_ib[6] we wmask_in[6] decoder_stage_7
  Xwmask_and_7 vdd vss we_i[7] we_ib[7] we wmask_in[7] decoder_stage_7
  Xcol_group_0 clk rstb vdd vss bl[0] bl[1] bl[2] bl[3] bl[4] bl[5] bl[6] bl[7] br[0] br[1] br[2] br[3] br[4] br[5] br[6] br[7] pc_b sel[0] sel[1] sel[2] sel[3] sel[4] sel[5] sel[6] sel[7] sel_b[0] sel_b[1] sel_b[2] sel_b[3] sel_b[4] sel_b[5] sel_b[6] sel_b[7] we_i[0] we_ib[0] din[0] dout[0] sense_en column
  Xcol_group_1 clk rstb vdd vss bl[8] bl[9] bl[10] bl[11] bl[12] bl[13] bl[14] bl[15] br[8] br[9] br[10] br[11] br[12] br[13] br[14] br[15] pc_b sel[0] sel[1] sel[2] sel[3] sel[4] sel[5] sel[6] sel[7] sel_b[0] sel_b[1] sel_b[2] sel_b[3] sel_b[4] sel_b[5] sel_b[6] sel_b[7] we_i[1] we_ib[1] din[1] dout[1] sense_en column
  Xcol_group_2 clk rstb vdd vss bl[16] bl[17] bl[18] bl[19] bl[20] bl[21] bl[22] bl[23] br[16] br[17] br[18] br[19] br[20] br[21] br[22] br[23] pc_b sel[0] sel[1] sel[2] sel[3] sel[4] sel[5] sel[6] sel[7] sel_b[0] sel_b[1] sel_b[2] sel_b[3] sel_b[4] sel_b[5] sel_b[6] sel_b[7] we_i[2] we_ib[2] din[2] dout[2] sense_en column
  Xcol_group_3 clk rstb vdd vss bl[24] bl[25] bl[26] bl[27] bl[28] bl[29] bl[30] bl[31] br[24] br[25] br[26] br[27] br[28] br[29] br[30] br[31] pc_b sel[0] sel[1] sel[2] sel[3] sel[4] sel[5] sel[6] sel[7] sel_b[0] sel_b[1] sel_b[2] sel_b[3] sel_b[4] sel_b[5] sel_b[6] sel_b[7] we_i[3] we_ib[3] din[3] dout[3] sense_en column
  Xcol_group_4 clk rstb vdd vss bl[32] bl[33] bl[34] bl[35] bl[36] bl[37] bl[38] bl[39] br[32] br[33] br[34] br[35] br[36] br[37] br[38] br[39] pc_b sel[0] sel[1] sel[2] sel[3] sel[4] sel[5] sel[6] sel[7] sel_b[0] sel_b[1] sel_b[2] sel_b[3] sel_b[4] sel_b[5] sel_b[6] sel_b[7] we_i[4] we_ib[4] din[4] dout[4] sense_en column
  Xcol_group_5 clk rstb vdd vss bl[40] bl[41] bl[42] bl[43] bl[44] bl[45] bl[46] bl[47] br[40] br[41] br[42] br[43] br[44] br[45] br[46] br[47] pc_b sel[0] sel[1] sel[2] sel[3] sel[4] sel[5] sel[6] sel[7] sel_b[0] sel_b[1] sel_b[2] sel_b[3] sel_b[4] sel_b[5] sel_b[6] sel_b[7] we_i[5] we_ib[5] din[5] dout[5] sense_en column
  Xcol_group_6 clk rstb vdd vss bl[48] bl[49] bl[50] bl[51] bl[52] bl[53] bl[54] bl[55] br[48] br[49] br[50] br[51] br[52] br[53] br[54] br[55] pc_b sel[0] sel[1] sel[2] sel[3] sel[4] sel[5] sel[6] sel[7] sel_b[0] sel_b[1] sel_b[2] sel_b[3] sel_b[4] sel_b[5] sel_b[6] sel_b[7] we_i[6] we_ib[6] din[6] dout[6] sense_en column
  Xcol_group_7 clk rstb vdd vss bl[56] bl[57] bl[58] bl[59] bl[60] bl[61] bl[62] bl[63] br[56] br[57] br[58] br[59] br[60] br[61] br[62] br[63] pc_b sel[0] sel[1] sel[2] sel[3] sel[4] sel[5] sel[6] sel[7] sel_b[0] sel_b[1] sel_b[2] sel_b[3] sel_b[4] sel_b[5] sel_b[6] sel_b[7] we_i[7] we_ib[7] din[7] dout[7] sense_en column

.ENDS col_peripherals

.SUBCKT mos_w850_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.850


.ENDS mos_w850_l150_m1_nf1_id1

.SUBCKT mos_w500_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.500


.ENDS mos_w500_l150_m1_nf1_id1

.SUBCKT precharge vdd bl br en_b

  Xbl_pull_up bl en_b vdd vdd mos_w850_l150_m1_nf1_id1
  Xbr_pull_up br en_b vdd vdd mos_w850_l150_m1_nf1_id1
  Xequalizer bl en_b br vdd mos_w500_l150_m1_nf1_id1

.ENDS precharge

.SUBCKT sram22_inner vdd vss clk we ce rstb addr[0] addr[1] addr[2] addr[3] addr[4] addr[5] addr[6] addr[7] addr[8] addr[9] wmask[0] wmask[1] wmask[2] wmask[3] wmask[4] wmask[5] wmask[6] wmask[7] din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] dout[0] dout[1] dout[2] dout[3] dout[4] dout[5] dout[6] dout[7]

  Xaddr_gate vdd vss addr_gated[0] addr_gated[1] addr_gated[2] addr_gated[3] addr_gated[4] addr_gated[5] addr_gated[6] addr_b_gated[0] addr_b_gated[1] addr_b_gated[2] addr_b_gated[3] addr_b_gated[4] addr_b_gated[5] addr_b_gated[6] addr_gate_y_b_noconn[0] addr_gate_y_b_noconn[1] addr_gate_y_b_noconn[2] addr_gate_y_b_noconn[3] addr_gate_y_b_noconn[4] addr_gate_y_b_noconn[5] addr_gate_y_b_noconn[6] addr_gate_y_b_noconn[7] addr_gate_y_b_noconn[8] addr_gate_y_b_noconn[9] addr_gate_y_b_noconn[10] addr_gate_y_b_noconn[11] addr_gate_y_b_noconn[12] addr_gate_y_b_noconn[13] wl_en addr_in[3] addr_in[4] addr_in[5] addr_in[6] addr_in[7] addr_in[8] addr_in[9] addr_in_b[3] addr_in_b[4] addr_in_b[5] addr_in_b[6] addr_in_b[7] addr_in_b[8] addr_in_b[9] decoder_stage
  Xdecoder vdd vss wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] wl_b[0] wl_b[1] wl_b[2] wl_b[3] wl_b[4] wl_b[5] wl_b[6] wl_b[7] wl_b[8] wl_b[9] wl_b[10] wl_b[11] wl_b[12] wl_b[13] wl_b[14] wl_b[15] wl_b[16] wl_b[17] wl_b[18] wl_b[19] wl_b[20] wl_b[21] wl_b[22] wl_b[23] wl_b[24] wl_b[25] wl_b[26] wl_b[27] wl_b[28] wl_b[29] wl_b[30] wl_b[31] wl_b[32] wl_b[33] wl_b[34] wl_b[35] wl_b[36] wl_b[37] wl_b[38] wl_b[39] wl_b[40] wl_b[41] wl_b[42] wl_b[43] wl_b[44] wl_b[45] wl_b[46] wl_b[47] wl_b[48] wl_b[49] wl_b[50] wl_b[51] wl_b[52] wl_b[53] wl_b[54] wl_b[55] wl_b[56] wl_b[57] wl_b[58] wl_b[59] wl_b[60] wl_b[61] wl_b[62] wl_b[63] wl_b[64] wl_b[65] wl_b[66] wl_b[67] wl_b[68] wl_b[69] wl_b[70] wl_b[71] wl_b[72] wl_b[73] wl_b[74] wl_b[75] wl_b[76] wl_b[77] wl_b[78] wl_b[79] wl_b[80] wl_b[81] wl_b[82] wl_b[83] wl_b[84] wl_b[85] wl_b[86] wl_b[87] wl_b[88] wl_b[89] wl_b[90] wl_b[91] wl_b[92] wl_b[93] wl_b[94] wl_b[95] wl_b[96] wl_b[97] wl_b[98] wl_b[99] wl_b[100] wl_b[101] wl_b[102] wl_b[103] wl_b[104] wl_b[105] wl_b[106] wl_b[107] wl_b[108] wl_b[109] wl_b[110] wl_b[111] wl_b[112] wl_b[113] wl_b[114] wl_b[115] wl_b[116] wl_b[117] wl_b[118] wl_b[119] wl_b[120] wl_b[121] wl_b[122] wl_b[123] wl_b[124] wl_b[125] wl_b[126] wl_b[127] addr_b_gated[0] addr_gated[0] addr_b_gated[1] addr_gated[1] addr_b_gated[2] addr_gated[2] addr_b_gated[3] addr_gated[3] addr_b_gated[4] addr_gated[4] addr_b_gated[5] addr_gated[5] addr_b_gated[6] addr_gated[6] decoder
  Xcolumn_decoder vdd vss col_sel[0] col_sel[1] col_sel[2] col_sel[3] col_sel[4] col_sel[5] col_sel[6] col_sel[7] col_sel_b[0] col_sel_b[1] col_sel_b[2] col_sel_b[3] col_sel_b[4] col_sel_b[5] col_sel_b[6] col_sel_b[7] addr_in_b[0] addr_in[0] addr_in_b[1] addr_in[1] addr_in_b[2] addr_in[2] decoder_1
  Xcontrol_logic clk ce_in we_in rstb rbl sense_en0 pc_b0 rwl wl_en0 write_driver_en0 vdd vss control_logic_replica_v2
  Xpc_b_buffer vdd vss pc_b pc pc_b0 decoder_stage_1
  Xwlen_buffer vdd vss wl_en wl_en_b wl_en0 decoder_stage_2
  Xwrite_driver_en_buffer vdd vss write_driver_en write_driver_en_b write_driver_en0 decoder_stage_3
  Xsense_en_buffer vdd vss sense_en sense_en_b sense_en0 decoder_stage_4
  Xaddr_we_ce_dffs vdd vss clk rstb addr[0] addr[1] addr[2] addr[3] addr[4] addr[5] addr[6] addr[7] addr[8] addr[9] we ce addr_in[0] addr_in[1] addr_in[2] addr_in[3] addr_in[4] addr_in[5] addr_in[6] addr_in[7] addr_in[8] addr_in[9] we_in ce_in addr_in_b[0] addr_in_b[1] addr_in_b[2] addr_in_b[3] addr_in_b[4] addr_in_b[5] addr_in_b[6] addr_in_b[7] addr_in_b[8] addr_in_b[9] we_in_b ce_in_b dff_array_12
  Xbitcell_array vdd vss vdd vdd bl[0] bl[1] bl[2] bl[3] bl[4] bl[5] bl[6] bl[7] bl[8] bl[9] bl[10] bl[11] bl[12] bl[13] bl[14] bl[15] bl[16] bl[17] bl[18] bl[19] bl[20] bl[21] bl[22] bl[23] bl[24] bl[25] bl[26] bl[27] bl[28] bl[29] bl[30] bl[31] bl[32] bl[33] bl[34] bl[35] bl[36] bl[37] bl[38] bl[39] bl[40] bl[41] bl[42] bl[43] bl[44] bl[45] bl[46] bl[47] bl[48] bl[49] bl[50] bl[51] bl[52] bl[53] bl[54] bl[55] bl[56] bl[57] bl[58] bl[59] bl[60] bl[61] bl[62] bl[63] br[0] br[1] br[2] br[3] br[4] br[5] br[6] br[7] br[8] br[9] br[10] br[11] br[12] br[13] br[14] br[15] br[16] br[17] br[18] br[19] br[20] br[21] br[22] br[23] br[24] br[25] br[26] br[27] br[28] br[29] br[30] br[31] br[32] br[33] br[34] br[35] br[36] br[37] br[38] br[39] br[40] br[41] br[42] br[43] br[44] br[45] br[46] br[47] br[48] br[49] br[50] br[51] br[52] br[53] br[54] br[55] br[56] br[57] br[58] br[59] br[60] br[61] br[62] br[63] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] sp_cell_array
  Xreplica_bitcell_array vdd vss rbl rbr rwl replica_cell_array
  Xcol_circuitry clk rstb vdd vss sense_en bl[0] bl[1] bl[2] bl[3] bl[4] bl[5] bl[6] bl[7] bl[8] bl[9] bl[10] bl[11] bl[12] bl[13] bl[14] bl[15] bl[16] bl[17] bl[18] bl[19] bl[20] bl[21] bl[22] bl[23] bl[24] bl[25] bl[26] bl[27] bl[28] bl[29] bl[30] bl[31] bl[32] bl[33] bl[34] bl[35] bl[36] bl[37] bl[38] bl[39] bl[40] bl[41] bl[42] bl[43] bl[44] bl[45] bl[46] bl[47] bl[48] bl[49] bl[50] bl[51] bl[52] bl[53] bl[54] bl[55] bl[56] bl[57] bl[58] bl[59] bl[60] bl[61] bl[62] bl[63] br[0] br[1] br[2] br[3] br[4] br[5] br[6] br[7] br[8] br[9] br[10] br[11] br[12] br[13] br[14] br[15] br[16] br[17] br[18] br[19] br[20] br[21] br[22] br[23] br[24] br[25] br[26] br[27] br[28] br[29] br[30] br[31] br[32] br[33] br[34] br[35] br[36] br[37] br[38] br[39] br[40] br[41] br[42] br[43] br[44] br[45] br[46] br[47] br[48] br[49] br[50] br[51] br[52] br[53] br[54] br[55] br[56] br[57] br[58] br[59] br[60] br[61] br[62] br[63] pc_b col_sel[0] col_sel[1] col_sel[2] col_sel[3] col_sel[4] col_sel[5] col_sel[6] col_sel[7] col_sel_b[0] col_sel_b[1] col_sel_b[2] col_sel_b[3] col_sel_b[4] col_sel_b[5] col_sel_b[6] col_sel_b[7] write_driver_en wmask[0] wmask[1] wmask[2] wmask[3] wmask[4] wmask[5] wmask[6] wmask[7] din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] dout[0] dout[1] dout[2] dout[3] dout[4] dout[5] dout[6] dout[7] col_peripherals
  Xreplica_precharge_0 vdd rbl rbr pc_b0 precharge
  Xreplica_precharge_1 vdd rbl rbr pc_b0 precharge
  Xreplica_mos vdd vss rbl replica_column_mos

.ENDS sram22_inner

.SUBCKT sram22_1024x8m8w1 vdd vss clk we ce rstb addr[0] addr[1] addr[2] addr[3] addr[4] addr[5] addr[6] addr[7] addr[8] addr[9] wmask[0] wmask[1] wmask[2] wmask[3] wmask[4] wmask[5] wmask[6] wmask[7] din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] dout[0] dout[1] dout[2] dout[3] dout[4] dout[5] dout[6] dout[7]

  X0 vdd vss clk we ce rstb addr[0] addr[1] addr[2] addr[3] addr[4] addr[5] addr[6] addr[7] addr[8] addr[9] wmask[0] wmask[1] wmask[2] wmask[3] wmask[4] wmask[5] wmask[6] wmask[7] din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] dout[0] dout[1] dout[2] dout[3] dout[4] dout[5] dout[6] dout[7] sram22_inner

.ENDS sram22_1024x8m8w1

