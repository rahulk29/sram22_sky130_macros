VERSION 5.8 ; 
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 
MACRO sram22_512x8m8w1
    CLASS BLOCK  ;
    FOREIGN sram22_512x8m8w1   ;
    SIZE 270.560 BY 297.080 ;
    SYMMETRY X Y R90 ;
    PIN dout[0] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.432400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 172.830 0.000 172.970 0.140 ;
        END 
    END dout[0] 
    PIN dout[1] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.432400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 183.730 0.000 183.870 0.140 ;
        END 
    END dout[1] 
    PIN dout[2] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.432400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 194.630 0.000 194.770 0.140 ;
        END 
    END dout[2] 
    PIN dout[3] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.432400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 205.530 0.000 205.670 0.140 ;
        END 
    END dout[3] 
    PIN dout[4] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.432400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 216.430 0.000 216.570 0.140 ;
        END 
    END dout[4] 
    PIN dout[5] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.432400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 227.330 0.000 227.470 0.140 ;
        END 
    END dout[5] 
    PIN dout[6] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.432400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 238.230 0.000 238.370 0.140 ;
        END 
    END dout[6] 
    PIN dout[7] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.432400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 249.130 0.000 249.270 0.140 ;
        END 
    END dout[7] 
    PIN din[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.802100 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.154000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 172.410 0.000 172.550 0.140 ;
        END 
    END din[0] 
    PIN din[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.802100 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.154000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 183.310 0.000 183.450 0.140 ;
        END 
    END din[1] 
    PIN din[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.802100 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.154000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 194.210 0.000 194.350 0.140 ;
        END 
    END din[2] 
    PIN din[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.802100 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.154000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 205.110 0.000 205.250 0.140 ;
        END 
    END din[3] 
    PIN din[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.802100 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.154000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 216.010 0.000 216.150 0.140 ;
        END 
    END din[4] 
    PIN din[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.802100 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.154000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 226.910 0.000 227.050 0.140 ;
        END 
    END din[5] 
    PIN din[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.802100 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.154000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 237.810 0.000 237.950 0.140 ;
        END 
    END din[6] 
    PIN din[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.802100 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.154000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 248.710 0.000 248.850 0.140 ;
        END 
    END din[7] 
    PIN wmask[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.612500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 172.060 0.000 172.200 0.140 ;
        END 
    END wmask[0] 
    PIN wmask[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.612500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 182.960 0.000 183.100 0.140 ;
        END 
    END wmask[1] 
    PIN wmask[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.612500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 193.860 0.000 194.000 0.140 ;
        END 
    END wmask[2] 
    PIN wmask[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.612500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 204.760 0.000 204.900 0.140 ;
        END 
    END wmask[3] 
    PIN wmask[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.612500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 215.660 0.000 215.800 0.140 ;
        END 
    END wmask[4] 
    PIN wmask[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.612500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 226.560 0.000 226.700 0.140 ;
        END 
    END wmask[5] 
    PIN wmask[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.612500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 237.460 0.000 237.600 0.140 ;
        END 
    END wmask[6] 
    PIN wmask[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.612500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 248.360 0.000 248.500 0.140 ;
        END 
    END wmask[7] 
    PIN addr[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.011900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 116.760 0.000 117.080 0.320 ;
        END 
    END addr[0] 
    PIN addr[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.011900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 110.640 0.000 110.960 0.320 ;
        END 
    END addr[1] 
    PIN addr[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.011900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 104.520 0.000 104.840 0.320 ;
        END 
    END addr[2] 
    PIN addr[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.011900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 98.400 0.000 98.720 0.320 ;
        END 
    END addr[3] 
    PIN addr[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.011900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 92.960 0.000 93.280 0.320 ;
        END 
    END addr[4] 
    PIN addr[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.011900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 86.840 0.000 87.160 0.320 ;
        END 
    END addr[5] 
    PIN addr[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.011900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 80.720 0.000 81.040 0.320 ;
        END 
    END addr[6] 
    PIN addr[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.011900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 74.600 0.000 74.920 0.320 ;
        END 
    END addr[7] 
    PIN addr[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.011900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 68.480 0.000 68.800 0.320 ;
        END 
    END addr[8] 
    PIN we 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.011900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 129.000 0.000 129.320 0.320 ;
        END 
    END we 
    PIN ce 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.011900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 122.880 0.000 123.200 0.320 ;
        END 
    END ce 
    PIN clk 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 10.323000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 132.400 0.000 132.720 0.320 ;
        END 
    END clk 
    PIN rstb 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 14.229000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 133.080 0.000 133.400 0.320 ;
        END 
    END rstb 
    PIN vdd 
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT 
            LAYER met2 ;
                RECT 0.160 5.920 172.160 6.240 ;
                RECT 250.040 5.920 270.400 6.240 ;
                RECT 0.160 7.280 270.400 7.600 ;
                RECT 0.160 8.640 270.400 8.960 ;
                RECT 0.160 10.000 132.040 10.320 ;
                RECT 260.920 10.000 270.400 10.320 ;
                RECT 0.160 11.360 159.240 11.680 ;
                RECT 260.920 11.360 270.400 11.680 ;
                RECT 0.160 12.720 159.240 13.040 ;
                RECT 260.920 12.720 270.400 13.040 ;
                RECT 0.160 14.080 159.240 14.400 ;
                RECT 260.920 14.080 270.400 14.400 ;
                RECT 0.160 15.440 159.240 15.760 ;
                RECT 260.920 15.440 270.400 15.760 ;
                RECT 0.160 16.800 159.240 17.120 ;
                RECT 260.920 16.800 270.400 17.120 ;
                RECT 0.160 18.160 159.240 18.480 ;
                RECT 260.920 18.160 270.400 18.480 ;
                RECT 0.160 19.520 159.240 19.840 ;
                RECT 260.920 19.520 270.400 19.840 ;
                RECT 0.160 20.880 64.040 21.200 ;
                RECT 133.760 20.880 159.240 21.200 ;
                RECT 260.920 20.880 270.400 21.200 ;
                RECT 0.160 22.240 159.240 22.560 ;
                RECT 260.920 22.240 270.400 22.560 ;
                RECT 0.160 23.600 159.240 23.920 ;
                RECT 260.920 23.600 270.400 23.920 ;
                RECT 0.160 24.960 64.040 25.280 ;
                RECT 133.080 24.960 159.240 25.280 ;
                RECT 260.920 24.960 270.400 25.280 ;
                RECT 0.160 26.320 159.240 26.640 ;
                RECT 260.920 26.320 270.400 26.640 ;
                RECT 0.160 27.680 158.560 28.000 ;
                RECT 260.920 27.680 270.400 28.000 ;
                RECT 0.160 29.040 159.240 29.360 ;
                RECT 260.920 29.040 270.400 29.360 ;
                RECT 0.160 30.400 159.240 30.720 ;
                RECT 260.920 30.400 270.400 30.720 ;
                RECT 0.160 31.760 159.240 32.080 ;
                RECT 260.920 31.760 270.400 32.080 ;
                RECT 0.160 33.120 159.240 33.440 ;
                RECT 260.920 33.120 270.400 33.440 ;
                RECT 0.160 34.480 159.240 34.800 ;
                RECT 260.920 34.480 270.400 34.800 ;
                RECT 0.160 35.840 159.240 36.160 ;
                RECT 260.920 35.840 270.400 36.160 ;
                RECT 0.160 37.200 159.240 37.520 ;
                RECT 260.920 37.200 270.400 37.520 ;
                RECT 0.160 38.560 159.240 38.880 ;
                RECT 260.920 38.560 270.400 38.880 ;
                RECT 0.160 39.920 159.240 40.240 ;
                RECT 260.920 39.920 270.400 40.240 ;
                RECT 0.160 41.280 93.960 41.600 ;
                RECT 104.520 41.280 159.240 41.600 ;
                RECT 260.920 41.280 270.400 41.600 ;
                RECT 0.160 42.640 92.600 42.960 ;
                RECT 110.640 42.640 159.240 42.960 ;
                RECT 260.920 42.640 270.400 42.960 ;
                RECT 0.160 44.000 91.240 44.320 ;
                RECT 116.760 44.000 159.240 44.320 ;
                RECT 260.920 44.000 270.400 44.320 ;
                RECT 0.160 45.360 71.520 45.680 ;
                RECT 133.760 45.360 159.240 45.680 ;
                RECT 260.920 45.360 270.400 45.680 ;
                RECT 0.160 46.720 70.840 47.040 ;
                RECT 129.680 46.720 159.240 47.040 ;
                RECT 260.920 46.720 270.400 47.040 ;
                RECT 0.160 48.080 159.240 48.400 ;
                RECT 260.920 48.080 270.400 48.400 ;
                RECT 0.160 49.440 125.920 49.760 ;
                RECT 131.720 49.440 159.240 49.760 ;
                RECT 260.920 49.440 270.400 49.760 ;
                RECT 0.160 50.800 125.920 51.120 ;
                RECT 131.720 50.800 159.240 51.120 ;
                RECT 260.920 50.800 270.400 51.120 ;
                RECT 0.160 52.160 125.920 52.480 ;
                RECT 260.920 52.160 270.400 52.480 ;
                RECT 0.160 53.520 67.440 53.840 ;
                RECT 78.000 53.520 125.920 53.840 ;
                RECT 260.920 53.520 270.400 53.840 ;
                RECT 0.160 54.880 68.800 55.200 ;
                RECT 74.600 54.880 81.720 55.200 ;
                RECT 84.800 54.880 125.920 55.200 ;
                RECT 131.720 54.880 159.240 55.200 ;
                RECT 260.920 54.880 270.400 55.200 ;
                RECT 0.160 56.240 70.160 56.560 ;
                RECT 73.240 56.240 159.240 56.560 ;
                RECT 260.920 56.240 270.400 56.560 ;
                RECT 0.160 57.600 159.240 57.920 ;
                RECT 260.920 57.600 270.400 57.920 ;
                RECT 0.160 58.960 76.280 59.280 ;
                RECT 84.800 58.960 159.240 59.280 ;
                RECT 260.920 58.960 270.400 59.280 ;
                RECT 0.160 60.320 68.800 60.640 ;
                RECT 78.000 60.320 159.240 60.640 ;
                RECT 260.920 60.320 270.400 60.640 ;
                RECT 0.160 61.680 72.880 62.000 ;
                RECT 77.320 61.680 91.240 62.000 ;
                RECT 99.760 61.680 106.200 62.000 ;
                RECT 131.040 61.680 159.240 62.000 ;
                RECT 260.920 61.680 270.400 62.000 ;
                RECT 0.160 63.040 92.600 63.360 ;
                RECT 98.400 63.040 106.200 63.360 ;
                RECT 140.560 63.040 159.240 63.360 ;
                RECT 260.920 63.040 270.400 63.360 ;
                RECT 0.160 64.400 68.800 64.720 ;
                RECT 78.000 64.400 93.960 64.720 ;
                RECT 97.720 64.400 106.200 64.720 ;
                RECT 140.560 64.400 159.240 64.720 ;
                RECT 260.920 64.400 270.400 64.720 ;
                RECT 0.160 65.760 75.600 66.080 ;
                RECT 84.120 65.760 106.200 66.080 ;
                RECT 139.200 65.760 159.240 66.080 ;
                RECT 260.920 65.760 270.400 66.080 ;
                RECT 0.160 67.120 106.200 67.440 ;
                RECT 143.280 67.120 159.240 67.440 ;
                RECT 260.920 67.120 270.400 67.440 ;
                RECT 0.160 68.480 76.280 68.800 ;
                RECT 82.080 68.480 106.200 68.800 ;
                RECT 143.280 68.480 159.240 68.800 ;
                RECT 260.920 68.480 270.400 68.800 ;
                RECT 0.160 69.840 79.000 70.160 ;
                RECT 84.800 69.840 106.200 70.160 ;
                RECT 141.920 69.840 159.240 70.160 ;
                RECT 260.920 69.840 270.400 70.160 ;
                RECT 0.160 71.200 72.880 71.520 ;
                RECT 78.000 71.200 106.200 71.520 ;
                RECT 146.000 71.200 159.240 71.520 ;
                RECT 260.920 71.200 270.400 71.520 ;
                RECT 0.160 72.560 106.200 72.880 ;
                RECT 144.640 72.560 159.240 72.880 ;
                RECT 260.920 72.560 270.400 72.880 ;
                RECT 0.160 73.920 66.760 74.240 ;
                RECT 89.560 73.920 106.200 74.240 ;
                RECT 146.000 73.920 159.240 74.240 ;
                RECT 260.920 73.920 270.400 74.240 ;
                RECT 0.160 75.280 76.280 75.600 ;
                RECT 84.800 75.280 106.200 75.600 ;
                RECT 148.720 75.280 159.240 75.600 ;
                RECT 260.920 75.280 270.400 75.600 ;
                RECT 0.160 76.640 75.600 76.960 ;
                RECT 78.000 76.640 85.120 76.960 ;
                RECT 91.600 76.640 106.200 76.960 ;
                RECT 131.040 76.640 159.240 76.960 ;
                RECT 260.920 76.640 270.400 76.960 ;
                RECT 0.160 78.000 67.440 78.320 ;
                RECT 80.720 78.000 106.200 78.320 ;
                RECT 147.360 78.000 159.240 78.320 ;
                RECT 260.920 78.000 270.400 78.320 ;
                RECT 0.160 79.360 75.600 79.680 ;
                RECT 84.800 79.360 106.200 79.680 ;
                RECT 131.040 79.360 159.240 79.680 ;
                RECT 260.920 79.360 270.400 79.680 ;
                RECT 0.160 80.720 73.560 81.040 ;
                RECT 77.320 80.720 106.200 81.040 ;
                RECT 151.440 80.720 159.240 81.040 ;
                RECT 260.920 80.720 270.400 81.040 ;
                RECT 0.160 82.080 68.800 82.400 ;
                RECT 73.240 82.080 76.280 82.400 ;
                RECT 84.800 82.080 106.200 82.400 ;
                RECT 151.440 82.080 159.240 82.400 ;
                RECT 260.920 82.080 270.400 82.400 ;
                RECT 0.160 83.440 71.520 83.760 ;
                RECT 75.280 83.440 106.200 83.760 ;
                RECT 154.160 83.440 159.240 83.760 ;
                RECT 260.920 83.440 270.400 83.760 ;
                RECT 0.160 84.800 68.800 85.120 ;
                RECT 71.880 84.800 106.200 85.120 ;
                RECT 152.800 84.800 159.240 85.120 ;
                RECT 260.920 84.800 270.400 85.120 ;
                RECT 0.160 86.160 72.880 86.480 ;
                RECT 78.000 86.160 106.200 86.480 ;
                RECT 154.160 86.160 159.240 86.480 ;
                RECT 260.920 86.160 270.400 86.480 ;
                RECT 0.160 87.520 68.800 87.840 ;
                RECT 83.440 87.520 106.200 87.840 ;
                RECT 131.040 87.520 159.240 87.840 ;
                RECT 260.920 87.520 270.400 87.840 ;
                RECT 0.160 88.880 106.200 89.200 ;
                RECT 156.880 88.880 159.240 89.200 ;
                RECT 260.920 88.880 270.400 89.200 ;
                RECT 0.160 90.240 75.600 90.560 ;
                RECT 77.320 90.240 106.200 90.560 ;
                RECT 156.880 90.240 159.240 90.560 ;
                RECT 260.920 90.240 270.400 90.560 ;
                RECT 0.160 91.600 76.280 91.920 ;
                RECT 78.680 91.600 106.200 91.920 ;
                RECT 155.520 91.600 159.240 91.920 ;
                RECT 260.920 91.600 270.400 91.920 ;
                RECT 0.160 92.960 67.440 93.280 ;
                RECT 74.600 92.960 75.600 93.280 ;
                RECT 77.320 92.960 106.200 93.280 ;
                RECT 260.920 92.960 270.400 93.280 ;
                RECT 0.160 94.320 67.440 94.640 ;
                RECT 78.000 94.320 106.200 94.640 ;
                RECT 260.920 94.320 270.400 94.640 ;
                RECT 0.160 95.680 70.160 96.000 ;
                RECT 84.800 95.680 106.200 96.000 ;
                RECT 131.040 95.680 159.240 96.000 ;
                RECT 260.920 95.680 270.400 96.000 ;
                RECT 0.160 97.040 75.600 97.360 ;
                RECT 78.680 97.040 82.400 97.360 ;
                RECT 84.800 97.040 159.240 97.360 ;
                RECT 260.920 97.040 270.400 97.360 ;
                RECT 0.160 98.400 159.240 98.720 ;
                RECT 260.920 98.400 270.400 98.720 ;
                RECT 0.160 99.760 134.760 100.080 ;
                RECT 260.920 99.760 270.400 100.080 ;
                RECT 0.160 101.120 63.360 101.440 ;
                RECT 80.720 101.120 156.520 101.440 ;
                RECT 260.920 101.120 270.400 101.440 ;
                RECT 0.160 102.480 45.680 102.800 ;
                RECT 63.720 102.480 153.800 102.800 ;
                RECT 260.920 102.480 270.400 102.800 ;
                RECT 0.160 103.840 45.680 104.160 ;
                RECT 63.720 103.840 151.080 104.160 ;
                RECT 260.920 103.840 270.400 104.160 ;
                RECT 0.160 105.200 45.680 105.520 ;
                RECT 63.720 105.200 148.360 105.520 ;
                RECT 260.920 105.200 270.400 105.520 ;
                RECT 0.160 106.560 45.680 106.880 ;
                RECT 63.720 106.560 79.000 106.880 ;
                RECT 86.840 106.560 145.640 106.880 ;
                RECT 260.920 106.560 270.400 106.880 ;
                RECT 0.160 107.920 45.680 108.240 ;
                RECT 63.720 107.920 72.200 108.240 ;
                RECT 84.800 107.920 140.200 108.240 ;
                RECT 260.920 107.920 270.400 108.240 ;
                RECT 0.160 109.280 45.680 109.600 ;
                RECT 63.720 109.280 137.480 109.600 ;
                RECT 260.920 109.280 270.400 109.600 ;
                RECT 0.160 110.640 45.680 110.960 ;
                RECT 63.720 110.640 66.760 110.960 ;
                RECT 71.880 110.640 137.480 110.960 ;
                RECT 260.920 110.640 270.400 110.960 ;
                RECT 0.160 112.000 45.680 112.320 ;
                RECT 63.720 112.000 159.240 112.320 ;
                RECT 260.920 112.000 270.400 112.320 ;
                RECT 0.160 113.360 45.680 113.680 ;
                RECT 63.720 113.360 159.240 113.680 ;
                RECT 260.920 113.360 270.400 113.680 ;
                RECT 0.160 114.720 45.680 115.040 ;
                RECT 63.720 114.720 159.240 115.040 ;
                RECT 260.920 114.720 270.400 115.040 ;
                RECT 0.160 116.080 45.680 116.400 ;
                RECT 63.720 116.080 159.240 116.400 ;
                RECT 260.920 116.080 270.400 116.400 ;
                RECT 0.160 117.440 45.680 117.760 ;
                RECT 64.400 117.440 82.400 117.760 ;
                RECT 84.800 117.440 125.240 117.760 ;
                RECT 131.040 117.440 159.240 117.760 ;
                RECT 260.920 117.440 270.400 117.760 ;
                RECT 0.160 118.800 45.680 119.120 ;
                RECT 63.720 118.800 125.240 119.120 ;
                RECT 131.040 118.800 159.240 119.120 ;
                RECT 260.920 118.800 270.400 119.120 ;
                RECT 0.160 120.160 45.680 120.480 ;
                RECT 63.720 120.160 68.800 120.480 ;
                RECT 73.920 120.160 125.240 120.480 ;
                RECT 131.040 120.160 159.240 120.480 ;
                RECT 260.920 120.160 270.400 120.480 ;
                RECT 0.160 121.520 45.680 121.840 ;
                RECT 63.720 121.520 125.240 121.840 ;
                RECT 131.040 121.520 159.240 121.840 ;
                RECT 260.920 121.520 270.400 121.840 ;
                RECT 0.160 122.880 45.680 123.200 ;
                RECT 63.720 122.880 125.240 123.200 ;
                RECT 131.040 122.880 159.240 123.200 ;
                RECT 260.920 122.880 270.400 123.200 ;
                RECT 0.160 124.240 45.680 124.560 ;
                RECT 63.720 124.240 159.240 124.560 ;
                RECT 260.920 124.240 270.400 124.560 ;
                RECT 0.160 125.600 45.680 125.920 ;
                RECT 63.720 125.600 71.520 125.920 ;
                RECT 74.600 125.600 75.600 125.920 ;
                RECT 84.120 125.600 138.840 125.920 ;
                RECT 260.920 125.600 270.400 125.920 ;
                RECT 0.160 126.960 45.680 127.280 ;
                RECT 63.720 126.960 68.800 127.280 ;
                RECT 71.880 126.960 141.560 127.280 ;
                RECT 260.920 126.960 270.400 127.280 ;
                RECT 0.160 128.320 45.680 128.640 ;
                RECT 63.720 128.320 144.280 128.640 ;
                RECT 260.920 128.320 270.400 128.640 ;
                RECT 0.160 129.680 45.680 130.000 ;
                RECT 63.720 129.680 108.240 130.000 ;
                RECT 130.360 129.680 147.000 130.000 ;
                RECT 260.920 129.680 270.400 130.000 ;
                RECT 0.160 131.040 45.680 131.360 ;
                RECT 63.720 131.040 108.240 131.360 ;
                RECT 130.360 131.040 149.720 131.360 ;
                RECT 260.920 131.040 270.400 131.360 ;
                RECT 0.160 132.400 45.680 132.720 ;
                RECT 63.720 132.400 108.240 132.720 ;
                RECT 130.360 132.400 152.440 132.720 ;
                RECT 260.920 132.400 270.400 132.720 ;
                RECT 0.160 133.760 45.680 134.080 ;
                RECT 63.720 133.760 108.240 134.080 ;
                RECT 130.360 133.760 155.160 134.080 ;
                RECT 260.920 133.760 270.400 134.080 ;
                RECT 0.160 135.120 45.680 135.440 ;
                RECT 63.720 135.120 108.240 135.440 ;
                RECT 260.920 135.120 270.400 135.440 ;
                RECT 0.160 136.480 70.160 136.800 ;
                RECT 74.600 136.480 108.240 136.800 ;
                RECT 260.920 136.480 270.400 136.800 ;
                RECT 0.160 137.840 108.240 138.160 ;
                RECT 130.360 137.840 159.240 138.160 ;
                RECT 260.920 137.840 270.400 138.160 ;
                RECT 0.160 139.200 26.640 139.520 ;
                RECT 45.360 139.200 108.240 139.520 ;
                RECT 130.360 139.200 159.240 139.520 ;
                RECT 260.920 139.200 270.400 139.520 ;
                RECT 0.160 140.560 26.640 140.880 ;
                RECT 45.360 140.560 72.880 140.880 ;
                RECT 78.680 140.560 108.240 140.880 ;
                RECT 130.360 140.560 159.240 140.880 ;
                RECT 260.920 140.560 270.400 140.880 ;
                RECT 0.160 141.920 26.640 142.240 ;
                RECT 45.360 141.920 51.120 142.240 ;
                RECT 58.960 141.920 108.240 142.240 ;
                RECT 130.360 141.920 159.240 142.240 ;
                RECT 260.920 141.920 270.400 142.240 ;
                RECT 0.160 143.280 26.640 143.600 ;
                RECT 63.040 143.280 108.240 143.600 ;
                RECT 130.360 143.280 159.240 143.600 ;
                RECT 260.920 143.280 270.400 143.600 ;
                RECT 0.160 144.640 26.640 144.960 ;
                RECT 63.040 144.640 108.240 144.960 ;
                RECT 260.920 144.640 270.400 144.960 ;
                RECT 0.160 146.000 26.640 146.320 ;
                RECT 45.360 146.000 51.120 146.320 ;
                RECT 58.960 146.000 67.440 146.320 ;
                RECT 77.320 146.000 108.240 146.320 ;
                RECT 260.920 146.000 270.400 146.320 ;
                RECT 0.160 147.360 18.480 147.680 ;
                RECT 58.280 147.360 108.240 147.680 ;
                RECT 130.360 147.360 270.400 147.680 ;
                RECT 0.160 148.720 57.920 149.040 ;
                RECT 105.200 148.720 270.400 149.040 ;
                RECT 0.160 150.080 156.520 150.400 ;
                RECT 263.640 150.080 270.400 150.400 ;
                RECT 0.160 151.440 156.520 151.760 ;
                RECT 263.640 151.440 270.400 151.760 ;
                RECT 0.160 152.800 156.520 153.120 ;
                RECT 263.640 152.800 270.400 153.120 ;
                RECT 0.160 154.160 62.000 154.480 ;
                RECT 68.480 154.160 70.160 154.480 ;
                RECT 82.760 154.160 115.720 154.480 ;
                RECT 263.640 154.160 270.400 154.480 ;
                RECT 0.160 155.520 59.960 155.840 ;
                RECT 82.080 155.520 99.400 155.840 ;
                RECT 105.200 155.520 115.720 155.840 ;
                RECT 263.640 155.520 270.400 155.840 ;
                RECT 0.160 156.880 59.960 157.200 ;
                RECT 80.720 156.880 95.320 157.200 ;
                RECT 105.200 156.880 115.720 157.200 ;
                RECT 263.640 156.880 270.400 157.200 ;
                RECT 0.160 158.240 59.960 158.560 ;
                RECT 70.520 158.240 95.320 158.560 ;
                RECT 105.200 158.240 115.720 158.560 ;
                RECT 263.640 158.240 270.400 158.560 ;
                RECT 0.160 159.600 95.320 159.920 ;
                RECT 105.200 159.600 115.720 159.920 ;
                RECT 263.640 159.600 270.400 159.920 ;
                RECT 0.160 160.960 59.960 161.280 ;
                RECT 70.520 160.960 95.320 161.280 ;
                RECT 105.200 160.960 115.720 161.280 ;
                RECT 263.640 160.960 270.400 161.280 ;
                RECT 0.160 162.320 59.960 162.640 ;
                RECT 70.520 162.320 115.720 162.640 ;
                RECT 263.640 162.320 270.400 162.640 ;
                RECT 0.160 163.680 95.320 164.000 ;
                RECT 105.200 163.680 115.720 164.000 ;
                RECT 263.640 163.680 270.400 164.000 ;
                RECT 0.160 165.040 95.320 165.360 ;
                RECT 105.200 165.040 115.720 165.360 ;
                RECT 263.640 165.040 270.400 165.360 ;
                RECT 0.160 166.400 95.320 166.720 ;
                RECT 105.200 166.400 115.720 166.720 ;
                RECT 263.640 166.400 270.400 166.720 ;
                RECT 0.160 167.760 18.480 168.080 ;
                RECT 55.560 167.760 68.800 168.080 ;
                RECT 71.200 167.760 95.320 168.080 ;
                RECT 105.200 167.760 115.720 168.080 ;
                RECT 263.640 167.760 270.400 168.080 ;
                RECT 0.160 169.120 17.800 169.440 ;
                RECT 55.560 169.120 68.800 169.440 ;
                RECT 71.880 169.120 95.320 169.440 ;
                RECT 105.200 169.120 115.720 169.440 ;
                RECT 263.640 169.120 270.400 169.440 ;
                RECT 0.160 170.480 17.120 170.800 ;
                RECT 55.560 170.480 115.720 170.800 ;
                RECT 263.640 170.480 270.400 170.800 ;
                RECT 0.160 171.840 16.440 172.160 ;
                RECT 55.560 171.840 96.000 172.160 ;
                RECT 105.200 171.840 115.720 172.160 ;
                RECT 263.640 171.840 270.400 172.160 ;
                RECT 0.160 173.200 95.320 173.520 ;
                RECT 105.200 173.200 115.720 173.520 ;
                RECT 263.640 173.200 270.400 173.520 ;
                RECT 0.160 174.560 15.760 174.880 ;
                RECT 55.560 174.560 95.320 174.880 ;
                RECT 105.200 174.560 115.720 174.880 ;
                RECT 263.640 174.560 270.400 174.880 ;
                RECT 0.160 175.920 15.080 176.240 ;
                RECT 55.560 175.920 95.320 176.240 ;
                RECT 105.200 175.920 115.720 176.240 ;
                RECT 263.640 175.920 270.400 176.240 ;
                RECT 0.160 177.280 95.320 177.600 ;
                RECT 105.200 177.280 115.720 177.600 ;
                RECT 263.640 177.280 270.400 177.600 ;
                RECT 0.160 178.640 14.400 178.960 ;
                RECT 55.560 178.640 115.720 178.960 ;
                RECT 263.640 178.640 270.400 178.960 ;
                RECT 0.160 180.000 13.720 180.320 ;
                RECT 55.560 180.000 68.800 180.320 ;
                RECT 73.920 180.000 95.320 180.320 ;
                RECT 105.200 180.000 115.720 180.320 ;
                RECT 263.640 180.000 270.400 180.320 ;
                RECT 0.160 181.360 95.320 181.680 ;
                RECT 105.200 181.360 115.720 181.680 ;
                RECT 263.640 181.360 270.400 181.680 ;
                RECT 0.160 182.720 13.040 183.040 ;
                RECT 55.560 182.720 68.800 183.040 ;
                RECT 73.240 182.720 95.320 183.040 ;
                RECT 105.200 182.720 115.720 183.040 ;
                RECT 263.640 182.720 270.400 183.040 ;
                RECT 0.160 184.080 12.360 184.400 ;
                RECT 55.560 184.080 68.800 184.400 ;
                RECT 72.560 184.080 95.320 184.400 ;
                RECT 105.200 184.080 115.720 184.400 ;
                RECT 263.640 184.080 270.400 184.400 ;
                RECT 0.160 185.440 11.680 185.760 ;
                RECT 55.560 185.440 68.800 185.760 ;
                RECT 71.880 185.440 95.320 185.760 ;
                RECT 104.520 185.440 115.720 185.760 ;
                RECT 263.640 185.440 270.400 185.760 ;
                RECT 0.160 186.800 11.000 187.120 ;
                RECT 55.560 186.800 99.400 187.120 ;
                RECT 105.200 186.800 115.720 187.120 ;
                RECT 263.640 186.800 270.400 187.120 ;
                RECT 0.160 188.160 96.680 188.480 ;
                RECT 105.200 188.160 115.720 188.480 ;
                RECT 263.640 188.160 270.400 188.480 ;
                RECT 0.160 189.520 96.680 189.840 ;
                RECT 105.200 189.520 115.720 189.840 ;
                RECT 263.640 189.520 270.400 189.840 ;
                RECT 0.160 190.880 96.680 191.200 ;
                RECT 105.200 190.880 115.720 191.200 ;
                RECT 263.640 190.880 270.400 191.200 ;
                RECT 0.160 192.240 96.680 192.560 ;
                RECT 105.200 192.240 115.720 192.560 ;
                RECT 263.640 192.240 270.400 192.560 ;
                RECT 0.160 193.600 73.560 193.920 ;
                RECT 82.760 193.600 115.720 193.920 ;
                RECT 263.640 193.600 270.400 193.920 ;
                RECT 0.160 194.960 72.200 195.280 ;
                RECT 82.080 194.960 101.440 195.280 ;
                RECT 105.200 194.960 115.720 195.280 ;
                RECT 263.640 194.960 270.400 195.280 ;
                RECT 0.160 196.320 70.840 196.640 ;
                RECT 80.720 196.320 95.320 196.640 ;
                RECT 105.200 196.320 115.720 196.640 ;
                RECT 263.640 196.320 270.400 196.640 ;
                RECT 0.160 197.680 95.320 198.000 ;
                RECT 105.200 197.680 115.720 198.000 ;
                RECT 263.640 197.680 270.400 198.000 ;
                RECT 0.160 199.040 95.320 199.360 ;
                RECT 105.200 199.040 115.720 199.360 ;
                RECT 263.640 199.040 270.400 199.360 ;
                RECT 0.160 200.400 95.320 200.720 ;
                RECT 105.200 200.400 115.720 200.720 ;
                RECT 263.640 200.400 270.400 200.720 ;
                RECT 0.160 201.760 95.320 202.080 ;
                RECT 97.720 201.760 115.720 202.080 ;
                RECT 263.640 201.760 270.400 202.080 ;
                RECT 0.160 203.120 96.680 203.440 ;
                RECT 105.200 203.120 115.720 203.440 ;
                RECT 263.640 203.120 270.400 203.440 ;
                RECT 0.160 204.480 95.320 204.800 ;
                RECT 105.200 204.480 115.720 204.800 ;
                RECT 263.640 204.480 270.400 204.800 ;
                RECT 0.160 205.840 95.320 206.160 ;
                RECT 105.200 205.840 115.720 206.160 ;
                RECT 263.640 205.840 270.400 206.160 ;
                RECT 0.160 207.200 95.320 207.520 ;
                RECT 105.200 207.200 115.720 207.520 ;
                RECT 263.640 207.200 270.400 207.520 ;
                RECT 0.160 208.560 95.320 208.880 ;
                RECT 105.200 208.560 115.720 208.880 ;
                RECT 263.640 208.560 270.400 208.880 ;
                RECT 0.160 209.920 115.720 210.240 ;
                RECT 263.640 209.920 270.400 210.240 ;
                RECT 0.160 211.280 96.680 211.600 ;
                RECT 105.200 211.280 115.720 211.600 ;
                RECT 263.640 211.280 270.400 211.600 ;
                RECT 0.160 212.640 95.320 212.960 ;
                RECT 105.200 212.640 115.720 212.960 ;
                RECT 263.640 212.640 270.400 212.960 ;
                RECT 0.160 214.000 95.320 214.320 ;
                RECT 105.200 214.000 115.720 214.320 ;
                RECT 263.640 214.000 270.400 214.320 ;
                RECT 0.160 215.360 95.320 215.680 ;
                RECT 105.200 215.360 115.720 215.680 ;
                RECT 263.640 215.360 270.400 215.680 ;
                RECT 0.160 216.720 95.320 217.040 ;
                RECT 105.200 216.720 115.720 217.040 ;
                RECT 263.640 216.720 270.400 217.040 ;
                RECT 0.160 218.080 115.720 218.400 ;
                RECT 263.640 218.080 270.400 218.400 ;
                RECT 0.160 219.440 95.320 219.760 ;
                RECT 105.200 219.440 115.720 219.760 ;
                RECT 263.640 219.440 270.400 219.760 ;
                RECT 0.160 220.800 95.320 221.120 ;
                RECT 105.200 220.800 115.720 221.120 ;
                RECT 263.640 220.800 270.400 221.120 ;
                RECT 0.160 222.160 95.320 222.480 ;
                RECT 105.200 222.160 115.720 222.480 ;
                RECT 263.640 222.160 270.400 222.480 ;
                RECT 0.160 223.520 95.320 223.840 ;
                RECT 105.200 223.520 115.720 223.840 ;
                RECT 263.640 223.520 270.400 223.840 ;
                RECT 0.160 224.880 95.320 225.200 ;
                RECT 105.200 224.880 115.720 225.200 ;
                RECT 263.640 224.880 270.400 225.200 ;
                RECT 0.160 226.240 115.720 226.560 ;
                RECT 263.640 226.240 270.400 226.560 ;
                RECT 0.160 227.600 97.360 227.920 ;
                RECT 105.200 227.600 115.720 227.920 ;
                RECT 263.640 227.600 270.400 227.920 ;
                RECT 0.160 228.960 97.360 229.280 ;
                RECT 105.200 228.960 115.720 229.280 ;
                RECT 263.640 228.960 270.400 229.280 ;
                RECT 0.160 230.320 97.360 230.640 ;
                RECT 105.200 230.320 115.720 230.640 ;
                RECT 263.640 230.320 270.400 230.640 ;
                RECT 0.160 231.680 97.360 232.000 ;
                RECT 105.200 231.680 115.720 232.000 ;
                RECT 263.640 231.680 270.400 232.000 ;
                RECT 0.160 233.040 115.720 233.360 ;
                RECT 263.640 233.040 270.400 233.360 ;
                RECT 0.160 234.400 99.400 234.720 ;
                RECT 105.200 234.400 115.720 234.720 ;
                RECT 263.640 234.400 270.400 234.720 ;
                RECT 0.160 235.760 98.040 236.080 ;
                RECT 105.200 235.760 115.720 236.080 ;
                RECT 263.640 235.760 270.400 236.080 ;
                RECT 0.160 237.120 98.040 237.440 ;
                RECT 105.200 237.120 115.720 237.440 ;
                RECT 263.640 237.120 270.400 237.440 ;
                RECT 0.160 238.480 98.040 238.800 ;
                RECT 105.200 238.480 115.720 238.800 ;
                RECT 263.640 238.480 270.400 238.800 ;
                RECT 0.160 239.840 98.040 240.160 ;
                RECT 105.200 239.840 115.720 240.160 ;
                RECT 263.640 239.840 270.400 240.160 ;
                RECT 0.160 241.200 115.720 241.520 ;
                RECT 263.640 241.200 270.400 241.520 ;
                RECT 0.160 242.560 101.440 242.880 ;
                RECT 105.200 242.560 115.720 242.880 ;
                RECT 263.640 242.560 270.400 242.880 ;
                RECT 0.160 243.920 102.120 244.240 ;
                RECT 105.200 243.920 115.720 244.240 ;
                RECT 263.640 243.920 270.400 244.240 ;
                RECT 0.160 245.280 98.040 245.600 ;
                RECT 105.200 245.280 115.720 245.600 ;
                RECT 263.640 245.280 270.400 245.600 ;
                RECT 0.160 246.640 98.040 246.960 ;
                RECT 105.200 246.640 115.720 246.960 ;
                RECT 263.640 246.640 270.400 246.960 ;
                RECT 0.160 248.000 98.040 248.320 ;
                RECT 105.200 248.000 115.720 248.320 ;
                RECT 263.640 248.000 270.400 248.320 ;
                RECT 0.160 249.360 115.720 249.680 ;
                RECT 263.640 249.360 270.400 249.680 ;
                RECT 0.160 250.720 98.720 251.040 ;
                RECT 105.200 250.720 115.720 251.040 ;
                RECT 263.640 250.720 270.400 251.040 ;
                RECT 0.160 252.080 98.720 252.400 ;
                RECT 105.200 252.080 115.720 252.400 ;
                RECT 263.640 252.080 270.400 252.400 ;
                RECT 0.160 253.440 100.080 253.760 ;
                RECT 105.200 253.440 115.720 253.760 ;
                RECT 263.640 253.440 270.400 253.760 ;
                RECT 0.160 254.800 98.720 255.120 ;
                RECT 105.200 254.800 115.720 255.120 ;
                RECT 263.640 254.800 270.400 255.120 ;
                RECT 0.160 256.160 98.720 256.480 ;
                RECT 105.200 256.160 115.720 256.480 ;
                RECT 263.640 256.160 270.400 256.480 ;
                RECT 0.160 257.520 115.720 257.840 ;
                RECT 263.640 257.520 270.400 257.840 ;
                RECT 0.160 258.880 98.720 259.200 ;
                RECT 105.200 258.880 115.720 259.200 ;
                RECT 263.640 258.880 270.400 259.200 ;
                RECT 0.160 260.240 98.720 260.560 ;
                RECT 105.200 260.240 115.720 260.560 ;
                RECT 263.640 260.240 270.400 260.560 ;
                RECT 0.160 261.600 98.720 261.920 ;
                RECT 105.200 261.600 115.720 261.920 ;
                RECT 263.640 261.600 270.400 261.920 ;
                RECT 0.160 262.960 102.800 263.280 ;
                RECT 105.200 262.960 115.720 263.280 ;
                RECT 263.640 262.960 270.400 263.280 ;
                RECT 0.160 264.320 98.720 264.640 ;
                RECT 105.200 264.320 115.720 264.640 ;
                RECT 263.640 264.320 270.400 264.640 ;
                RECT 0.160 265.680 115.720 266.000 ;
                RECT 263.640 265.680 270.400 266.000 ;
                RECT 0.160 267.040 98.720 267.360 ;
                RECT 105.200 267.040 115.720 267.360 ;
                RECT 263.640 267.040 270.400 267.360 ;
                RECT 0.160 268.400 98.720 268.720 ;
                RECT 105.200 268.400 115.720 268.720 ;
                RECT 263.640 268.400 270.400 268.720 ;
                RECT 0.160 269.760 98.720 270.080 ;
                RECT 105.200 269.760 115.720 270.080 ;
                RECT 263.640 269.760 270.400 270.080 ;
                RECT 0.160 271.120 98.720 271.440 ;
                RECT 105.200 271.120 115.720 271.440 ;
                RECT 263.640 271.120 270.400 271.440 ;
                RECT 0.160 272.480 115.720 272.800 ;
                RECT 263.640 272.480 270.400 272.800 ;
                RECT 0.160 273.840 101.440 274.160 ;
                RECT 105.200 273.840 115.720 274.160 ;
                RECT 263.640 273.840 270.400 274.160 ;
                RECT 0.160 275.200 98.720 275.520 ;
                RECT 105.200 275.200 115.720 275.520 ;
                RECT 263.640 275.200 270.400 275.520 ;
                RECT 0.160 276.560 98.720 276.880 ;
                RECT 105.200 276.560 115.720 276.880 ;
                RECT 263.640 276.560 270.400 276.880 ;
                RECT 0.160 277.920 98.720 278.240 ;
                RECT 105.200 277.920 115.720 278.240 ;
                RECT 263.640 277.920 270.400 278.240 ;
                RECT 0.160 279.280 98.720 279.600 ;
                RECT 105.200 279.280 115.720 279.600 ;
                RECT 263.640 279.280 270.400 279.600 ;
                RECT 0.160 280.640 115.720 280.960 ;
                RECT 263.640 280.640 270.400 280.960 ;
                RECT 0.160 282.000 115.720 282.320 ;
                RECT 263.640 282.000 270.400 282.320 ;
                RECT 0.160 283.360 156.520 283.680 ;
                RECT 263.640 283.360 270.400 283.680 ;
                RECT 0.160 284.720 156.520 285.040 ;
                RECT 263.640 284.720 270.400 285.040 ;
                RECT 0.160 286.080 270.400 286.400 ;
                RECT 0.160 287.440 270.400 287.760 ;
                RECT 0.160 288.800 270.400 289.120 ;
                RECT 0.160 290.160 270.400 290.480 ;
                RECT 0.160 291.520 270.400 291.840 ;
                RECT 0.160 0.160 270.400 1.520 ;
                RECT 0.160 295.560 270.400 296.920 ;
                RECT 160.660 32.015 166.460 33.385 ;
                RECT 253.360 32.015 259.160 33.385 ;
                RECT 160.660 36.485 166.460 37.425 ;
                RECT 253.360 36.485 259.160 37.425 ;
                RECT 160.660 40.675 166.460 41.885 ;
                RECT 253.360 40.675 259.160 41.885 ;
                RECT 160.660 45.275 166.460 46.485 ;
                RECT 253.360 45.275 259.160 46.485 ;
                RECT 160.660 85.575 259.160 85.865 ;
                RECT 160.660 53.100 259.160 54.900 ;
                RECT 160.660 80.150 259.160 82.240 ;
                RECT 160.660 72.470 259.160 73.270 ;
                RECT 160.660 114.215 259.160 116.015 ;
                RECT 160.660 64.570 259.160 65.370 ;
                RECT 160.660 67.580 259.160 68.380 ;
                RECT 160.660 140.205 259.160 142.805 ;
                RECT 160.660 16.260 259.160 18.060 ;
                RECT 120.860 153.875 122.780 281.855 ;
                RECT 124.700 153.875 126.620 281.855 ;
                RECT 139.690 153.875 141.610 281.855 ;
                RECT 143.530 153.875 145.450 281.855 ;
                RECT 147.370 153.875 149.290 281.855 ;
                RECT 151.210 153.875 153.130 281.855 ;
                RECT 109.235 61.175 111.155 96.575 ;
                RECT 115.995 61.175 117.915 96.575 ;
                RECT 124.705 61.175 126.625 96.575 ;
                RECT 128.545 61.175 130.465 96.575 ;
                RECT 112.440 129.020 114.360 147.240 ;
                RECT 119.715 129.020 121.465 147.240 ;
                RECT 127.895 129.020 129.815 147.240 ;
                RECT 128.755 117.860 130.675 123.020 ;
                RECT 129.055 50.015 130.805 55.175 ;
                RECT 60.480 156.145 69.640 156.895 ;
                RECT 60.480 160.900 69.640 162.820 ;
                RECT 46.620 143.930 62.660 144.730 ;
                RECT 27.420 143.505 44.660 146.215 ;
        END 
    END vdd 
    PIN vss 
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT 
            LAYER met2 ;
                RECT 2.880 5.240 172.160 5.560 ;
                RECT 250.040 5.240 267.680 5.560 ;
                RECT 2.880 6.600 267.680 6.920 ;
                RECT 2.880 7.960 267.680 8.280 ;
                RECT 2.880 9.320 132.720 9.640 ;
                RECT 165.040 9.320 267.680 9.640 ;
                RECT 2.880 10.680 159.240 11.000 ;
                RECT 260.920 10.680 267.680 11.000 ;
                RECT 2.880 12.040 159.240 12.360 ;
                RECT 260.920 12.040 267.680 12.360 ;
                RECT 2.880 13.400 159.240 13.720 ;
                RECT 260.920 13.400 267.680 13.720 ;
                RECT 2.880 14.760 159.240 15.080 ;
                RECT 260.920 14.760 267.680 15.080 ;
                RECT 2.880 16.120 159.240 16.440 ;
                RECT 260.920 16.120 267.680 16.440 ;
                RECT 2.880 17.480 159.240 17.800 ;
                RECT 260.920 17.480 267.680 17.800 ;
                RECT 2.880 18.840 159.240 19.160 ;
                RECT 260.920 18.840 267.680 19.160 ;
                RECT 2.880 20.200 64.040 20.520 ;
                RECT 133.760 20.200 159.240 20.520 ;
                RECT 260.920 20.200 267.680 20.520 ;
                RECT 2.880 21.560 159.240 21.880 ;
                RECT 260.920 21.560 267.680 21.880 ;
                RECT 2.880 22.920 159.240 23.240 ;
                RECT 260.920 22.920 267.680 23.240 ;
                RECT 2.880 24.280 64.040 24.600 ;
                RECT 133.080 24.280 159.240 24.600 ;
                RECT 260.920 24.280 267.680 24.600 ;
                RECT 2.880 25.640 159.240 25.960 ;
                RECT 260.920 25.640 267.680 25.960 ;
                RECT 2.880 27.000 159.240 27.320 ;
                RECT 260.920 27.000 267.680 27.320 ;
                RECT 2.880 28.360 158.560 28.680 ;
                RECT 260.920 28.360 267.680 28.680 ;
                RECT 2.880 29.720 159.240 30.040 ;
                RECT 260.920 29.720 267.680 30.040 ;
                RECT 2.880 31.080 159.240 31.400 ;
                RECT 260.920 31.080 267.680 31.400 ;
                RECT 2.880 32.440 159.240 32.760 ;
                RECT 260.920 32.440 267.680 32.760 ;
                RECT 2.880 33.800 159.240 34.120 ;
                RECT 260.920 33.800 267.680 34.120 ;
                RECT 2.880 35.160 159.240 35.480 ;
                RECT 260.920 35.160 267.680 35.480 ;
                RECT 2.880 36.520 159.240 36.840 ;
                RECT 260.920 36.520 267.680 36.840 ;
                RECT 2.880 37.880 159.240 38.200 ;
                RECT 260.920 37.880 267.680 38.200 ;
                RECT 2.880 39.240 159.240 39.560 ;
                RECT 260.920 39.240 267.680 39.560 ;
                RECT 2.880 40.600 94.640 40.920 ;
                RECT 105.880 40.600 159.240 40.920 ;
                RECT 260.920 40.600 267.680 40.920 ;
                RECT 2.880 41.960 93.280 42.280 ;
                RECT 112.000 41.960 159.240 42.280 ;
                RECT 260.920 41.960 267.680 42.280 ;
                RECT 2.880 43.320 91.920 43.640 ;
                RECT 118.120 43.320 159.240 43.640 ;
                RECT 260.920 43.320 267.680 43.640 ;
                RECT 2.880 44.680 68.800 45.000 ;
                RECT 133.080 44.680 159.240 45.000 ;
                RECT 260.920 44.680 267.680 45.000 ;
                RECT 2.880 46.040 70.160 46.360 ;
                RECT 123.560 46.040 159.240 46.360 ;
                RECT 260.920 46.040 267.680 46.360 ;
                RECT 2.880 47.400 159.240 47.720 ;
                RECT 260.920 47.400 267.680 47.720 ;
                RECT 2.880 48.760 159.240 49.080 ;
                RECT 260.920 48.760 267.680 49.080 ;
                RECT 2.880 50.120 125.920 50.440 ;
                RECT 131.720 50.120 159.240 50.440 ;
                RECT 260.920 50.120 267.680 50.440 ;
                RECT 2.880 51.480 125.920 51.800 ;
                RECT 260.920 51.480 267.680 51.800 ;
                RECT 2.880 52.840 67.440 53.160 ;
                RECT 78.000 52.840 125.920 53.160 ;
                RECT 260.920 52.840 267.680 53.160 ;
                RECT 2.880 54.200 68.800 54.520 ;
                RECT 70.520 54.200 89.880 54.520 ;
                RECT 122.880 54.200 125.920 54.520 ;
                RECT 131.720 54.200 159.240 54.520 ;
                RECT 260.920 54.200 267.680 54.520 ;
                RECT 2.880 55.560 70.160 55.880 ;
                RECT 74.600 55.560 81.720 55.880 ;
                RECT 84.800 55.560 159.240 55.880 ;
                RECT 260.920 55.560 267.680 55.880 ;
                RECT 2.880 56.920 70.160 57.240 ;
                RECT 73.240 56.920 159.240 57.240 ;
                RECT 260.920 56.920 267.680 57.240 ;
                RECT 2.880 58.280 76.280 58.600 ;
                RECT 84.800 58.280 159.240 58.600 ;
                RECT 260.920 58.280 267.680 58.600 ;
                RECT 2.880 59.640 71.520 59.960 ;
                RECT 78.000 59.640 159.240 59.960 ;
                RECT 260.920 59.640 267.680 59.960 ;
                RECT 2.880 61.000 68.800 61.320 ;
                RECT 78.000 61.000 106.200 61.320 ;
                RECT 131.040 61.000 159.240 61.320 ;
                RECT 260.920 61.000 267.680 61.320 ;
                RECT 2.880 62.360 91.920 62.680 ;
                RECT 99.080 62.360 106.200 62.680 ;
                RECT 131.040 62.360 159.240 62.680 ;
                RECT 260.920 62.360 267.680 62.680 ;
                RECT 2.880 63.720 68.800 64.040 ;
                RECT 78.000 63.720 93.280 64.040 ;
                RECT 97.720 63.720 106.200 64.040 ;
                RECT 139.200 63.720 159.240 64.040 ;
                RECT 260.920 63.720 267.680 64.040 ;
                RECT 2.880 65.080 76.280 65.400 ;
                RECT 84.120 65.080 94.640 65.400 ;
                RECT 97.040 65.080 106.200 65.400 ;
                RECT 140.560 65.080 159.240 65.400 ;
                RECT 260.920 65.080 267.680 65.400 ;
                RECT 2.880 66.440 75.600 66.760 ;
                RECT 78.000 66.440 106.200 66.760 ;
                RECT 143.280 66.440 159.240 66.760 ;
                RECT 260.920 66.440 267.680 66.760 ;
                RECT 2.880 67.800 106.200 68.120 ;
                RECT 141.920 67.800 159.240 68.120 ;
                RECT 260.920 67.800 267.680 68.120 ;
                RECT 2.880 69.160 76.280 69.480 ;
                RECT 84.800 69.160 106.200 69.480 ;
                RECT 143.280 69.160 159.240 69.480 ;
                RECT 260.920 69.160 267.680 69.480 ;
                RECT 2.880 70.520 72.880 70.840 ;
                RECT 78.000 70.520 106.200 70.840 ;
                RECT 131.040 70.520 159.240 70.840 ;
                RECT 260.920 70.520 267.680 70.840 ;
                RECT 2.880 71.880 75.600 72.200 ;
                RECT 78.000 71.880 106.200 72.200 ;
                RECT 146.000 71.880 159.240 72.200 ;
                RECT 260.920 71.880 267.680 72.200 ;
                RECT 2.880 73.240 106.200 73.560 ;
                RECT 146.000 73.240 159.240 73.560 ;
                RECT 260.920 73.240 267.680 73.560 ;
                RECT 2.880 74.600 66.760 74.920 ;
                RECT 89.560 74.600 106.200 74.920 ;
                RECT 144.640 74.600 159.240 74.920 ;
                RECT 260.920 74.600 267.680 74.920 ;
                RECT 2.880 75.960 85.120 76.280 ;
                RECT 90.920 75.960 106.200 76.280 ;
                RECT 148.720 75.960 159.240 76.280 ;
                RECT 260.920 75.960 267.680 76.280 ;
                RECT 2.880 77.320 75.600 77.640 ;
                RECT 78.000 77.320 87.840 77.640 ;
                RECT 91.600 77.320 106.200 77.640 ;
                RECT 148.720 77.320 159.240 77.640 ;
                RECT 260.920 77.320 267.680 77.640 ;
                RECT 2.880 78.680 67.440 79.000 ;
                RECT 80.720 78.680 106.200 79.000 ;
                RECT 131.040 78.680 159.240 79.000 ;
                RECT 260.920 78.680 267.680 79.000 ;
                RECT 2.880 80.040 75.600 80.360 ;
                RECT 84.800 80.040 106.200 80.360 ;
                RECT 151.440 80.040 159.240 80.360 ;
                RECT 260.920 80.040 267.680 80.360 ;
                RECT 2.880 81.400 73.560 81.720 ;
                RECT 84.800 81.400 106.200 81.720 ;
                RECT 131.040 81.400 159.240 81.720 ;
                RECT 260.920 81.400 267.680 81.720 ;
                RECT 2.880 82.760 68.800 83.080 ;
                RECT 75.280 82.760 106.200 83.080 ;
                RECT 150.080 82.760 159.240 83.080 ;
                RECT 260.920 82.760 267.680 83.080 ;
                RECT 2.880 84.120 106.200 84.440 ;
                RECT 154.160 84.120 159.240 84.440 ;
                RECT 260.920 84.120 267.680 84.440 ;
                RECT 2.880 85.480 68.800 85.800 ;
                RECT 71.880 85.480 106.200 85.800 ;
                RECT 154.160 85.480 159.240 85.800 ;
                RECT 260.920 85.480 267.680 85.800 ;
                RECT 2.880 86.840 68.800 87.160 ;
                RECT 78.000 86.840 106.200 87.160 ;
                RECT 152.800 86.840 159.240 87.160 ;
                RECT 260.920 86.840 267.680 87.160 ;
                RECT 2.880 88.200 72.880 88.520 ;
                RECT 83.440 88.200 106.200 88.520 ;
                RECT 156.880 88.200 159.240 88.520 ;
                RECT 260.920 88.200 267.680 88.520 ;
                RECT 2.880 89.560 75.600 89.880 ;
                RECT 77.320 89.560 106.200 89.880 ;
                RECT 155.520 89.560 159.240 89.880 ;
                RECT 260.920 89.560 267.680 89.880 ;
                RECT 2.880 90.920 76.280 91.240 ;
                RECT 78.680 90.920 106.200 91.240 ;
                RECT 156.880 90.920 159.240 91.240 ;
                RECT 260.920 90.920 267.680 91.240 ;
                RECT 2.880 92.280 106.200 92.600 ;
                RECT 260.920 92.280 267.680 92.600 ;
                RECT 2.880 93.640 67.440 93.960 ;
                RECT 77.320 93.640 106.200 93.960 ;
                RECT 260.920 93.640 267.680 93.960 ;
                RECT 2.880 95.000 67.440 95.320 ;
                RECT 84.800 95.000 106.200 95.320 ;
                RECT 260.920 95.000 267.680 95.320 ;
                RECT 2.880 96.360 75.600 96.680 ;
                RECT 78.680 96.360 106.200 96.680 ;
                RECT 131.040 96.360 159.240 96.680 ;
                RECT 260.920 96.360 267.680 96.680 ;
                RECT 2.880 97.720 82.400 98.040 ;
                RECT 84.800 97.720 159.240 98.040 ;
                RECT 260.920 97.720 267.680 98.040 ;
                RECT 2.880 99.080 134.760 99.400 ;
                RECT 260.920 99.080 267.680 99.400 ;
                RECT 2.880 100.440 63.360 100.760 ;
                RECT 77.320 100.440 156.520 100.760 ;
                RECT 260.920 100.440 267.680 100.760 ;
                RECT 2.880 101.800 45.680 102.120 ;
                RECT 63.720 101.800 73.560 102.120 ;
                RECT 80.720 101.800 153.800 102.120 ;
                RECT 260.920 101.800 267.680 102.120 ;
                RECT 2.880 103.160 45.680 103.480 ;
                RECT 63.720 103.160 151.080 103.480 ;
                RECT 260.920 103.160 267.680 103.480 ;
                RECT 2.880 104.520 45.680 104.840 ;
                RECT 63.720 104.520 148.360 104.840 ;
                RECT 260.920 104.520 267.680 104.840 ;
                RECT 2.880 105.880 45.680 106.200 ;
                RECT 63.720 105.880 79.000 106.200 ;
                RECT 86.840 105.880 145.640 106.200 ;
                RECT 260.920 105.880 267.680 106.200 ;
                RECT 2.880 107.240 45.680 107.560 ;
                RECT 63.720 107.240 142.920 107.560 ;
                RECT 260.920 107.240 267.680 107.560 ;
                RECT 2.880 108.600 45.680 108.920 ;
                RECT 63.720 108.600 72.200 108.920 ;
                RECT 84.800 108.600 140.200 108.920 ;
                RECT 260.920 108.600 267.680 108.920 ;
                RECT 2.880 109.960 45.680 110.280 ;
                RECT 63.720 109.960 68.800 110.280 ;
                RECT 71.880 109.960 137.480 110.280 ;
                RECT 260.920 109.960 267.680 110.280 ;
                RECT 2.880 111.320 45.680 111.640 ;
                RECT 63.720 111.320 66.760 111.640 ;
                RECT 70.520 111.320 159.240 111.640 ;
                RECT 260.920 111.320 267.680 111.640 ;
                RECT 2.880 112.680 45.680 113.000 ;
                RECT 63.720 112.680 159.240 113.000 ;
                RECT 260.920 112.680 267.680 113.000 ;
                RECT 2.880 114.040 45.680 114.360 ;
                RECT 63.720 114.040 159.240 114.360 ;
                RECT 260.920 114.040 267.680 114.360 ;
                RECT 2.880 115.400 45.680 115.720 ;
                RECT 63.720 115.400 159.240 115.720 ;
                RECT 260.920 115.400 267.680 115.720 ;
                RECT 2.880 116.760 45.680 117.080 ;
                RECT 64.400 116.760 82.400 117.080 ;
                RECT 84.800 116.760 159.240 117.080 ;
                RECT 260.920 116.760 267.680 117.080 ;
                RECT 2.880 118.120 45.680 118.440 ;
                RECT 63.720 118.120 90.560 118.440 ;
                RECT 131.040 118.120 159.240 118.440 ;
                RECT 260.920 118.120 267.680 118.440 ;
                RECT 2.880 119.480 45.680 119.800 ;
                RECT 63.720 119.480 68.800 119.800 ;
                RECT 73.920 119.480 125.240 119.800 ;
                RECT 131.040 119.480 159.240 119.800 ;
                RECT 260.920 119.480 267.680 119.800 ;
                RECT 2.880 120.840 45.680 121.160 ;
                RECT 63.720 120.840 125.240 121.160 ;
                RECT 131.040 120.840 159.240 121.160 ;
                RECT 260.920 120.840 267.680 121.160 ;
                RECT 2.880 122.200 45.680 122.520 ;
                RECT 63.720 122.200 125.240 122.520 ;
                RECT 131.040 122.200 159.240 122.520 ;
                RECT 260.920 122.200 267.680 122.520 ;
                RECT 2.880 123.560 45.680 123.880 ;
                RECT 63.720 123.560 159.240 123.880 ;
                RECT 260.920 123.560 267.680 123.880 ;
                RECT 2.880 124.920 45.680 125.240 ;
                RECT 63.720 124.920 71.520 125.240 ;
                RECT 74.600 124.920 138.840 125.240 ;
                RECT 260.920 124.920 267.680 125.240 ;
                RECT 2.880 126.280 45.680 126.600 ;
                RECT 63.720 126.280 68.800 126.600 ;
                RECT 84.120 126.280 138.840 126.600 ;
                RECT 260.920 126.280 267.680 126.600 ;
                RECT 2.880 127.640 45.680 127.960 ;
                RECT 63.720 127.640 141.560 127.960 ;
                RECT 260.920 127.640 267.680 127.960 ;
                RECT 2.880 129.000 45.680 129.320 ;
                RECT 63.720 129.000 108.240 129.320 ;
                RECT 130.360 129.000 144.280 129.320 ;
                RECT 260.920 129.000 267.680 129.320 ;
                RECT 2.880 130.360 45.680 130.680 ;
                RECT 63.720 130.360 108.240 130.680 ;
                RECT 130.360 130.360 149.720 130.680 ;
                RECT 260.920 130.360 267.680 130.680 ;
                RECT 2.880 131.720 45.680 132.040 ;
                RECT 63.720 131.720 108.240 132.040 ;
                RECT 130.360 131.720 152.440 132.040 ;
                RECT 260.920 131.720 267.680 132.040 ;
                RECT 2.880 133.080 45.680 133.400 ;
                RECT 63.720 133.080 108.240 133.400 ;
                RECT 130.360 133.080 155.160 133.400 ;
                RECT 260.920 133.080 267.680 133.400 ;
                RECT 2.880 134.440 45.680 134.760 ;
                RECT 63.720 134.440 108.240 134.760 ;
                RECT 130.360 134.440 157.880 134.760 ;
                RECT 260.920 134.440 267.680 134.760 ;
                RECT 2.880 135.800 70.160 136.120 ;
                RECT 74.600 135.800 108.240 136.120 ;
                RECT 260.920 135.800 267.680 136.120 ;
                RECT 2.880 137.160 108.240 137.480 ;
                RECT 130.360 137.160 159.240 137.480 ;
                RECT 260.920 137.160 267.680 137.480 ;
                RECT 2.880 138.520 108.240 138.840 ;
                RECT 130.360 138.520 159.240 138.840 ;
                RECT 260.920 138.520 267.680 138.840 ;
                RECT 2.880 139.880 26.640 140.200 ;
                RECT 45.360 139.880 108.240 140.200 ;
                RECT 130.360 139.880 159.240 140.200 ;
                RECT 260.920 139.880 267.680 140.200 ;
                RECT 2.880 141.240 26.640 141.560 ;
                RECT 45.360 141.240 72.880 141.560 ;
                RECT 78.680 141.240 108.240 141.560 ;
                RECT 130.360 141.240 159.240 141.560 ;
                RECT 260.920 141.240 267.680 141.560 ;
                RECT 2.880 142.600 26.640 142.920 ;
                RECT 45.360 142.600 51.120 142.920 ;
                RECT 58.960 142.600 108.240 142.920 ;
                RECT 130.360 142.600 159.240 142.920 ;
                RECT 260.920 142.600 267.680 142.920 ;
                RECT 2.880 143.960 26.640 144.280 ;
                RECT 63.040 143.960 108.240 144.280 ;
                RECT 130.360 143.960 159.240 144.280 ;
                RECT 260.920 143.960 267.680 144.280 ;
                RECT 2.880 145.320 26.640 145.640 ;
                RECT 45.360 145.320 108.240 145.640 ;
                RECT 260.920 145.320 267.680 145.640 ;
                RECT 2.880 146.680 18.480 147.000 ;
                RECT 58.960 146.680 67.440 147.000 ;
                RECT 77.320 146.680 108.240 147.000 ;
                RECT 130.360 146.680 159.240 147.000 ;
                RECT 260.920 146.680 267.680 147.000 ;
                RECT 2.880 148.040 51.120 148.360 ;
                RECT 71.880 148.040 267.680 148.360 ;
                RECT 2.880 149.400 66.760 149.720 ;
                RECT 70.520 149.400 267.680 149.720 ;
                RECT 2.880 150.760 156.520 151.080 ;
                RECT 263.640 150.760 267.680 151.080 ;
                RECT 2.880 152.120 156.520 152.440 ;
                RECT 263.640 152.120 267.680 152.440 ;
                RECT 2.880 153.480 62.000 153.800 ;
                RECT 68.480 153.480 115.720 153.800 ;
                RECT 263.640 153.480 267.680 153.800 ;
                RECT 2.880 154.840 59.960 155.160 ;
                RECT 82.080 154.840 115.720 155.160 ;
                RECT 263.640 154.840 267.680 155.160 ;
                RECT 2.880 156.200 59.960 156.520 ;
                RECT 81.400 156.200 95.320 156.520 ;
                RECT 105.200 156.200 115.720 156.520 ;
                RECT 263.640 156.200 267.680 156.520 ;
                RECT 2.880 157.560 73.560 157.880 ;
                RECT 80.720 157.560 95.320 157.880 ;
                RECT 105.200 157.560 115.720 157.880 ;
                RECT 263.640 157.560 267.680 157.880 ;
                RECT 2.880 158.920 59.960 159.240 ;
                RECT 70.520 158.920 95.320 159.240 ;
                RECT 105.200 158.920 115.720 159.240 ;
                RECT 263.640 158.920 267.680 159.240 ;
                RECT 2.880 160.280 59.960 160.600 ;
                RECT 70.520 160.280 95.320 160.600 ;
                RECT 105.200 160.280 115.720 160.600 ;
                RECT 263.640 160.280 267.680 160.600 ;
                RECT 2.880 161.640 59.960 161.960 ;
                RECT 70.520 161.640 95.320 161.960 ;
                RECT 105.200 161.640 115.720 161.960 ;
                RECT 263.640 161.640 267.680 161.960 ;
                RECT 2.880 163.000 59.960 163.320 ;
                RECT 70.520 163.000 115.720 163.320 ;
                RECT 263.640 163.000 267.680 163.320 ;
                RECT 2.880 164.360 95.320 164.680 ;
                RECT 105.200 164.360 115.720 164.680 ;
                RECT 263.640 164.360 267.680 164.680 ;
                RECT 2.880 165.720 95.320 166.040 ;
                RECT 105.200 165.720 115.720 166.040 ;
                RECT 263.640 165.720 267.680 166.040 ;
                RECT 2.880 167.080 18.480 167.400 ;
                RECT 55.560 167.080 95.320 167.400 ;
                RECT 105.200 167.080 115.720 167.400 ;
                RECT 263.640 167.080 267.680 167.400 ;
                RECT 2.880 168.440 17.800 168.760 ;
                RECT 55.560 168.440 95.320 168.760 ;
                RECT 105.200 168.440 115.720 168.760 ;
                RECT 263.640 168.440 267.680 168.760 ;
                RECT 2.880 169.800 95.320 170.120 ;
                RECT 102.480 169.800 115.720 170.120 ;
                RECT 263.640 169.800 267.680 170.120 ;
                RECT 2.880 171.160 17.120 171.480 ;
                RECT 55.560 171.160 68.800 171.480 ;
                RECT 72.560 171.160 99.400 171.480 ;
                RECT 105.200 171.160 115.720 171.480 ;
                RECT 263.640 171.160 267.680 171.480 ;
                RECT 2.880 172.520 16.440 172.840 ;
                RECT 55.560 172.520 68.800 172.840 ;
                RECT 73.240 172.520 95.320 172.840 ;
                RECT 105.200 172.520 115.720 172.840 ;
                RECT 263.640 172.520 267.680 172.840 ;
                RECT 2.880 173.880 95.320 174.200 ;
                RECT 105.200 173.880 115.720 174.200 ;
                RECT 263.640 173.880 267.680 174.200 ;
                RECT 2.880 175.240 15.760 175.560 ;
                RECT 55.560 175.240 68.800 175.560 ;
                RECT 73.920 175.240 95.320 175.560 ;
                RECT 105.200 175.240 115.720 175.560 ;
                RECT 263.640 175.240 267.680 175.560 ;
                RECT 2.880 176.600 15.080 176.920 ;
                RECT 55.560 176.600 68.800 176.920 ;
                RECT 74.600 176.600 95.320 176.920 ;
                RECT 105.200 176.600 115.720 176.920 ;
                RECT 263.640 176.600 267.680 176.920 ;
                RECT 2.880 177.960 14.400 178.280 ;
                RECT 55.560 177.960 68.800 178.280 ;
                RECT 74.600 177.960 95.320 178.280 ;
                RECT 103.840 177.960 115.720 178.280 ;
                RECT 263.640 177.960 267.680 178.280 ;
                RECT 2.880 179.320 13.720 179.640 ;
                RECT 55.560 179.320 101.440 179.640 ;
                RECT 105.200 179.320 115.720 179.640 ;
                RECT 263.640 179.320 267.680 179.640 ;
                RECT 2.880 180.680 95.320 181.000 ;
                RECT 105.200 180.680 115.720 181.000 ;
                RECT 263.640 180.680 267.680 181.000 ;
                RECT 2.880 182.040 13.040 182.360 ;
                RECT 55.560 182.040 95.320 182.360 ;
                RECT 105.200 182.040 115.720 182.360 ;
                RECT 263.640 182.040 267.680 182.360 ;
                RECT 2.880 183.400 12.360 183.720 ;
                RECT 55.560 183.400 95.320 183.720 ;
                RECT 105.200 183.400 115.720 183.720 ;
                RECT 263.640 183.400 267.680 183.720 ;
                RECT 2.880 184.760 11.680 185.080 ;
                RECT 55.560 184.760 95.320 185.080 ;
                RECT 105.200 184.760 115.720 185.080 ;
                RECT 263.640 184.760 267.680 185.080 ;
                RECT 2.880 186.120 115.720 186.440 ;
                RECT 263.640 186.120 267.680 186.440 ;
                RECT 2.880 187.480 11.000 187.800 ;
                RECT 55.560 187.480 68.800 187.800 ;
                RECT 71.200 187.480 96.680 187.800 ;
                RECT 105.200 187.480 115.720 187.800 ;
                RECT 263.640 187.480 267.680 187.800 ;
                RECT 2.880 188.840 100.080 189.160 ;
                RECT 105.200 188.840 115.720 189.160 ;
                RECT 263.640 188.840 267.680 189.160 ;
                RECT 2.880 190.200 100.080 190.520 ;
                RECT 105.200 190.200 115.720 190.520 ;
                RECT 263.640 190.200 267.680 190.520 ;
                RECT 2.880 191.560 96.680 191.880 ;
                RECT 105.200 191.560 115.720 191.880 ;
                RECT 263.640 191.560 267.680 191.880 ;
                RECT 2.880 192.920 96.680 193.240 ;
                RECT 105.200 192.920 115.720 193.240 ;
                RECT 263.640 192.920 267.680 193.240 ;
                RECT 2.880 194.280 72.880 194.600 ;
                RECT 82.080 194.280 115.720 194.600 ;
                RECT 263.640 194.280 267.680 194.600 ;
                RECT 2.880 195.640 71.520 195.960 ;
                RECT 81.400 195.640 96.680 195.960 ;
                RECT 105.200 195.640 115.720 195.960 ;
                RECT 263.640 195.640 267.680 195.960 ;
                RECT 2.880 197.000 70.160 197.320 ;
                RECT 80.720 197.000 95.320 197.320 ;
                RECT 105.200 197.000 115.720 197.320 ;
                RECT 263.640 197.000 267.680 197.320 ;
                RECT 2.880 198.360 95.320 198.680 ;
                RECT 105.200 198.360 115.720 198.680 ;
                RECT 263.640 198.360 267.680 198.680 ;
                RECT 2.880 199.720 95.320 200.040 ;
                RECT 105.200 199.720 115.720 200.040 ;
                RECT 263.640 199.720 267.680 200.040 ;
                RECT 2.880 201.080 95.320 201.400 ;
                RECT 105.200 201.080 115.720 201.400 ;
                RECT 263.640 201.080 267.680 201.400 ;
                RECT 2.880 202.440 115.720 202.760 ;
                RECT 263.640 202.440 267.680 202.760 ;
                RECT 2.880 203.800 95.320 204.120 ;
                RECT 105.200 203.800 115.720 204.120 ;
                RECT 263.640 203.800 267.680 204.120 ;
                RECT 2.880 205.160 95.320 205.480 ;
                RECT 105.200 205.160 115.720 205.480 ;
                RECT 263.640 205.160 267.680 205.480 ;
                RECT 2.880 206.520 95.320 206.840 ;
                RECT 105.200 206.520 115.720 206.840 ;
                RECT 263.640 206.520 267.680 206.840 ;
                RECT 2.880 207.880 95.320 208.200 ;
                RECT 105.200 207.880 115.720 208.200 ;
                RECT 263.640 207.880 267.680 208.200 ;
                RECT 2.880 209.240 95.320 209.560 ;
                RECT 98.400 209.240 115.720 209.560 ;
                RECT 263.640 209.240 267.680 209.560 ;
                RECT 2.880 210.600 101.440 210.920 ;
                RECT 105.200 210.600 115.720 210.920 ;
                RECT 263.640 210.600 267.680 210.920 ;
                RECT 2.880 211.960 95.320 212.280 ;
                RECT 105.200 211.960 115.720 212.280 ;
                RECT 263.640 211.960 267.680 212.280 ;
                RECT 2.880 213.320 95.320 213.640 ;
                RECT 105.200 213.320 115.720 213.640 ;
                RECT 263.640 213.320 267.680 213.640 ;
                RECT 2.880 214.680 95.320 215.000 ;
                RECT 105.200 214.680 115.720 215.000 ;
                RECT 263.640 214.680 267.680 215.000 ;
                RECT 2.880 216.040 95.320 216.360 ;
                RECT 105.200 216.040 115.720 216.360 ;
                RECT 263.640 216.040 267.680 216.360 ;
                RECT 2.880 217.400 95.320 217.720 ;
                RECT 99.760 217.400 115.720 217.720 ;
                RECT 263.640 217.400 267.680 217.720 ;
                RECT 2.880 218.760 99.400 219.080 ;
                RECT 105.200 218.760 115.720 219.080 ;
                RECT 263.640 218.760 267.680 219.080 ;
                RECT 2.880 220.120 95.320 220.440 ;
                RECT 105.200 220.120 115.720 220.440 ;
                RECT 263.640 220.120 267.680 220.440 ;
                RECT 2.880 221.480 95.320 221.800 ;
                RECT 105.200 221.480 115.720 221.800 ;
                RECT 263.640 221.480 267.680 221.800 ;
                RECT 2.880 222.840 95.320 223.160 ;
                RECT 105.200 222.840 115.720 223.160 ;
                RECT 263.640 222.840 267.680 223.160 ;
                RECT 2.880 224.200 95.320 224.520 ;
                RECT 105.200 224.200 115.720 224.520 ;
                RECT 263.640 224.200 267.680 224.520 ;
                RECT 2.880 225.560 115.720 225.880 ;
                RECT 263.640 225.560 267.680 225.880 ;
                RECT 2.880 226.920 97.360 227.240 ;
                RECT 105.200 226.920 115.720 227.240 ;
                RECT 263.640 226.920 267.680 227.240 ;
                RECT 2.880 228.280 102.120 228.600 ;
                RECT 105.200 228.280 115.720 228.600 ;
                RECT 263.640 228.280 267.680 228.600 ;
                RECT 2.880 229.640 97.360 229.960 ;
                RECT 105.200 229.640 115.720 229.960 ;
                RECT 263.640 229.640 267.680 229.960 ;
                RECT 2.880 231.000 97.360 231.320 ;
                RECT 105.200 231.000 115.720 231.320 ;
                RECT 263.640 231.000 267.680 231.320 ;
                RECT 2.880 232.360 97.360 232.680 ;
                RECT 105.200 232.360 115.720 232.680 ;
                RECT 263.640 232.360 267.680 232.680 ;
                RECT 2.880 233.720 115.720 234.040 ;
                RECT 263.640 233.720 267.680 234.040 ;
                RECT 2.880 235.080 98.040 235.400 ;
                RECT 105.200 235.080 115.720 235.400 ;
                RECT 263.640 235.080 267.680 235.400 ;
                RECT 2.880 236.440 98.040 236.760 ;
                RECT 105.200 236.440 115.720 236.760 ;
                RECT 263.640 236.440 267.680 236.760 ;
                RECT 2.880 237.800 100.080 238.120 ;
                RECT 105.200 237.800 115.720 238.120 ;
                RECT 263.640 237.800 267.680 238.120 ;
                RECT 2.880 239.160 100.760 239.480 ;
                RECT 105.200 239.160 115.720 239.480 ;
                RECT 263.640 239.160 267.680 239.480 ;
                RECT 2.880 240.520 98.040 240.840 ;
                RECT 105.200 240.520 115.720 240.840 ;
                RECT 263.640 240.520 267.680 240.840 ;
                RECT 2.880 241.880 115.720 242.200 ;
                RECT 263.640 241.880 267.680 242.200 ;
                RECT 2.880 243.240 98.040 243.560 ;
                RECT 105.200 243.240 115.720 243.560 ;
                RECT 263.640 243.240 267.680 243.560 ;
                RECT 2.880 244.600 98.040 244.920 ;
                RECT 105.200 244.600 115.720 244.920 ;
                RECT 263.640 244.600 267.680 244.920 ;
                RECT 2.880 245.960 98.040 246.280 ;
                RECT 105.200 245.960 115.720 246.280 ;
                RECT 263.640 245.960 267.680 246.280 ;
                RECT 2.880 247.320 98.040 247.640 ;
                RECT 105.200 247.320 115.720 247.640 ;
                RECT 263.640 247.320 267.680 247.640 ;
                RECT 2.880 248.680 115.720 249.000 ;
                RECT 263.640 248.680 267.680 249.000 ;
                RECT 2.880 250.040 99.400 250.360 ;
                RECT 105.200 250.040 115.720 250.360 ;
                RECT 263.640 250.040 267.680 250.360 ;
                RECT 2.880 251.400 98.720 251.720 ;
                RECT 105.200 251.400 115.720 251.720 ;
                RECT 263.640 251.400 267.680 251.720 ;
                RECT 2.880 252.760 98.720 253.080 ;
                RECT 105.200 252.760 115.720 253.080 ;
                RECT 263.640 252.760 267.680 253.080 ;
                RECT 2.880 254.120 98.720 254.440 ;
                RECT 105.200 254.120 115.720 254.440 ;
                RECT 263.640 254.120 267.680 254.440 ;
                RECT 2.880 255.480 98.720 255.800 ;
                RECT 105.200 255.480 115.720 255.800 ;
                RECT 263.640 255.480 267.680 255.800 ;
                RECT 2.880 256.840 115.720 257.160 ;
                RECT 263.640 256.840 267.680 257.160 ;
                RECT 2.880 258.200 101.440 258.520 ;
                RECT 105.200 258.200 115.720 258.520 ;
                RECT 263.640 258.200 267.680 258.520 ;
                RECT 2.880 259.560 98.720 259.880 ;
                RECT 105.200 259.560 115.720 259.880 ;
                RECT 263.640 259.560 267.680 259.880 ;
                RECT 2.880 260.920 98.720 261.240 ;
                RECT 105.200 260.920 115.720 261.240 ;
                RECT 263.640 260.920 267.680 261.240 ;
                RECT 2.880 262.280 98.720 262.600 ;
                RECT 105.200 262.280 115.720 262.600 ;
                RECT 263.640 262.280 267.680 262.600 ;
                RECT 2.880 263.640 98.720 263.960 ;
                RECT 105.200 263.640 115.720 263.960 ;
                RECT 263.640 263.640 267.680 263.960 ;
                RECT 2.880 265.000 115.720 265.320 ;
                RECT 263.640 265.000 267.680 265.320 ;
                RECT 2.880 266.360 98.720 266.680 ;
                RECT 105.200 266.360 115.720 266.680 ;
                RECT 263.640 266.360 267.680 266.680 ;
                RECT 2.880 267.720 100.080 268.040 ;
                RECT 105.200 267.720 115.720 268.040 ;
                RECT 263.640 267.720 267.680 268.040 ;
                RECT 2.880 269.080 98.720 269.400 ;
                RECT 105.200 269.080 115.720 269.400 ;
                RECT 263.640 269.080 267.680 269.400 ;
                RECT 2.880 270.440 98.720 270.760 ;
                RECT 105.200 270.440 115.720 270.760 ;
                RECT 263.640 270.440 267.680 270.760 ;
                RECT 2.880 271.800 98.720 272.120 ;
                RECT 105.200 271.800 115.720 272.120 ;
                RECT 263.640 271.800 267.680 272.120 ;
                RECT 2.880 273.160 115.720 273.480 ;
                RECT 263.640 273.160 267.680 273.480 ;
                RECT 2.880 274.520 98.720 274.840 ;
                RECT 105.200 274.520 115.720 274.840 ;
                RECT 263.640 274.520 267.680 274.840 ;
                RECT 2.880 275.880 98.720 276.200 ;
                RECT 105.200 275.880 115.720 276.200 ;
                RECT 263.640 275.880 267.680 276.200 ;
                RECT 2.880 277.240 102.120 277.560 ;
                RECT 105.200 277.240 115.720 277.560 ;
                RECT 263.640 277.240 267.680 277.560 ;
                RECT 2.880 278.600 98.720 278.920 ;
                RECT 105.200 278.600 115.720 278.920 ;
                RECT 263.640 278.600 267.680 278.920 ;
                RECT 2.880 279.960 98.720 280.280 ;
                RECT 105.200 279.960 115.720 280.280 ;
                RECT 263.640 279.960 267.680 280.280 ;
                RECT 2.880 281.320 115.720 281.640 ;
                RECT 263.640 281.320 267.680 281.640 ;
                RECT 2.880 282.680 156.520 283.000 ;
                RECT 263.640 282.680 267.680 283.000 ;
                RECT 2.880 284.040 156.520 284.360 ;
                RECT 263.640 284.040 267.680 284.360 ;
                RECT 2.880 285.400 156.520 285.720 ;
                RECT 263.640 285.400 267.680 285.720 ;
                RECT 2.880 286.760 267.680 287.080 ;
                RECT 2.880 288.120 267.680 288.440 ;
                RECT 2.880 289.480 267.680 289.800 ;
                RECT 2.880 290.840 267.680 291.160 ;
                RECT 2.880 2.880 267.680 4.240 ;
                RECT 2.880 292.840 267.680 294.200 ;
                RECT 160.660 29.370 166.460 30.490 ;
                RECT 253.360 29.370 259.160 30.490 ;
                RECT 160.660 35.070 166.460 35.520 ;
                RECT 253.360 35.070 259.160 35.520 ;
                RECT 160.660 38.950 166.460 39.510 ;
                RECT 253.360 38.950 259.160 39.510 ;
                RECT 160.660 43.550 166.460 44.110 ;
                RECT 253.360 43.550 259.160 44.110 ;
                RECT 160.660 56.840 259.160 58.640 ;
                RECT 160.660 68.900 259.160 69.700 ;
                RECT 160.660 77.030 259.160 79.120 ;
                RECT 160.660 65.890 259.160 66.690 ;
                RECT 160.660 121.410 259.160 122.815 ;
                RECT 160.660 73.790 259.160 74.590 ;
                RECT 160.660 98.135 259.160 98.425 ;
                RECT 160.660 70.580 259.160 71.380 ;
                RECT 160.660 20.000 259.160 21.800 ;
                RECT 116.500 153.875 118.250 281.855 ;
                RECT 129.855 153.875 131.775 281.855 ;
                RECT 133.695 153.875 135.615 281.855 ;
                RECT 106.610 61.175 107.500 96.575 ;
                RECT 113.370 61.175 114.260 96.575 ;
                RECT 120.560 61.175 122.310 96.575 ;
                RECT 108.845 129.020 109.955 147.240 ;
                RECT 117.220 129.020 118.110 147.240 ;
                RECT 123.765 129.020 125.085 147.240 ;
                RECT 126.130 117.860 127.020 123.020 ;
                RECT 126.560 50.015 127.450 55.175 ;
                RECT 60.480 154.940 69.640 155.310 ;
                RECT 60.480 158.275 69.640 159.165 ;
                RECT 27.420 139.250 44.660 139.920 ;
                RECT 27.420 140.610 44.660 142.300 ;
        END 
    END vss 
    OBS 
        LAYER met1 ;
            RECT 0.000 0.000 270.560 297.080 ;
        LAYER met2 ;
            RECT 0.000 0.000 270.560 297.080 ;
    END 
END sram22_512x8m8w1 
END LIBRARY 

