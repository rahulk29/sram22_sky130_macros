VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sramgen_sram_4096x32m8w8_replica_v1
  CLASS BLOCK ;
  ORIGIN 93.555 1025.97 ;
  FOREIGN sramgen_sram_4096x32m8w8_replica_v1 -93.555 -1025.97 ;
  SIZE 756.015 BY 1037.685 ;
  SYMMETRY X Y R90 ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT -88.2 -1025.57 -87.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -86.6 -1025.57 -86.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -85 -1025.57 -84.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -83.4 -1025.57 -83 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -81.8 -993.54 -81.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -80.2 -1012.62 -79.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -78.6 -1025.57 -78.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -77 -1007.32 -76.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -77 -1025.57 -76.6 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -75.4 -1008.38 -75 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -73.8 -1012.62 -73.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -73.8 -1025.57 -73.4 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -72.2 -1025.57 -71.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -70.6 -1006.26 -70.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -70.6 -1025.57 -70.2 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -69 -1012.62 -68.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -67.4 -1012.62 -67 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -67.4 -1025.57 -67 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -65.8 -1025.57 -65.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -64.2 -1006.26 -63.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -64.2 -1025.57 -63.8 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -62.6 -1012.62 -62.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -61 -1025.57 -60.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -59.4 -1004.14 -59 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -59.4 -1025.57 -59 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -57.8 -1012.62 -57.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -56.2 -1012.62 -55.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -56.2 -1025.57 -55.8 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -54.6 -1025.57 -54.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -53 -1003.08 -52.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -53 -1025.57 -52.6 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -51.4 -1012.62 -51 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.8 -1012.62 -49.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.8 -1025.57 -49.4 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -48.2 -1025.57 -47.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -46.6 -1003.08 -46.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -46.6 -1025.57 -46.2 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -45 -1012.62 -44.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -45 -1025.57 -44.6 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.4 -1025.57 -43 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -41.8 -1002.02 -41.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -41.8 -1025.57 -41.4 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -40.2 -1012.62 -39.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.6 -1012.62 -38.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.6 -1025.57 -38.2 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -37 -1025.57 -36.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -35.4 -1000.96 -35 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -35.4 -1025.57 -35 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -33.8 -1012.62 -33.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -32.2 -1025.57 -31.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.6 -999.9 -30.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.6 -1025.57 -30.2 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -29 -999.9 -28.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -29 -1025.57 -28.6 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -27.4 -1012.62 -27 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -27.4 -1025.57 -27 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -25.8 -1025.57 -25.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -24.2 -998.84 -23.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -24.2 -1025.57 -23.8 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -22.6 -1012.62 -22.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -21 -1012.62 -20.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -21 -1025.57 -20.6 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.4 -1025.57 -19 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.8 -997.78 -17.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.8 -1025.57 -17.4 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -16.2 -1012.62 -15.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -14.6 -1025.57 -14.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -13 -996.72 -12.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -13 -1025.57 -12.6 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.4 -996.72 -11 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.4 -1025.57 -11 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.8 -818.64 -9.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.8 -1012.62 -9.4 -975.94 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.8 -1025.57 -9.4 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -8.2 -1025.57 -7.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -6.6 -992.48 -6.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -6.6 -1025.57 -6.2 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -5 -1025.57 -4.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -3.4 -1025.57 -3 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.8 2.86 -1.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.8 -1025.57 -1.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.2 2.86 0.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.2 -1025.57 0.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.4 2.86 1.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.4 -1025.57 1.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 3 2.86 3.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 3 -1025.57 3.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.6 2.86 5 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.6 -1025.57 5 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.2 2.86 6.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.2 -1025.57 6.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.8 2.86 8.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.8 -1025.57 8.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.4 2.86 9.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.4 -1025.57 9.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 11 2.86 11.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 11 -865.28 11.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 11 -1025.57 11.4 -973.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.6 2.86 13 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.6 -828.18 13 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.6 -902.38 13 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.2 2.86 14.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.2 -839.84 14.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.2 -1025.57 14.6 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.8 2.86 16.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.8 -1025.57 16.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.4 2.86 17.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.4 -1025.57 17.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 19 2.86 19.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 19 -1025.57 19.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.6 2.86 21 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.6 -1025.57 21 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.2 2.86 22.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.2 -907.68 22.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.8 2.86 24.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.8 -907.68 24.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.4 2.86 25.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.4 -1025.57 25.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 27 2.86 27.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 27 -1025.57 27.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.6 2.86 29 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.6 -1025.57 29 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.2 2.86 30.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.2 -1025.57 30.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.8 2.86 32.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.8 -1025.57 32.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.4 2.86 33.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.4 -828.18 33.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.4 -902.38 33.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 35 2.86 35.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 35 -828.18 35.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 35 -1025.57 35.4 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.6 2.86 37 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.6 -844.08 37 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.6 -1025.57 37 -926.12 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.2 2.86 38.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.2 -1025.57 38.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.8 2.86 40.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.8 -1025.57 40.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.4 2.86 41.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.4 -1025.57 41.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 43 2.86 43.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 43 -1025.57 43.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.6 2.86 45 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.6 -1025.57 45 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.2 2.86 46.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.2 -1025.57 46.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.8 2.86 48.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.8 -1025.57 48.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.4 2.86 49.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.4 -1025.57 49.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 51 2.86 51.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 51 -1025.57 51.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.6 2.86 53 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.6 -828.18 53 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.6 -902.38 53 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.2 2.86 54.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.2 -839.84 54.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.2 -1025.57 54.6 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.8 2.86 56.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.8 -1025.57 56.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.4 2.86 57.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.4 -1025.57 57.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 59 2.86 59.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 59 -1025.57 59.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.6 2.86 61 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.6 -1025.57 61 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.2 2.86 62.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.2 -907.68 62.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.8 2.86 64.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.8 -907.68 64.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.8 -1025.57 64.2 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.4 2.86 65.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.4 -1025.57 65.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 67 2.86 67.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 67 -1025.57 67.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.6 2.86 69 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.6 -1025.57 69 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.2 2.86 70.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.2 -1025.57 70.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.8 2.86 72.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.8 -1025.57 72.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.4 2.86 73.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.4 -828.18 73.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.4 -902.38 73.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 75 2.86 75.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 75 -828.18 75.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 75 -1025.57 75.4 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.6 2.86 77 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.6 -1025.57 77 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.2 2.86 78.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.2 -1025.57 78.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.8 2.86 80.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.8 -1025.57 80.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.4 2.86 81.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.4 -1025.57 81.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 83 2.86 83.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 83 -1025.57 83.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.6 2.86 85 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.6 -1025.57 85 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.2 2.86 86.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.2 -1025.57 86.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.8 2.86 88.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.8 -1025.57 88.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.4 2.86 89.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.4 -1025.57 89.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 91 2.86 91.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 91 -1025.57 91.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.6 2.86 93 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.6 -828.18 93 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.6 -902.38 93 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.2 2.86 94.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.2 -839.84 94.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.2 -1025.57 94.6 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.8 2.86 96.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.8 -1025.57 96.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.4 2.86 97.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.4 -1025.57 97.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 99 2.86 99.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 99 -1025.57 99.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.6 2.86 101 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.6 -1025.57 101 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.2 2.86 102.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.2 -907.68 102.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.8 2.86 104.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.8 -907.68 104.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.8 -1025.57 104.2 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.4 2.86 105.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.4 -1025.57 105.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 107 2.86 107.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 107 -1025.57 107.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.6 2.86 109 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.6 -1025.57 109 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.2 2.86 110.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.2 -1025.57 110.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.8 2.86 112.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.8 -1025.57 112.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.4 2.86 113.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.4 -828.18 113.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.4 -902.38 113.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 115 2.86 115.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 115 -828.18 115.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 115 -1025.57 115.4 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.6 2.86 117 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.6 -1025.57 117 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.2 2.86 118.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.2 -1025.57 118.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.8 2.86 120.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.8 -1025.57 120.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.4 2.86 121.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.4 -1025.57 121.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 123 2.86 123.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 123 -1025.57 123.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.6 2.86 125 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.6 -1025.57 125 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.2 2.86 126.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.2 -1025.57 126.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.8 2.86 128.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.8 -1025.57 128.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.4 2.86 129.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.4 -1025.57 129.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 131 2.86 131.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 131 -1025.57 131.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.6 2.86 133 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.6 -828.18 133 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.6 -902.38 133 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.2 2.86 134.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.2 -839.84 134.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.2 -1025.57 134.6 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.8 2.86 136.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.8 -1025.57 136.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.4 2.86 137.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.4 -1025.57 137.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 139 2.86 139.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 139 -1025.57 139.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.6 2.86 141 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.6 -1025.57 141 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.2 2.86 142.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.2 -907.68 142.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.8 2.86 144.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.8 -907.68 144.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.8 -1025.57 144.2 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.4 2.86 145.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.4 -1025.57 145.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 147 2.86 147.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 147 -1025.57 147.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.6 2.86 149 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.6 -1025.57 149 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.2 2.86 150.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.2 -1025.57 150.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.8 2.86 152.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.8 -1025.57 152.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.4 2.86 153.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.4 -828.18 153.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.4 -902.38 153.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 155 2.86 155.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 155 -828.18 155.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 155 -1025.57 155.4 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.6 2.86 157 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.6 -1025.57 157 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.2 2.86 158.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.2 -1025.57 158.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.8 2.86 160.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.8 -1025.57 160.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.4 2.86 161.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.4 -1025.57 161.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 163 2.86 163.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 163 -1025.57 163.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.6 2.86 165 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.6 -1025.57 165 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.2 2.86 166.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.2 -1025.57 166.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.8 2.86 168.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.8 -1025.57 168.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.4 2.86 169.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.4 -1025.57 169.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 171 2.86 171.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 171 -1025.57 171.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.6 2.86 173 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.6 -828.18 173 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.6 -902.38 173 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.2 2.86 174.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.2 -839.84 174.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.2 -1025.57 174.6 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.8 2.86 176.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.8 -1025.57 176.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.4 2.86 177.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.4 -1025.57 177.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 179 2.86 179.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 179 -1025.57 179.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.6 2.86 181 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.6 -1025.57 181 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.2 2.86 182.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.2 -907.68 182.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.8 2.86 184.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.8 -907.68 184.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.4 2.86 185.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.4 -1025.57 185.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 187 2.86 187.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 187 -1025.57 187.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.6 2.86 189 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.6 -1025.57 189 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.2 2.86 190.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.2 -1025.57 190.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 191.8 2.86 192.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 191.8 -1025.57 192.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.4 2.86 193.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.4 -828.18 193.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.4 -902.38 193.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 195 2.86 195.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 195 -828.18 195.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 195 -1025.57 195.4 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.6 2.86 197 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.6 -844.08 197 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.6 -1025.57 197 -926.12 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.2 2.86 198.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.2 -1025.57 198.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.8 2.86 200.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.8 -1025.57 200.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.4 2.86 201.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.4 -1025.57 201.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 203 2.86 203.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 203 -1025.57 203.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.6 2.86 205 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.6 -1025.57 205 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 206.2 2.86 206.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 206.2 -1025.57 206.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.8 2.86 208.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.8 -1025.57 208.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.4 2.86 209.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.4 -1025.57 209.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 211 2.86 211.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 211 -1025.57 211.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 212.6 2.86 213 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 212.6 -828.18 213 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 212.6 -902.38 213 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.2 2.86 214.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.2 -839.84 214.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.2 -1025.57 214.6 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 215.8 2.86 216.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 215.8 -1025.57 216.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 217.4 2.86 217.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 217.4 -1025.57 217.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 219 2.86 219.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 219 -1025.57 219.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.6 2.86 221 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.6 -1025.57 221 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.2 2.86 222.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.2 -907.68 222.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 223.8 2.86 224.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 223.8 -907.68 224.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 223.8 -1025.57 224.2 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 225.4 2.86 225.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 225.4 -1025.57 225.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 227 2.86 227.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 227 -1025.57 227.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.6 2.86 229 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.6 -1025.57 229 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 230.2 2.86 230.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 230.2 -1025.57 230.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.8 2.86 232.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.8 -1025.57 232.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.4 2.86 233.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.4 -828.18 233.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.4 -902.38 233.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 235 2.86 235.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 235 -828.18 235.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 235 -1025.57 235.4 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 236.6 2.86 237 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 236.6 -1025.57 237 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 238.2 2.86 238.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 238.2 -1025.57 238.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.8 2.86 240.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.8 -1025.57 240.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.4 2.86 241.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.4 -1025.57 241.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 243 2.86 243.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 243 -1025.57 243.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 244.6 2.86 245 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 244.6 -1025.57 245 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 246.2 2.86 246.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 246.2 -1025.57 246.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 247.8 2.86 248.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 247.8 -1025.57 248.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.4 2.86 249.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.4 -1025.57 249.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 251 2.86 251.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 251 -1025.57 251.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.6 2.86 253 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.6 -828.18 253 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.6 -902.38 253 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.2 2.86 254.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.2 -839.84 254.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.2 -1025.57 254.6 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 255.8 2.86 256.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 255.8 -1025.57 256.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 257.4 2.86 257.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 257.4 -1025.57 257.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 259 2.86 259.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 259 -1025.57 259.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.6 2.86 261 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.6 -1025.57 261 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.2 2.86 262.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.2 -907.68 262.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 263.8 2.86 264.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 263.8 -907.68 264.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 263.8 -1025.57 264.2 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 265.4 2.86 265.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 265.4 -1025.57 265.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 267 2.86 267.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 267 -1025.57 267.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 268.6 2.86 269 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 268.6 -1025.57 269 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 270.2 2.86 270.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 270.2 -1025.57 270.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.8 2.86 272.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.8 -1025.57 272.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.4 2.86 273.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.4 -828.18 273.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.4 -902.38 273.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 275 2.86 275.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 275 -828.18 275.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 275 -1025.57 275.4 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 276.6 2.86 277 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 276.6 -1025.57 277 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 278.2 2.86 278.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 278.2 -1025.57 278.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.8 2.86 280.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.8 -1025.57 280.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 281.4 2.86 281.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 281.4 -1025.57 281.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 283 2.86 283.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 283 -1025.57 283.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.6 2.86 285 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.6 -1025.57 285 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.2 2.86 286.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.2 -1025.57 286.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 287.8 2.86 288.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 287.8 -1025.57 288.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 289.4 2.86 289.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 289.4 -1025.57 289.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 291 2.86 291.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 291 -1025.57 291.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.6 2.86 293 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.6 -828.18 293 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.6 -902.38 293 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.2 2.86 294.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.2 -839.84 294.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.2 -1025.57 294.6 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 295.8 2.86 296.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 295.8 -1025.57 296.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 297.4 2.86 297.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 297.4 -1025.57 297.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 299 2.86 299.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 299 -1025.57 299.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 300.6 2.86 301 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 300.6 -1025.57 301 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 302.2 2.86 302.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 302.2 -907.68 302.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.8 2.86 304.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.8 -907.68 304.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.8 -1025.57 304.2 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.4 2.86 305.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.4 -1025.57 305.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 307 2.86 307.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 307 -1025.57 307.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 308.6 2.86 309 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 308.6 -1025.57 309 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 310.2 2.86 310.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 310.2 -1025.57 310.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.8 2.86 312.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.8 -1025.57 312.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.4 2.86 313.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.4 -828.18 313.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.4 -902.38 313.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 315 2.86 315.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 315 -828.18 315.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 315 -1025.57 315.4 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.6 2.86 317 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.6 -1025.57 317 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.2 2.86 318.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.2 -1025.57 318.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 319.8 2.86 320.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 319.8 -1025.57 320.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 321.4 2.86 321.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 321.4 -1025.57 321.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 323 2.86 323.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 323 -1025.57 323.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.6 2.86 325 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.6 -1025.57 325 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.2 2.86 326.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.2 -1025.57 326.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 327.8 2.86 328.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 327.8 -1025.57 328.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 329.4 2.86 329.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 329.4 -1025.57 329.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 331 2.86 331.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 331 -1025.57 331.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 332.6 2.86 333 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 332.6 -828.18 333 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 332.6 -902.38 333 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 334.2 2.86 334.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 334.2 -839.84 334.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 334.2 -1025.57 334.6 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.8 2.86 336.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.8 -1025.57 336.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.4 2.86 337.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.4 -1025.57 337.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 339 2.86 339.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 339 -1025.57 339.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 340.6 2.86 341 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 340.6 -1025.57 341 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 342.2 2.86 342.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 342.2 -907.68 342.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 343.8 2.86 344.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 343.8 -907.68 344.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.4 2.86 345.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.4 -1025.57 345.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 347 2.86 347.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 347 -1025.57 347.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 348.6 2.86 349 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 348.6 -1025.57 349 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.2 2.86 350.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.2 -1025.57 350.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 351.8 2.86 352.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 351.8 -1025.57 352.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 353.4 2.86 353.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 353.4 -828.18 353.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 353.4 -902.38 353.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 355 2.86 355.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 355 -828.18 355.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 355 -1025.57 355.4 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 356.6 2.86 357 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 356.6 -844.08 357 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 356.6 -1025.57 357 -926.12 ;
    END
    PORT
      LAYER met3 ;
        RECT 358.2 2.86 358.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 358.2 -1025.57 358.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 359.8 2.86 360.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 359.8 -1025.57 360.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 361.4 2.86 361.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 361.4 -1025.57 361.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 363 2.86 363.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 363 -1025.57 363.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 364.6 2.86 365 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 364.6 -1025.57 365 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 366.2 2.86 366.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 366.2 -1025.57 366.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 367.8 2.86 368.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 367.8 -1025.57 368.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 369.4 2.86 369.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 369.4 -1025.57 369.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 371 2.86 371.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 371 -1025.57 371.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 372.6 2.86 373 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 372.6 -828.18 373 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 372.6 -902.38 373 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 374.2 2.86 374.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 374.2 -839.84 374.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 374.2 -1025.57 374.6 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 375.8 2.86 376.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 375.8 -1025.57 376.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 377.4 2.86 377.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 377.4 -1025.57 377.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 379 2.86 379.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 379 -1025.57 379.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 380.6 2.86 381 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 380.6 -1025.57 381 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 382.2 2.86 382.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 382.2 -907.68 382.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 383.8 2.86 384.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 383.8 -907.68 384.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 383.8 -1025.57 384.2 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 385.4 2.86 385.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 385.4 -1025.57 385.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 387 2.86 387.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 387 -1025.57 387.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 388.6 2.86 389 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 388.6 -1025.57 389 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 390.2 2.86 390.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 390.2 -1025.57 390.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 391.8 2.86 392.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 391.8 -1025.57 392.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 393.4 2.86 393.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 393.4 -828.18 393.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 393.4 -902.38 393.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 395 2.86 395.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 395 -828.18 395.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 395 -1025.57 395.4 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 396.6 2.86 397 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 396.6 -1025.57 397 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 398.2 2.86 398.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 398.2 -1025.57 398.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 399.8 2.86 400.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 399.8 -1025.57 400.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 401.4 2.86 401.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 401.4 -1025.57 401.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 403 2.86 403.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 403 -1025.57 403.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 404.6 2.86 405 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 404.6 -1025.57 405 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 406.2 2.86 406.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 406.2 -1025.57 406.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 407.8 2.86 408.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 407.8 -1025.57 408.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 409.4 2.86 409.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 409.4 -1025.57 409.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 411 2.86 411.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 411 -1025.57 411.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 412.6 2.86 413 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 412.6 -828.18 413 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 412.6 -902.38 413 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 414.2 2.86 414.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 414.2 -839.84 414.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 414.2 -1025.57 414.6 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 415.8 2.86 416.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 415.8 -1025.57 416.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 417.4 2.86 417.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 417.4 -1025.57 417.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 419 2.86 419.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 419 -1025.57 419.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 420.6 2.86 421 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 420.6 -1025.57 421 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 422.2 2.86 422.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 422.2 -907.68 422.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 423.8 2.86 424.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 423.8 -907.68 424.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 423.8 -1025.57 424.2 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 425.4 2.86 425.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 425.4 -1025.57 425.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 427 2.86 427.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 427 -1025.57 427.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 428.6 2.86 429 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 428.6 -1025.57 429 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 430.2 2.86 430.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 430.2 -1025.57 430.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 431.8 2.86 432.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 431.8 -1025.57 432.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 433.4 2.86 433.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 433.4 -828.18 433.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 433.4 -902.38 433.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 435 2.86 435.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 435 -828.18 435.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 435 -1025.57 435.4 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 436.6 2.86 437 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 436.6 -1025.57 437 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 438.2 2.86 438.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 438.2 -1025.57 438.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 439.8 2.86 440.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 439.8 -1025.57 440.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 441.4 2.86 441.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 441.4 -1025.57 441.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 443 2.86 443.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 443 -1025.57 443.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 444.6 2.86 445 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 444.6 -1025.57 445 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 446.2 2.86 446.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 446.2 -1025.57 446.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 447.8 2.86 448.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 447.8 -1025.57 448.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 449.4 2.86 449.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 449.4 -1025.57 449.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 451 2.86 451.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 451 -1025.57 451.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 452.6 2.86 453 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 452.6 -828.18 453 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 452.6 -902.38 453 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 454.2 2.86 454.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 454.2 -839.84 454.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 454.2 -1025.57 454.6 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 455.8 2.86 456.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 455.8 -1025.57 456.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 457.4 2.86 457.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 457.4 -1025.57 457.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 459 2.86 459.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 459 -1025.57 459.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 460.6 2.86 461 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 460.6 -1025.57 461 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 462.2 2.86 462.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 462.2 -907.68 462.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 463.8 2.86 464.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 463.8 -907.68 464.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 463.8 -1025.57 464.2 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 465.4 2.86 465.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 465.4 -1025.57 465.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 467 2.86 467.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 467 -1025.57 467.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 468.6 2.86 469 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 468.6 -1025.57 469 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 470.2 2.86 470.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 470.2 -1025.57 470.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 471.8 2.86 472.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 471.8 -1025.57 472.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 473.4 2.86 473.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 473.4 -828.18 473.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 473.4 -902.38 473.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 475 2.86 475.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 475 -828.18 475.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 475 -1025.57 475.4 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 476.6 2.86 477 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 476.6 -1025.57 477 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 478.2 2.86 478.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 478.2 -1025.57 478.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 479.8 2.86 480.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 479.8 -1025.57 480.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 481.4 2.86 481.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 481.4 -1025.57 481.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 483 2.86 483.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 483 -1025.57 483.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 484.6 2.86 485 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 484.6 -1025.57 485 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 486.2 2.86 486.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 486.2 -1025.57 486.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 487.8 2.86 488.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 487.8 -1025.57 488.2 -818 ;
        RECT 487.75 -905.075 488.2 -904.745 ;
        RECT 487.75 -919.215 488.2 -918.885 ;
    END
    PORT
      LAYER met3 ;
        RECT 489.4 2.86 489.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 489.4 -1025.57 489.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 491 2.86 491.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 491 -1025.57 491.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 492.6 2.86 493 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 492.6 -828.18 493 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 492.6 -902.38 493 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 494.2 2.86 494.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 494.2 -839.84 494.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 494.2 -1025.57 494.6 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 495.8 2.86 496.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 495.8 -1025.57 496.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 497.4 2.86 497.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 497.4 -1025.57 497.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 499 2.86 499.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 499 -1025.57 499.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 500.6 2.86 501 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 500.6 -1025.57 501 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 502.2 2.86 502.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 502.2 -907.68 502.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 503.8 2.86 504.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 503.8 -907.68 504.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 505.4 2.86 505.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 505.4 -1025.57 505.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 507 2.86 507.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 507 -1025.57 507.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 508.6 2.86 509 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 508.6 -1025.57 509 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 510.2 2.86 510.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 510.2 -1025.57 510.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 511.8 2.86 512.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 511.8 -1025.57 512.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 513.4 2.86 513.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 513.4 -828.18 513.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 513.4 -902.38 513.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 515 2.86 515.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 515 -828.18 515.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 515 -1025.57 515.4 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 516.6 2.86 517 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 516.6 -844.08 517 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 516.6 -1025.57 517 -926.12 ;
    END
    PORT
      LAYER met3 ;
        RECT 518.2 2.86 518.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 518.2 -1025.57 518.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 519.8 2.86 520.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 519.8 -1025.57 520.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 521.4 2.86 521.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 521.4 -1025.57 521.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 523 2.86 523.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 523 -1025.57 523.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 524.6 2.86 525 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 524.6 -1025.57 525 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 526.2 2.86 526.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 526.2 -1025.57 526.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 527.8 2.86 528.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 527.8 -1025.57 528.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 529.4 2.86 529.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 529.4 -1025.57 529.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 531 2.86 531.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 531 -1025.57 531.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 532.6 2.86 533 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 532.6 -828.18 533 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 532.6 -902.38 533 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 534.2 2.86 534.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 534.2 -839.84 534.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 534.2 -1025.57 534.6 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 535.8 2.86 536.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 535.8 -1025.57 536.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 537.4 2.86 537.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 537.4 -1025.57 537.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 539 2.86 539.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 539 -1025.57 539.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 540.6 2.86 541 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 540.6 -1025.57 541 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 542.2 2.86 542.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 542.2 -907.68 542.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 543.8 2.86 544.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 543.8 -907.68 544.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 543.8 -1025.57 544.2 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 545.4 2.86 545.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 545.4 -1025.57 545.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 547 2.86 547.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 547 -1025.57 547.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 548.6 2.86 549 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 548.6 -1025.57 549 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 550.2 2.86 550.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 550.2 -1025.57 550.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 551.8 2.86 552.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 551.8 -1025.57 552.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 553.4 2.86 553.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 553.4 -828.18 553.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 553.4 -902.38 553.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 555 2.86 555.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 555 -828.18 555.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 555 -1025.57 555.4 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 556.6 2.86 557 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 556.6 -1025.57 557 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 558.2 2.86 558.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 558.2 -1025.57 558.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 559.8 2.86 560.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 559.8 -1025.57 560.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 561.4 2.86 561.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 561.4 -1025.57 561.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 563 2.86 563.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 563 -1025.57 563.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 564.6 2.86 565 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 564.6 -1025.57 565 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 566.2 2.86 566.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 566.2 -1025.57 566.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 567.8 2.86 568.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 567.8 -1025.57 568.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 569.4 2.86 569.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 569.4 -1025.57 569.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 571 2.86 571.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 571 -1025.57 571.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 572.6 2.86 573 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 572.6 -828.18 573 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 572.6 -902.38 573 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 574.2 2.86 574.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 574.2 -839.84 574.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 574.2 -1025.57 574.6 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 575.8 2.86 576.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 575.8 -1025.57 576.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 577.4 2.86 577.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 577.4 -1025.57 577.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 579 2.86 579.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 579 -1025.57 579.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 580.6 2.86 581 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 580.6 -1025.57 581 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 582.2 2.86 582.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 582.2 -907.68 582.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 583.8 2.86 584.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 583.8 -907.68 584.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 583.8 -1025.57 584.2 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 585.4 2.86 585.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 585.4 -1025.57 585.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 587 2.86 587.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 587 -1025.57 587.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 588.6 2.86 589 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 588.6 -1025.57 589 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 590.2 2.86 590.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 590.2 -1025.57 590.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 591.8 2.86 592.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 591.8 -1025.57 592.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 593.4 2.86 593.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 593.4 -828.18 593.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 593.4 -902.38 593.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 595 2.86 595.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 595 -828.18 595.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 595 -1025.57 595.4 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 596.6 2.86 597 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 596.6 -1025.57 597 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 598.2 2.86 598.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 598.2 -1025.57 598.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 599.8 2.86 600.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 599.8 -1025.57 600.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 601.4 2.86 601.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 601.4 -1025.57 601.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 603 2.86 603.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 603 -1025.57 603.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 604.6 2.86 605 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 604.6 -1025.57 605 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 606.2 2.86 606.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 606.2 -1025.57 606.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 607.8 2.86 608.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 607.8 -1025.57 608.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 609.4 2.86 609.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 609.4 -1025.57 609.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 611 2.86 611.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 611 -1025.57 611.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 612.6 2.86 613 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 612.6 -828.18 613 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 612.6 -902.38 613 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 614.2 2.86 614.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 614.2 -839.84 614.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 614.2 -1025.57 614.6 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 615.8 2.86 616.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 615.8 -1025.57 616.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 617.4 2.86 617.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 617.4 -1025.57 617.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 619 2.86 619.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 619 -1025.57 619.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 620.6 2.86 621 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 620.6 -1025.57 621 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 622.2 2.86 622.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 622.2 -907.68 622.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 623.8 2.86 624.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 623.8 -907.68 624.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 623.8 -1025.57 624.2 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 625.4 2.86 625.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 625.4 -1025.57 625.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 627 2.86 627.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 627 -1025.57 627.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 628.6 2.86 629 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 628.6 -1025.57 629 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 630.2 2.86 630.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 630.2 -1025.57 630.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 631.8 2.86 632.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 631.8 -1025.57 632.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 633.4 2.86 633.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 633.4 -828.18 633.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 633.4 -902.38 633.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 635 2.86 635.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 635 -828.18 635.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 635 -1025.57 635.4 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 636.6 2.86 637 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 636.6 -1025.57 637 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 638.2 2.86 638.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 638.2 -1025.57 638.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 639.8 2.86 640.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 639.8 -1025.57 640.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 641.4 2.86 641.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 641.4 -1025.57 641.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 643 2.86 643.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 643 -1025.57 643.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 644.6 2.86 645 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 644.6 -1025.57 645 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 646.2 2.86 646.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 646.2 -1025.57 646.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 647.8 2.86 648.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 647.8 -1025.57 648.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 649.4 2.86 649.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 649.4 -1025.57 649.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 651 -1025.57 651.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 652.6 -1025.57 653 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 654.2 -1025.57 654.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 655.8 -1025.57 656.2 11.315 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT -87.4 -1024.03 -87 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -85.8 -1024.03 -85.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -84.2 -1024.03 -83.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -82.6 -1024.03 -82.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -81 -993.54 -80.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -79.4 -1012.62 -79 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -79.4 -1024.03 -79 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -77.8 -1024.03 -77.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -76.2 -1007.32 -75.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -76.2 -1024.03 -75.8 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -74.6 -1012.62 -74.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -73 -1024.03 -72.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -71.4 -1006.26 -71 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -71.4 -1024.03 -71 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -69.8 -1007.32 -69.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -69.8 -1024.03 -69.4 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -68.2 -1012.62 -67.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -68.2 -1024.03 -67.8 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -66.6 -1024.03 -66.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -65 -1005.2 -64.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -65 -1024.03 -64.6 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -63.4 -1012.62 -63 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -61.8 -1012.62 -61.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -61.8 -1024.03 -61.4 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -60.2 -1024.03 -59.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -58.6 -1004.14 -58.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -58.6 -1024.03 -58.2 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -57 -1012.62 -56.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -55.4 -1024.03 -55 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.8 -1003.08 -53.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.8 -1024.03 -53.4 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -52.2 -1004.14 -51.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -50.6 -1012.62 -50.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -50.6 -1024.03 -50.2 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -49 -1024.03 -48.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.4 -1002.02 -47 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.4 -1024.03 -47 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.8 -1012.62 -45.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -44.2 -1012.62 -43.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -44.2 -1024.03 -43.8 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -42.6 -1024.03 -42.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -41 -1002.02 -40.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -41 -1024.03 -40.6 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -39.4 -1012.62 -39 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -37.8 -1024.03 -37.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.2 -1000.96 -35.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.2 -1024.03 -35.8 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -34.6 -1000.96 -34.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -33 -1012.62 -32.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -33 -1024.03 -32.6 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -31.4 -1024.03 -31 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.8 -999.9 -29.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.8 -1024.03 -29.4 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -28.2 -1012.62 -27.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.6 -1012.62 -26.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.6 -1024.03 -26.2 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -25 -1024.03 -24.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.4 -998.84 -23 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.4 -1024.03 -23 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.8 -1012.62 -21.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -20.2 -1024.03 -19.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.6 -997.78 -18.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.6 -1024.03 -18.2 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -17 -997.78 -16.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.4 -1012.62 -15 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.4 -1024.03 -15 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -13.8 -1024.03 -13.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -12.2 -996.72 -11.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -12.2 -1024.03 -11.8 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -10.6 -818.64 -10.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -10.6 -1012.62 -10.2 -975.94 ;
    END
    PORT
      LAYER met3 ;
        RECT -9 -1012.62 -8.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -9 -1024.03 -8.6 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -7.4 -1024.03 -7 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.8 -992.48 -5.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.8 -1024.03 -5.4 -1015.16 ;
        RECT -5.825 -1017.025 -5.4 -1016.695 ;
    END
    PORT
      LAYER met3 ;
        RECT -4.2 -1024.03 -3.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -2.6 -1024.03 -2.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -1 2.86 -0.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -1 -1024.03 -0.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.6 2.86 1 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.6 -1024.03 1 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.2 2.86 2.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.2 -1024.03 2.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.8 2.86 4.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.8 -1024.03 4.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.4 2.86 5.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.4 -1024.03 5.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 7 2.86 7.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 7 -1024.03 7.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.6 2.86 9 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.6 -1024.03 9 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.2 2.86 10.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.2 -1024.03 10.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.8 2.86 12.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.8 -1024.03 12.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.4 2.86 13.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.4 -828.18 13.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.4 -902.38 13.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 15 2.86 15.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 15 -828.18 15.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 15 -1024.03 15.4 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.6 2.86 17 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.6 -1024.03 17 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.2 2.86 18.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.2 -1024.03 18.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.8 2.86 20.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.8 -1024.03 20.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.4 2.86 21.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.4 -907.68 21.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 23 2.86 23.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 23 -907.68 23.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.6 2.86 25 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.6 -923.58 25 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.2 2.86 26.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.2 -1024.03 26.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.8 2.86 28.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.8 -1024.03 28.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.4 2.86 29.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.4 -1024.03 29.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 31 2.86 31.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 31 -1024.03 31.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.6 2.86 33 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.6 -828.18 33 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.6 -902.38 33 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.2 2.86 34.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.2 -839.84 34.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.2 -1024.03 34.6 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.8 2.86 36.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.8 -844.08 36.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.8 -1024.03 36.2 -926.12 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.4 2.86 37.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.4 -1024.03 37.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 39 2.86 39.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 39 -1024.03 39.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.6 2.86 41 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.6 -1024.03 41 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.2 2.86 42.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.2 -1024.03 42.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.8 2.86 44.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.8 -1024.03 44.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.4 2.86 45.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.4 -1024.03 45.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 47 2.86 47.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 47 -1024.03 47.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.6 2.86 49 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.6 -1024.03 49 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.2 2.86 50.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.2 -1024.03 50.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.8 2.86 52.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.8 -1024.03 52.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.4 2.86 53.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.4 -828.18 53.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.4 -902.38 53.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 55 2.86 55.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 55 -828.18 55.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 55 -1024.03 55.4 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.6 2.86 57 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.6 -1024.03 57 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.2 2.86 58.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.2 -1024.03 58.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.8 2.86 60.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.8 -1024.03 60.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.4 2.86 61.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.4 -907.68 61.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 63 2.86 63.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 63 -907.68 63.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.6 2.86 65 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.6 -1024.03 65 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.2 2.86 66.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.2 -1024.03 66.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.8 2.86 68.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.8 -1024.03 68.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.4 2.86 69.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.4 -1024.03 69.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 71 2.86 71.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 71 -1024.03 71.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.6 2.86 73 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.6 -828.18 73 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.6 -902.38 73 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.2 2.86 74.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.2 -839.84 74.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.2 -1024.03 74.6 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.8 2.86 76.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.8 -1024.03 76.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.4 2.86 77.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.4 -1024.03 77.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 79 2.86 79.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 79 -1024.03 79.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.6 2.86 81 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.6 -1024.03 81 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.2 2.86 82.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.2 -1024.03 82.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.8 2.86 84.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.8 -1024.03 84.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.4 2.86 85.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.4 -1024.03 85.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 87 2.86 87.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 87 -1024.03 87.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.6 2.86 89 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.6 -1024.03 89 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.2 2.86 90.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.2 -1024.03 90.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.8 2.86 92.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.8 -1024.03 92.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.4 2.86 93.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.4 -828.18 93.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.4 -902.38 93.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 95 2.86 95.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 95 -828.18 95.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 95 -1024.03 95.4 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.6 2.86 97 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.6 -1024.03 97 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.2 2.86 98.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.2 -1024.03 98.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.8 2.86 100.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.8 -1024.03 100.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.4 2.86 101.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.4 -907.68 101.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 103 2.86 103.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 103 -907.68 103.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.6 2.86 105 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.6 -1024.03 105 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.2 2.86 106.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.2 -1024.03 106.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.8 2.86 108.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.8 -1024.03 108.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.4 2.86 109.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.4 -1024.03 109.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 111 2.86 111.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 111 -1024.03 111.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.6 2.86 113 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.6 -828.18 113 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.6 -902.38 113 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.2 2.86 114.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.2 -839.84 114.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.2 -1024.03 114.6 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.8 2.86 116.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.8 -1024.03 116.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.4 2.86 117.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.4 -1024.03 117.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 119 2.86 119.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 119 -1024.03 119.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.6 2.86 121 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.6 -1024.03 121 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.2 2.86 122.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.2 -1024.03 122.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.8 2.86 124.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.8 -1024.03 124.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.4 2.86 125.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.4 -1024.03 125.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 127 2.86 127.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 127 -1024.03 127.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.6 2.86 129 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.6 -1024.03 129 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.2 2.86 130.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.2 -1024.03 130.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.8 2.86 132.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.8 -1024.03 132.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.4 2.86 133.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.4 -828.18 133.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.4 -902.38 133.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 135 2.86 135.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 135 -828.18 135.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 135 -1024.03 135.4 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.6 2.86 137 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.6 -1024.03 137 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.2 2.86 138.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.2 -1024.03 138.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.8 2.86 140.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.8 -1024.03 140.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.4 2.86 141.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.4 -907.68 141.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 143 2.86 143.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 143 -907.68 143.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.6 2.86 145 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.6 -1024.03 145 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.2 2.86 146.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.2 -1024.03 146.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.8 2.86 148.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.8 -1024.03 148.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.4 2.86 149.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.4 -1024.03 149.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 151 2.86 151.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 151 -1024.03 151.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.6 2.86 153 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.6 -828.18 153 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.6 -902.38 153 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.2 2.86 154.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.2 -839.84 154.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.2 -1024.03 154.6 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.8 2.86 156.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.8 -1024.03 156.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 157.4 2.86 157.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 157.4 -1024.03 157.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 159 2.86 159.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 159 -1024.03 159.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.6 2.86 161 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.6 -1024.03 161 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 162.2 2.86 162.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 162.2 -1024.03 162.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.8 2.86 164.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.8 -1024.03 164.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.4 2.86 165.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.4 -1024.03 165.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 167 2.86 167.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 167 -1024.03 167.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.6 2.86 169 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.6 -1024.03 169 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.2 2.86 170.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.2 -1024.03 170.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.8 2.86 172.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.8 -1024.03 172.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.4 2.86 173.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.4 -828.18 173.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.4 -902.38 173.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 175 2.86 175.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 175 -828.18 175.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 175 -1024.03 175.4 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 176.6 2.86 177 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 176.6 -1024.03 177 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.2 2.86 178.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.2 -1024.03 178.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.8 2.86 180.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.8 -1024.03 180.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 181.4 2.86 181.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 181.4 -907.68 181.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 183 2.86 183.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 183 -907.68 183.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.6 2.86 185 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.6 -923.58 185 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.2 2.86 186.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.2 -1024.03 186.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 187.8 2.86 188.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 187.8 -1024.03 188.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.4 2.86 189.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.4 -1024.03 189.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 191 2.86 191.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 191 -1024.03 191.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.6 2.86 193 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.6 -828.18 193 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.6 -902.38 193 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.2 2.86 194.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.2 -839.84 194.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.2 -1024.03 194.6 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.8 2.86 196.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.8 -844.08 196.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.8 -1024.03 196.2 -926.12 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.4 2.86 197.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.4 -1024.03 197.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 199 2.86 199.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 199 -1024.03 199.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.6 2.86 201 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.6 -1024.03 201 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 202.2 2.86 202.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 202.2 -1024.03 202.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.8 2.86 204.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.8 -1024.03 204.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.4 2.86 205.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.4 -1024.03 205.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 207 2.86 207.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 207 -1024.03 207.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 208.6 2.86 209 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 208.6 -1024.03 209 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 210.2 2.86 210.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 210.2 -1024.03 210.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.8 2.86 212.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.8 -1024.03 212.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 213.4 2.86 213.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 213.4 -828.18 213.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 213.4 -902.38 213.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 215 2.86 215.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 215 -828.18 215.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 215 -1024.03 215.4 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.6 2.86 217 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.6 -1024.03 217 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.2 2.86 218.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.2 -1024.03 218.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 219.8 2.86 220.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 219.8 -1024.03 220.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 221.4 2.86 221.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 221.4 -907.68 221.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 223 2.86 223.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 223 -907.68 223.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.6 2.86 225 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.6 -1024.03 225 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.2 2.86 226.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.2 -1024.03 226.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 227.8 2.86 228.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 227.8 -1024.03 228.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 229.4 2.86 229.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 229.4 -1024.03 229.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 231 2.86 231.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 231 -1024.03 231.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 232.6 2.86 233 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 232.6 -828.18 233 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 232.6 -902.38 233 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.2 2.86 234.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.2 -839.84 234.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.2 -1024.03 234.6 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.8 2.86 236.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.8 -1024.03 236.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.4 2.86 237.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.4 -1024.03 237.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 239 2.86 239.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 239 -1024.03 239.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 240.6 2.86 241 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 240.6 -1024.03 241 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 242.2 2.86 242.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 242.2 -1024.03 242.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.8 2.86 244.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.8 -1024.03 244.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.4 2.86 245.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.4 -1024.03 245.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 247 2.86 247.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 247 -1024.03 247.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.6 2.86 249 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.6 -1024.03 249 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.2 2.86 250.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.2 -1024.03 250.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 251.8 2.86 252.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 251.8 -1024.03 252.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 253.4 2.86 253.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 253.4 -828.18 253.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 253.4 -902.38 253.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 255 2.86 255.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 255 -828.18 255.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 255 -1024.03 255.4 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.6 2.86 257 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.6 -1024.03 257 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.2 2.86 258.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.2 -1024.03 258.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 259.8 2.86 260.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 259.8 -1024.03 260.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 261.4 2.86 261.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 261.4 -907.68 261.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 263 2.86 263.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 263 -907.68 263.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.6 2.86 265 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.6 -1024.03 265 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 266.2 2.86 266.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 266.2 -1024.03 266.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.8 2.86 268.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.8 -1024.03 268.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.4 2.86 269.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.4 -1024.03 269.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 271 2.86 271.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 271 -1024.03 271.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 272.6 2.86 273 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 272.6 -828.18 273 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 272.6 -902.38 273 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 274.2 2.86 274.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 274.2 -839.84 274.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 274.2 -1024.03 274.6 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.8 2.86 276.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.8 -1024.03 276.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.4 2.86 277.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.4 -1024.03 277.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 279 2.86 279.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 279 -1024.03 279.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 280.6 2.86 281 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 280.6 -1024.03 281 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.2 2.86 282.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.2 -1024.03 282.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 283.8 2.86 284.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 283.8 -1024.03 284.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 285.4 2.86 285.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 285.4 -1024.03 285.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 287 2.86 287.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 287 -1024.03 287.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.6 2.86 289 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.6 -1024.03 289 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.2 2.86 290.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.2 -1024.03 290.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 291.8 2.86 292.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 291.8 -1024.03 292.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 293.4 2.86 293.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 293.4 -828.18 293.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 293.4 -902.38 293.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 295 2.86 295.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 295 -828.18 295.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 295 -1024.03 295.4 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.6 2.86 297 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.6 -1024.03 297 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 298.2 2.86 298.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 298.2 -1024.03 298.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.8 2.86 300.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.8 -1024.03 300.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.4 2.86 301.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.4 -907.68 301.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 303 2.86 303.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 303 -907.68 303.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 304.6 2.86 305 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 304.6 -1024.03 305 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 306.2 2.86 306.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 306.2 -1024.03 306.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.8 2.86 308.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.8 -1024.03 308.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.4 2.86 309.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.4 -1024.03 309.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 311 2.86 311.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 311 -1024.03 311.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 312.6 2.86 313 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 312.6 -828.18 313 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 312.6 -902.38 313 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 314.2 2.86 314.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 314.2 -839.84 314.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 314.2 -1024.03 314.6 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 315.8 2.86 316.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 315.8 -1024.03 316.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 317.4 2.86 317.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 317.4 -1024.03 317.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 319 2.86 319.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 319 -1024.03 319.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.6 2.86 321 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.6 -1024.03 321 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.2 2.86 322.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.2 -1024.03 322.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 323.8 2.86 324.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 323.8 -1024.03 324.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 325.4 2.86 325.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 325.4 -1024.03 325.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 327 2.86 327.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 327 -1024.03 327.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.6 2.86 329 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.6 -1024.03 329 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.2 2.86 330.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.2 -1024.03 330.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 331.8 2.86 332.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 331.8 -1024.03 332.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.4 2.86 333.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.4 -828.18 333.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.4 -902.38 333.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 335 2.86 335.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 335 -828.18 335.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 335 -1024.03 335.4 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 336.6 2.86 337 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 336.6 -1024.03 337 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 338.2 2.86 338.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 338.2 -1024.03 338.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.8 2.86 340.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.8 -1024.03 340.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 341.4 2.86 341.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 341.4 -907.68 341.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 343 2.86 343.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 343 -907.68 343.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 344.6 2.86 345 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 344.6 -923.58 345 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 346.2 2.86 346.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 346.2 -1024.03 346.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.8 2.86 348.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.8 -1024.03 348.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 349.4 2.86 349.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 349.4 -1024.03 349.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 351 2.86 351.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 351 -1024.03 351.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.6 2.86 353 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.6 -828.18 353 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.6 -902.38 353 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.2 2.86 354.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.2 -839.84 354.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.2 -1024.03 354.6 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 355.8 2.86 356.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 355.8 -844.08 356.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 355.8 -1024.03 356.2 -926.12 ;
    END
    PORT
      LAYER met3 ;
        RECT 357.4 2.86 357.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 357.4 -1024.03 357.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 359 2.86 359.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 359 -1024.03 359.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 360.6 2.86 361 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 360.6 -1024.03 361 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 362.2 2.86 362.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 362.2 -1024.03 362.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 363.8 2.86 364.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 363.8 -1024.03 364.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 365.4 2.86 365.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 365.4 -1024.03 365.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 367 2.86 367.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 367 -1024.03 367.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 368.6 2.86 369 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 368.6 -1024.03 369 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 370.2 2.86 370.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 370.2 -1024.03 370.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 371.8 2.86 372.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 371.8 -1024.03 372.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 373.4 2.86 373.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 373.4 -828.18 373.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 373.4 -902.38 373.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 375 2.86 375.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 375 -828.18 375.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 375 -1024.03 375.4 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 376.6 2.86 377 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 376.6 -1024.03 377 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 378.2 2.86 378.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 378.2 -1024.03 378.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 379.8 2.86 380.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 379.8 -1024.03 380.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 381.4 2.86 381.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 381.4 -907.68 381.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 383 2.86 383.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 383 -907.68 383.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 384.6 2.86 385 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 384.6 -1024.03 385 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 386.2 2.86 386.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 386.2 -1024.03 386.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 387.8 2.86 388.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 387.8 -1024.03 388.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 389.4 2.86 389.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 389.4 -1024.03 389.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 391 2.86 391.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 391 -1024.03 391.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 392.6 2.86 393 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 392.6 -828.18 393 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 392.6 -902.38 393 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 394.2 2.86 394.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 394.2 -839.84 394.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 394.2 -1024.03 394.6 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 395.8 2.86 396.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 395.8 -1024.03 396.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 397.4 2.86 397.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 397.4 -1024.03 397.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 399 2.86 399.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 399 -1024.03 399.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 400.6 2.86 401 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 400.6 -1024.03 401 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 402.2 2.86 402.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 402.2 -1024.03 402.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 403.8 2.86 404.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 403.8 -1024.03 404.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 405.4 2.86 405.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 405.4 -1024.03 405.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 407 2.86 407.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 407 -1024.03 407.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 408.6 2.86 409 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 408.6 -1024.03 409 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 410.2 2.86 410.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 410.2 -1024.03 410.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 411.8 2.86 412.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 411.8 -1024.03 412.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 413.4 2.86 413.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 413.4 -828.18 413.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 413.4 -902.38 413.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 415 2.86 415.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 415 -828.18 415.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 415 -1024.03 415.4 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 416.6 2.86 417 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 416.6 -1024.03 417 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 418.2 2.86 418.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 418.2 -1024.03 418.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 419.8 2.86 420.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 419.8 -1024.03 420.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 421.4 2.86 421.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 421.4 -907.68 421.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 423 2.86 423.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 423 -907.68 423.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 424.6 2.86 425 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 424.6 -1024.03 425 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 426.2 2.86 426.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 426.2 -1024.03 426.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 427.8 2.86 428.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 427.8 -1024.03 428.2 -818 ;
        RECT 427.75 -928.085 428.2 -927.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 429.4 2.86 429.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 429.4 -1024.03 429.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 431 2.86 431.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 431 -1024.03 431.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 432.6 2.86 433 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 432.6 -828.18 433 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 432.6 -902.38 433 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 434.2 2.86 434.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 434.2 -839.84 434.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 434.2 -1024.03 434.6 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 435.8 2.86 436.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 435.8 -1024.03 436.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 437.4 2.86 437.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 437.4 -1024.03 437.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 439 2.86 439.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 439 -1024.03 439.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 440.6 2.86 441 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 440.6 -1024.03 441 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 442.2 2.86 442.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 442.2 -1024.03 442.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 443.8 2.86 444.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 443.8 -1024.03 444.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 445.4 2.86 445.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 445.4 -1024.03 445.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 447 2.86 447.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 447 -1024.03 447.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 448.6 2.86 449 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 448.6 -1024.03 449 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 450.2 2.86 450.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 450.2 -1024.03 450.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 451.8 2.86 452.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 451.8 -1024.03 452.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 453.4 2.86 453.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 453.4 -828.18 453.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 453.4 -902.38 453.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 455 2.86 455.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 455 -828.18 455.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 455 -1024.03 455.4 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 456.6 2.86 457 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 456.6 -1024.03 457 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 458.2 2.86 458.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 458.2 -1024.03 458.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 459.8 2.86 460.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 459.8 -1024.03 460.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 461.4 2.86 461.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 461.4 -907.68 461.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 463 2.86 463.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 463 -907.68 463.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 464.6 2.86 465 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 464.6 -1024.03 465 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 466.2 2.86 466.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 466.2 -1024.03 466.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 467.8 2.86 468.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 467.8 -1024.03 468.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 469.4 2.86 469.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 469.4 -1024.03 469.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 471 2.86 471.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 471 -1024.03 471.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 472.6 2.86 473 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 472.6 -828.18 473 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 472.6 -902.38 473 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 474.2 2.86 474.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 474.2 -839.84 474.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 474.2 -1024.03 474.6 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 475.8 2.86 476.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 475.8 -1024.03 476.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 477.4 2.86 477.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 477.4 -1024.03 477.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 479 2.86 479.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 479 -1024.03 479.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 480.6 2.86 481 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 480.6 -1024.03 481 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 482.2 2.86 482.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 482.2 -1024.03 482.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 483.8 2.86 484.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 483.8 -1024.03 484.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 485.4 2.86 485.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 485.4 -1024.03 485.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 487 2.86 487.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 487 -1024.03 487.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 488.6 2.86 489 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 488.6 -1024.03 489 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 490.2 2.86 490.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 490.2 -1024.03 490.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 491.8 2.86 492.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 491.8 -1024.03 492.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 493.4 2.86 493.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 493.4 -828.18 493.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 493.4 -902.38 493.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 495 2.86 495.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 495 -828.18 495.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 495 -1024.03 495.4 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 496.6 2.86 497 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 496.6 -1024.03 497 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 498.2 2.86 498.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 498.2 -1024.03 498.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 499.8 2.86 500.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 499.8 -1024.03 500.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 501.4 2.86 501.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 501.4 -907.68 501.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 503 2.86 503.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 503 -907.68 503.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 504.6 2.86 505 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 504.6 -923.58 505 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 506.2 2.86 506.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 506.2 -1024.03 506.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 507.8 2.86 508.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 507.8 -1024.03 508.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 509.4 2.86 509.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 509.4 -1024.03 509.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 511 2.86 511.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 511 -1024.03 511.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 512.6 2.86 513 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 512.6 -828.18 513 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 512.6 -902.38 513 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 514.2 2.86 514.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 514.2 -839.84 514.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 514.2 -1024.03 514.6 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 515.8 2.86 516.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 515.8 -844.08 516.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 515.8 -1024.03 516.2 -926.12 ;
    END
    PORT
      LAYER met3 ;
        RECT 517.4 2.86 517.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 517.4 -1024.03 517.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 519 2.86 519.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 519 -1024.03 519.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 520.6 2.86 521 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 520.6 -1024.03 521 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 522.2 2.86 522.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 522.2 -1024.03 522.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 523.8 2.86 524.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 523.8 -1024.03 524.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 525.4 2.86 525.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 525.4 -1024.03 525.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 527 2.86 527.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 527 -1024.03 527.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 528.6 2.86 529 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 528.6 -1024.03 529 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 530.2 2.86 530.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 530.2 -1024.03 530.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 531.8 2.86 532.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 531.8 -1024.03 532.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 533.4 2.86 533.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 533.4 -828.18 533.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 533.4 -902.38 533.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 535 2.86 535.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 535 -828.18 535.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 535 -1024.03 535.4 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 536.6 2.86 537 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 536.6 -1024.03 537 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 538.2 2.86 538.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 538.2 -1024.03 538.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 539.8 2.86 540.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 539.8 -1024.03 540.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 541.4 2.86 541.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 541.4 -907.68 541.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 543 2.86 543.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 543 -907.68 543.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 544.6 2.86 545 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 544.6 -1024.03 545 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 546.2 2.86 546.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 546.2 -1024.03 546.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 547.8 2.86 548.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 547.8 -1024.03 548.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 549.4 2.86 549.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 549.4 -1024.03 549.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 551 2.86 551.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 551 -1024.03 551.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 552.6 2.86 553 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 552.6 -828.18 553 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 552.6 -902.38 553 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 554.2 2.86 554.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 554.2 -839.84 554.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 554.2 -1024.03 554.6 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 555.8 2.86 556.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 555.8 -1024.03 556.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 557.4 2.86 557.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 557.4 -1024.03 557.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 559 2.86 559.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 559 -1024.03 559.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 560.6 2.86 561 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 560.6 -1024.03 561 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 562.2 2.86 562.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 562.2 -1024.03 562.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 563.8 2.86 564.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 563.8 -1024.03 564.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 565.4 2.86 565.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 565.4 -1024.03 565.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 567 2.86 567.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 567 -1024.03 567.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 568.6 2.86 569 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 568.6 -1024.03 569 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 570.2 2.86 570.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 570.2 -1024.03 570.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 571.8 2.86 572.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 571.8 -1024.03 572.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 573.4 2.86 573.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 573.4 -828.18 573.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 573.4 -902.38 573.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 575 2.86 575.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 575 -828.18 575.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 575 -1024.03 575.4 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 576.6 2.86 577 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 576.6 -1024.03 577 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 578.2 2.86 578.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 578.2 -1024.03 578.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 579.8 2.86 580.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 579.8 -1024.03 580.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 581.4 2.86 581.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 581.4 -907.68 581.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 583 2.86 583.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 583 -907.68 583.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 584.6 2.86 585 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 584.6 -1024.03 585 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 586.2 2.86 586.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 586.2 -1024.03 586.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 587.8 2.86 588.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 587.8 -1024.03 588.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 589.4 2.86 589.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 589.4 -1024.03 589.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 591 2.86 591.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 591 -1024.03 591.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 592.6 2.86 593 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 592.6 -828.18 593 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 592.6 -902.38 593 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 594.2 2.86 594.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 594.2 -839.84 594.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 594.2 -1024.03 594.6 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 595.8 2.86 596.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 595.8 -1024.03 596.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 597.4 2.86 597.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 597.4 -1024.03 597.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 599 2.86 599.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 599 -1024.03 599.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 600.6 2.86 601 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 600.6 -1024.03 601 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 602.2 2.86 602.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 602.2 -1024.03 602.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 603.8 2.86 604.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 603.8 -1024.03 604.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 605.4 2.86 605.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 605.4 -1024.03 605.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 607 2.86 607.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 607 -1024.03 607.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 608.6 2.86 609 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 608.6 -1024.03 609 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 610.2 2.86 610.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 610.2 -1024.03 610.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 611.8 2.86 612.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 611.8 -1024.03 612.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 613.4 2.86 613.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 613.4 -828.18 613.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 613.4 -902.38 613.8 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 615 2.86 615.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 615 -828.18 615.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 615 -1024.03 615.4 -909.16 ;
    END
    PORT
      LAYER met3 ;
        RECT 616.6 2.86 617 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 616.6 -1024.03 617 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 618.2 2.86 618.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 618.2 -1024.03 618.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 619.8 2.86 620.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 619.8 -1024.03 620.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 621.4 2.86 621.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 621.4 -907.68 621.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 623 2.86 623.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 623 -907.68 623.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 624.6 2.86 625 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 624.6 -1024.03 625 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 626.2 2.86 626.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 626.2 -1024.03 626.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 627.8 2.86 628.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 627.8 -1024.03 628.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 629.4 2.86 629.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 629.4 -1024.03 629.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 631 2.86 631.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 631 -1024.03 631.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 632.6 2.86 633 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 632.6 -828.18 633 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 632.6 -902.38 633 -893.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 634.2 2.86 634.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 634.2 -839.84 634.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 634.2 -1024.03 634.6 -916.58 ;
    END
    PORT
      LAYER met3 ;
        RECT 635.8 2.86 636.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 635.8 -1024.03 636.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 637.4 2.86 637.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 637.4 -1024.03 637.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 639 2.86 639.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 639 -1024.03 639.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 640.6 2.86 641 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 640.6 -1024.03 641 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 642.2 2.86 642.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 642.2 -1024.03 642.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 643.8 2.86 644.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 643.8 -1024.03 644.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 645.4 2.86 645.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 645.4 -1024.03 645.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 647 2.86 647.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 647 -1024.03 647.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 648.6 2.86 649 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 648.6 -1024.03 649 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 650.2 2.86 650.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 650.2 -1024.03 650.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 651.8 -1024.03 652.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 653.4 -1024.03 653.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 655 -1024.03 655.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 656.6 -1024.03 657 9.775 ;
    END
  END vss
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -16.46 -1025.97 -16.16 -1025.67 ;
    END
  END addr[0]
  PIN addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -74.86 -1025.97 -74.56 -1025.67 ;
    END
  END addr[10]
  PIN addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -80.7 -1025.97 -80.4 -1025.67 ;
    END
  END addr[11]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -22.3 -1025.97 -22 -1025.67 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -28.14 -1025.97 -27.84 -1025.67 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -33.98 -1025.97 -33.68 -1025.67 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -39.82 -1025.97 -39.52 -1025.67 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -45.66 -1025.97 -45.36 -1025.67 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -51.5 -1025.97 -51.2 -1025.67 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -57.34 -1025.97 -57.04 -1025.67 ;
    END
  END addr[7]
  PIN addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -63.18 -1025.97 -62.88 -1025.67 ;
    END
  END addr[8]
  PIN addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -69.02 -1025.97 -68.72 -1025.67 ;
    END
  END addr[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -81.72 -1025.97 -81.3 -1025.55 ;
    END
  END clk
  PIN din[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.015 -1025.97 22.315 -1025.67 ;
    END
  END din[0]
  PIN din[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 222.015 -1025.97 222.315 -1025.67 ;
    END
  END din[10]
  PIN din[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 222.63 -1025.97 222.93 -1025.67 ;
    END
  END din[11]
  PIN din[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.015 -1025.97 262.315 -1025.67 ;
    END
  END din[12]
  PIN din[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.63 -1025.97 262.93 -1025.67 ;
    END
  END din[13]
  PIN din[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 302.015 -1025.97 302.315 -1025.67 ;
    END
  END din[14]
  PIN din[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 302.63 -1025.97 302.93 -1025.67 ;
    END
  END din[15]
  PIN din[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 342.015 -1025.97 342.315 -1025.67 ;
    END
  END din[16]
  PIN din[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 342.63 -1025.97 342.93 -1025.67 ;
    END
  END din[17]
  PIN din[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 382.015 -1025.97 382.315 -1025.67 ;
    END
  END din[18]
  PIN din[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 382.63 -1025.97 382.93 -1025.67 ;
    END
  END din[19]
  PIN din[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.63 -1025.97 22.93 -1025.67 ;
    END
  END din[1]
  PIN din[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 422.015 -1025.97 422.315 -1025.67 ;
    END
  END din[20]
  PIN din[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 422.63 -1025.97 422.93 -1025.67 ;
    END
  END din[21]
  PIN din[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 462.015 -1025.97 462.315 -1025.67 ;
    END
  END din[22]
  PIN din[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 462.63 -1025.97 462.93 -1025.67 ;
    END
  END din[23]
  PIN din[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 502.015 -1025.97 502.315 -1025.67 ;
    END
  END din[24]
  PIN din[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 502.63 -1025.97 502.93 -1025.67 ;
    END
  END din[25]
  PIN din[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 542.015 -1025.97 542.315 -1025.67 ;
    END
  END din[26]
  PIN din[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 542.63 -1025.97 542.93 -1025.67 ;
    END
  END din[27]
  PIN din[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.015 -1025.97 582.315 -1025.67 ;
    END
  END din[28]
  PIN din[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.63 -1025.97 582.93 -1025.67 ;
    END
  END din[29]
  PIN din[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 62.015 -1025.97 62.315 -1025.67 ;
    END
  END din[2]
  PIN din[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 622.015 -1025.97 622.315 -1025.67 ;
    END
  END din[30]
  PIN din[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 622.63 -1025.97 622.93 -1025.67 ;
    END
  END din[31]
  PIN din[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 62.63 -1025.97 62.93 -1025.67 ;
    END
  END din[3]
  PIN din[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 102.015 -1025.97 102.315 -1025.67 ;
    END
  END din[4]
  PIN din[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 102.63 -1025.97 102.93 -1025.67 ;
    END
  END din[5]
  PIN din[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 142.015 -1025.97 142.315 -1025.67 ;
    END
  END din[6]
  PIN din[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 142.63 -1025.97 142.93 -1025.67 ;
    END
  END din[7]
  PIN din[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 182.015 -1025.97 182.315 -1025.67 ;
    END
  END din[8]
  PIN din[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 182.63 -1025.97 182.93 -1025.67 ;
    END
  END din[9]
  PIN dout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 13.285 -1025.97 13.585 -1025.67 ;
    END
  END dout[0]
  PIN dout[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.285 -1025.97 213.585 -1025.67 ;
    END
  END dout[10]
  PIN dout[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 233.285 -1025.97 233.585 -1025.67 ;
    END
  END dout[11]
  PIN dout[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 253.285 -1025.97 253.585 -1025.67 ;
    END
  END dout[12]
  PIN dout[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.285 -1025.97 273.585 -1025.67 ;
    END
  END dout[13]
  PIN dout[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 293.285 -1025.97 293.585 -1025.67 ;
    END
  END dout[14]
  PIN dout[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.285 -1025.97 313.585 -1025.67 ;
    END
  END dout[15]
  PIN dout[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 333.285 -1025.97 333.585 -1025.67 ;
    END
  END dout[16]
  PIN dout[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 353.285 -1025.97 353.585 -1025.67 ;
    END
  END dout[17]
  PIN dout[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 373.285 -1025.97 373.585 -1025.67 ;
    END
  END dout[18]
  PIN dout[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.285 -1025.97 393.585 -1025.67 ;
    END
  END dout[19]
  PIN dout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 33.285 -1025.97 33.585 -1025.67 ;
    END
  END dout[1]
  PIN dout[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 413.285 -1025.97 413.585 -1025.67 ;
    END
  END dout[20]
  PIN dout[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 433.285 -1025.97 433.585 -1025.67 ;
    END
  END dout[21]
  PIN dout[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 453.285 -1025.97 453.585 -1025.67 ;
    END
  END dout[22]
  PIN dout[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 473.285 -1025.97 473.585 -1025.67 ;
    END
  END dout[23]
  PIN dout[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 493.285 -1025.97 493.585 -1025.67 ;
    END
  END dout[24]
  PIN dout[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 513.285 -1025.97 513.585 -1025.67 ;
    END
  END dout[25]
  PIN dout[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 533.285 -1025.97 533.585 -1025.67 ;
    END
  END dout[26]
  PIN dout[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 553.285 -1025.97 553.585 -1025.67 ;
    END
  END dout[27]
  PIN dout[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 573.285 -1025.97 573.585 -1025.67 ;
    END
  END dout[28]
  PIN dout[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 593.285 -1025.97 593.585 -1025.67 ;
    END
  END dout[29]
  PIN dout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 53.285 -1025.97 53.585 -1025.67 ;
    END
  END dout[2]
  PIN dout[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.285 -1025.97 613.585 -1025.67 ;
    END
  END dout[30]
  PIN dout[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 633.285 -1025.97 633.585 -1025.67 ;
    END
  END dout[31]
  PIN dout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 73.285 -1025.97 73.585 -1025.67 ;
    END
  END dout[3]
  PIN dout[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 93.285 -1025.97 93.585 -1025.67 ;
    END
  END dout[4]
  PIN dout[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 113.285 -1025.97 113.585 -1025.67 ;
    END
  END dout[5]
  PIN dout[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.285 -1025.97 133.585 -1025.67 ;
    END
  END dout[6]
  PIN dout[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 153.285 -1025.97 153.585 -1025.67 ;
    END
  END dout[7]
  PIN dout[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 173.285 -1025.97 173.585 -1025.67 ;
    END
  END dout[8]
  PIN dout[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 193.285 -1025.97 193.585 -1025.67 ;
    END
  END dout[9]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -10.62 -1025.97 -10.32 -1025.67 ;
    END
  END we
  PIN wmask[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 24.125 -1025.97 24.425 -1025.67 ;
    END
  END wmask[0]
  PIN wmask[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 184.125 -1025.97 184.425 -1025.67 ;
    END
  END wmask[1]
  PIN wmask[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 344.125 -1025.97 344.425 -1025.67 ;
    END
  END wmask[2]
  PIN wmask[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 504.125 -1025.97 504.425 -1025.67 ;
    END
  END wmask[3]
  OBS
    LAYER met1 SPACING 0.14 ;
      RECT -93.555 -1025.97 662.46 11.715 ;
    LAYER met2 SPACING 0.14 ;
      RECT -93.555 -1025.97 662.46 11.715 ;
    LAYER met3 SPACING 0.3 ;
      RECT 635.115 -876.73 635.445 -876.4 ;
      RECT 635.13 -892.16 635.43 -876.4 ;
      RECT 635.115 -892.16 635.445 -891.83 ;
      RECT 635.13 -872.945 635.43 -829.2 ;
      RECT 635.115 -831.175 635.445 -830.845 ;
      RECT 635.115 -872.535 635.445 -872.205 ;
      RECT 634.515 -916.05 634.815 -840.46 ;
      RECT 634.5 -840.835 634.83 -840.505 ;
      RECT 634.5 -860.315 634.83 -859.985 ;
      RECT 634.5 -916.05 634.83 -915.72 ;
      RECT 633.9 -855.655 634.2 -841.09 ;
      RECT 633.885 -841.465 634.215 -841.135 ;
      RECT 633.885 -855.655 634.215 -855.325 ;
      RECT 633.27 -903.135 633.6 -902.805 ;
      RECT 633.285 -1025.18 633.585 -902.805 ;
      RECT 633.27 -877.19 633.6 -876.86 ;
      RECT 633.285 -892.16 633.585 -876.86 ;
      RECT 633.27 -892.16 633.6 -891.83 ;
      RECT 633.285 -872.965 633.585 -829.2 ;
      RECT 633.27 -829.575 633.6 -829.245 ;
      RECT 633.27 -872.965 633.6 -872.635 ;
      RECT 623.245 -908.525 623.575 -908.195 ;
      RECT 623.26 -1017.91 623.56 -908.195 ;
      RECT 623.245 -915.765 623.575 -915.435 ;
      RECT 623.245 -1017.865 623.575 -1017.535 ;
      RECT 622.615 -914.965 622.945 -914.635 ;
      RECT 622.63 -1025.18 622.93 -914.635 ;
      RECT 622 -909.325 622.33 -908.995 ;
      RECT 622.015 -1025.18 622.315 -908.995 ;
      RECT 615.115 -876.73 615.445 -876.4 ;
      RECT 615.13 -892.16 615.43 -876.4 ;
      RECT 615.115 -892.16 615.445 -891.83 ;
      RECT 615.13 -872.945 615.43 -829.2 ;
      RECT 615.115 -831.175 615.445 -830.845 ;
      RECT 615.115 -872.535 615.445 -872.205 ;
      RECT 614.515 -908.04 614.815 -840.46 ;
      RECT 614.5 -840.835 614.83 -840.505 ;
      RECT 614.5 -860.315 614.83 -859.985 ;
      RECT 614.5 -908.04 614.83 -907.71 ;
      RECT 613.9 -855.655 614.2 -841.09 ;
      RECT 613.885 -841.465 614.215 -841.135 ;
      RECT 613.885 -855.655 614.215 -855.325 ;
      RECT 613.27 -903.135 613.6 -902.805 ;
      RECT 613.285 -1025.18 613.585 -902.805 ;
      RECT 613.27 -877.19 613.6 -876.86 ;
      RECT 613.285 -892.16 613.585 -876.86 ;
      RECT 613.27 -892.16 613.6 -891.83 ;
      RECT 613.285 -872.965 613.585 -829.2 ;
      RECT 613.27 -829.575 613.6 -829.245 ;
      RECT 613.27 -872.965 613.6 -872.635 ;
      RECT 595.115 -876.73 595.445 -876.4 ;
      RECT 595.13 -892.16 595.43 -876.4 ;
      RECT 595.115 -892.16 595.445 -891.83 ;
      RECT 595.13 -872.945 595.43 -829.2 ;
      RECT 595.115 -831.175 595.445 -830.845 ;
      RECT 595.115 -872.535 595.445 -872.205 ;
      RECT 594.515 -916.05 594.815 -840.46 ;
      RECT 594.5 -840.835 594.83 -840.505 ;
      RECT 594.5 -860.315 594.83 -859.985 ;
      RECT 594.5 -916.05 594.83 -915.72 ;
      RECT 593.9 -855.655 594.2 -841.09 ;
      RECT 593.885 -841.465 594.215 -841.135 ;
      RECT 593.885 -855.655 594.215 -855.325 ;
      RECT 593.27 -903.135 593.6 -902.805 ;
      RECT 593.285 -1025.18 593.585 -902.805 ;
      RECT 593.27 -877.19 593.6 -876.86 ;
      RECT 593.285 -892.16 593.585 -876.86 ;
      RECT 593.27 -892.16 593.6 -891.83 ;
      RECT 593.285 -872.965 593.585 -829.2 ;
      RECT 593.27 -829.575 593.6 -829.245 ;
      RECT 593.27 -872.965 593.6 -872.635 ;
      RECT 583.245 -908.525 583.575 -908.195 ;
      RECT 583.26 -1017.91 583.56 -908.195 ;
      RECT 583.245 -915.765 583.575 -915.435 ;
      RECT 583.245 -1017.865 583.575 -1017.535 ;
      RECT 582.615 -914.965 582.945 -914.635 ;
      RECT 582.63 -1025.18 582.93 -914.635 ;
      RECT 582 -909.325 582.33 -908.995 ;
      RECT 582.015 -1025.18 582.315 -908.995 ;
      RECT 575.115 -876.73 575.445 -876.4 ;
      RECT 575.13 -892.16 575.43 -876.4 ;
      RECT 575.115 -892.16 575.445 -891.83 ;
      RECT 575.13 -872.945 575.43 -829.2 ;
      RECT 575.115 -831.175 575.445 -830.845 ;
      RECT 575.115 -872.535 575.445 -872.205 ;
      RECT 574.515 -908.04 574.815 -840.46 ;
      RECT 574.5 -840.835 574.83 -840.505 ;
      RECT 574.5 -860.315 574.83 -859.985 ;
      RECT 574.5 -908.04 574.83 -907.71 ;
      RECT 573.9 -855.655 574.2 -841.09 ;
      RECT 573.885 -841.465 574.215 -841.135 ;
      RECT 573.885 -855.655 574.215 -855.325 ;
      RECT 573.27 -903.135 573.6 -902.805 ;
      RECT 573.285 -1025.18 573.585 -902.805 ;
      RECT 573.27 -877.19 573.6 -876.86 ;
      RECT 573.285 -892.16 573.585 -876.86 ;
      RECT 573.27 -892.16 573.6 -891.83 ;
      RECT 573.285 -872.965 573.585 -829.2 ;
      RECT 573.27 -829.575 573.6 -829.245 ;
      RECT 573.27 -872.965 573.6 -872.635 ;
      RECT 555.115 -876.73 555.445 -876.4 ;
      RECT 555.13 -892.16 555.43 -876.4 ;
      RECT 555.115 -892.16 555.445 -891.83 ;
      RECT 555.13 -872.945 555.43 -829.2 ;
      RECT 555.115 -831.175 555.445 -830.845 ;
      RECT 555.115 -872.535 555.445 -872.205 ;
      RECT 554.515 -916.05 554.815 -840.46 ;
      RECT 554.5 -840.835 554.83 -840.505 ;
      RECT 554.5 -860.315 554.83 -859.985 ;
      RECT 554.5 -916.05 554.83 -915.72 ;
      RECT 553.9 -855.655 554.2 -841.09 ;
      RECT 553.885 -841.465 554.215 -841.135 ;
      RECT 553.885 -855.655 554.215 -855.325 ;
      RECT 553.27 -903.135 553.6 -902.805 ;
      RECT 553.285 -1025.18 553.585 -902.805 ;
      RECT 553.27 -877.19 553.6 -876.86 ;
      RECT 553.285 -892.16 553.585 -876.86 ;
      RECT 553.27 -892.16 553.6 -891.83 ;
      RECT 553.285 -872.965 553.585 -829.2 ;
      RECT 553.27 -829.575 553.6 -829.245 ;
      RECT 553.27 -872.965 553.6 -872.635 ;
      RECT 543.245 -908.525 543.575 -908.195 ;
      RECT 543.26 -1017.91 543.56 -908.195 ;
      RECT 543.245 -915.765 543.575 -915.435 ;
      RECT 543.245 -1017.865 543.575 -1017.535 ;
      RECT 542.615 -914.965 542.945 -914.635 ;
      RECT 542.63 -1025.18 542.93 -914.635 ;
      RECT 542 -909.325 542.33 -908.995 ;
      RECT 542.015 -1025.18 542.315 -908.995 ;
      RECT 535.115 -876.73 535.445 -876.4 ;
      RECT 535.13 -892.16 535.43 -876.4 ;
      RECT 535.115 -892.16 535.445 -891.83 ;
      RECT 535.13 -872.945 535.43 -829.2 ;
      RECT 535.115 -831.175 535.445 -830.845 ;
      RECT 535.115 -872.535 535.445 -872.205 ;
      RECT 534.515 -908.04 534.815 -840.46 ;
      RECT 534.5 -840.835 534.83 -840.505 ;
      RECT 534.5 -860.315 534.83 -859.985 ;
      RECT 534.5 -908.04 534.83 -907.71 ;
      RECT 533.9 -855.655 534.2 -841.09 ;
      RECT 533.885 -841.465 534.215 -841.135 ;
      RECT 533.885 -855.655 534.215 -855.325 ;
      RECT 533.27 -903.135 533.6 -902.805 ;
      RECT 533.285 -1025.18 533.585 -902.805 ;
      RECT 533.27 -877.19 533.6 -876.86 ;
      RECT 533.285 -892.16 533.585 -876.86 ;
      RECT 533.27 -892.16 533.6 -891.83 ;
      RECT 533.285 -872.965 533.585 -829.2 ;
      RECT 533.27 -829.575 533.6 -829.245 ;
      RECT 533.27 -872.965 533.6 -872.635 ;
      RECT 516.3 -924.89 516.6 -845.185 ;
      RECT 516.285 -845.56 516.615 -845.23 ;
      RECT 516.285 -924.89 516.615 -924.56 ;
      RECT 515.115 -876.73 515.445 -876.4 ;
      RECT 515.13 -892.16 515.43 -876.4 ;
      RECT 515.115 -892.16 515.445 -891.83 ;
      RECT 515.13 -872.945 515.43 -829.2 ;
      RECT 515.115 -831.175 515.445 -830.845 ;
      RECT 515.115 -872.535 515.445 -872.205 ;
      RECT 514.515 -916.05 514.815 -840.46 ;
      RECT 514.5 -840.835 514.83 -840.505 ;
      RECT 514.5 -860.315 514.83 -859.985 ;
      RECT 514.5 -916.05 514.83 -915.72 ;
      RECT 513.9 -855.655 514.2 -841.09 ;
      RECT 513.885 -841.465 514.215 -841.135 ;
      RECT 513.885 -855.655 514.215 -855.325 ;
      RECT 513.27 -903.135 513.6 -902.805 ;
      RECT 513.285 -1025.18 513.585 -902.805 ;
      RECT 513.27 -877.19 513.6 -876.86 ;
      RECT 513.285 -892.16 513.585 -876.86 ;
      RECT 513.27 -892.16 513.6 -891.83 ;
      RECT 513.285 -872.965 513.585 -829.2 ;
      RECT 513.27 -829.575 513.6 -829.245 ;
      RECT 513.27 -872.965 513.6 -872.635 ;
      RECT 504.11 -925.265 504.44 -924.935 ;
      RECT 504.125 -1025.18 504.425 -924.935 ;
      RECT 503.245 -908.525 503.575 -908.195 ;
      RECT 503.26 -1017.91 503.56 -908.195 ;
      RECT 503.245 -915.765 503.575 -915.435 ;
      RECT 503.245 -924.465 503.575 -924.135 ;
      RECT 503.245 -1017.865 503.575 -1017.535 ;
      RECT 502.615 -914.965 502.945 -914.635 ;
      RECT 502.63 -1025.18 502.93 -914.635 ;
      RECT 502 -909.325 502.33 -908.995 ;
      RECT 502.015 -1025.18 502.315 -908.995 ;
      RECT 495.115 -876.73 495.445 -876.4 ;
      RECT 495.13 -892.16 495.43 -876.4 ;
      RECT 495.115 -892.16 495.445 -891.83 ;
      RECT 495.13 -872.945 495.43 -829.2 ;
      RECT 495.115 -831.175 495.445 -830.845 ;
      RECT 495.115 -872.535 495.445 -872.205 ;
      RECT 494.515 -908.04 494.815 -840.46 ;
      RECT 494.5 -840.835 494.83 -840.505 ;
      RECT 494.5 -860.315 494.83 -859.985 ;
      RECT 494.5 -908.04 494.83 -907.71 ;
      RECT 493.9 -855.655 494.2 -841.09 ;
      RECT 493.885 -841.465 494.215 -841.135 ;
      RECT 493.885 -855.655 494.215 -855.325 ;
      RECT 493.27 -903.135 493.6 -902.805 ;
      RECT 493.285 -1025.18 493.585 -902.805 ;
      RECT 493.27 -877.19 493.6 -876.86 ;
      RECT 493.285 -892.16 493.585 -876.86 ;
      RECT 493.27 -892.16 493.6 -891.83 ;
      RECT 493.285 -872.965 493.585 -829.2 ;
      RECT 493.27 -829.575 493.6 -829.245 ;
      RECT 493.27 -872.965 493.6 -872.635 ;
      RECT 475.115 -876.73 475.445 -876.4 ;
      RECT 475.13 -892.16 475.43 -876.4 ;
      RECT 475.115 -892.16 475.445 -891.83 ;
      RECT 475.13 -872.945 475.43 -829.2 ;
      RECT 475.115 -831.175 475.445 -830.845 ;
      RECT 475.115 -872.535 475.445 -872.205 ;
      RECT 474.515 -916.05 474.815 -840.46 ;
      RECT 474.5 -840.835 474.83 -840.505 ;
      RECT 474.5 -860.315 474.83 -859.985 ;
      RECT 474.5 -916.05 474.83 -915.72 ;
      RECT 473.9 -855.655 474.2 -841.09 ;
      RECT 473.885 -841.465 474.215 -841.135 ;
      RECT 473.885 -855.655 474.215 -855.325 ;
      RECT 473.27 -903.135 473.6 -902.805 ;
      RECT 473.285 -1025.18 473.585 -902.805 ;
      RECT 473.27 -877.19 473.6 -876.86 ;
      RECT 473.285 -892.16 473.585 -876.86 ;
      RECT 473.27 -892.16 473.6 -891.83 ;
      RECT 473.285 -872.965 473.585 -829.2 ;
      RECT 473.27 -829.575 473.6 -829.245 ;
      RECT 473.27 -872.965 473.6 -872.635 ;
      RECT 463.245 -908.525 463.575 -908.195 ;
      RECT 463.26 -1017.91 463.56 -908.195 ;
      RECT 463.245 -915.765 463.575 -915.435 ;
      RECT 463.245 -1017.865 463.575 -1017.535 ;
      RECT 462.615 -914.965 462.945 -914.635 ;
      RECT 462.63 -1025.18 462.93 -914.635 ;
      RECT 462 -909.325 462.33 -908.995 ;
      RECT 462.015 -1025.18 462.315 -908.995 ;
      RECT 455.115 -876.73 455.445 -876.4 ;
      RECT 455.13 -892.16 455.43 -876.4 ;
      RECT 455.115 -892.16 455.445 -891.83 ;
      RECT 455.13 -872.945 455.43 -829.2 ;
      RECT 455.115 -831.175 455.445 -830.845 ;
      RECT 455.115 -872.535 455.445 -872.205 ;
      RECT 454.515 -908.04 454.815 -840.46 ;
      RECT 454.5 -840.835 454.83 -840.505 ;
      RECT 454.5 -860.315 454.83 -859.985 ;
      RECT 454.5 -908.04 454.83 -907.71 ;
      RECT 453.9 -855.655 454.2 -841.09 ;
      RECT 453.885 -841.465 454.215 -841.135 ;
      RECT 453.885 -855.655 454.215 -855.325 ;
      RECT 453.27 -903.135 453.6 -902.805 ;
      RECT 453.285 -1025.18 453.585 -902.805 ;
      RECT 453.27 -877.19 453.6 -876.86 ;
      RECT 453.285 -892.16 453.585 -876.86 ;
      RECT 453.27 -892.16 453.6 -891.83 ;
      RECT 453.285 -872.965 453.585 -829.2 ;
      RECT 453.27 -829.575 453.6 -829.245 ;
      RECT 453.27 -872.965 453.6 -872.635 ;
      RECT 435.115 -876.73 435.445 -876.4 ;
      RECT 435.13 -892.16 435.43 -876.4 ;
      RECT 435.115 -892.16 435.445 -891.83 ;
      RECT 435.13 -872.945 435.43 -829.2 ;
      RECT 435.115 -831.175 435.445 -830.845 ;
      RECT 435.115 -872.535 435.445 -872.205 ;
      RECT 434.515 -916.05 434.815 -840.46 ;
      RECT 434.5 -840.835 434.83 -840.505 ;
      RECT 434.5 -860.315 434.83 -859.985 ;
      RECT 434.5 -916.05 434.83 -915.72 ;
      RECT 433.9 -855.655 434.2 -841.09 ;
      RECT 433.885 -841.465 434.215 -841.135 ;
      RECT 433.885 -855.655 434.215 -855.325 ;
      RECT 433.27 -903.135 433.6 -902.805 ;
      RECT 433.285 -1025.18 433.585 -902.805 ;
      RECT 433.27 -877.19 433.6 -876.86 ;
      RECT 433.285 -892.16 433.585 -876.86 ;
      RECT 433.27 -892.16 433.6 -891.83 ;
      RECT 433.285 -872.965 433.585 -829.2 ;
      RECT 433.27 -829.575 433.6 -829.245 ;
      RECT 433.27 -872.965 433.6 -872.635 ;
      RECT 423.245 -908.525 423.575 -908.195 ;
      RECT 423.26 -1017.91 423.56 -908.195 ;
      RECT 423.245 -915.765 423.575 -915.435 ;
      RECT 423.245 -1017.865 423.575 -1017.535 ;
      RECT 422.615 -914.965 422.945 -914.635 ;
      RECT 422.63 -1025.18 422.93 -914.635 ;
      RECT 422 -909.325 422.33 -908.995 ;
      RECT 422.015 -1025.18 422.315 -908.995 ;
      RECT 415.115 -876.73 415.445 -876.4 ;
      RECT 415.13 -892.16 415.43 -876.4 ;
      RECT 415.115 -892.16 415.445 -891.83 ;
      RECT 415.13 -872.945 415.43 -829.2 ;
      RECT 415.115 -831.175 415.445 -830.845 ;
      RECT 415.115 -872.535 415.445 -872.205 ;
      RECT 414.515 -908.04 414.815 -840.46 ;
      RECT 414.5 -840.835 414.83 -840.505 ;
      RECT 414.5 -860.315 414.83 -859.985 ;
      RECT 414.5 -908.04 414.83 -907.71 ;
      RECT 413.9 -855.655 414.2 -841.09 ;
      RECT 413.885 -841.465 414.215 -841.135 ;
      RECT 413.885 -855.655 414.215 -855.325 ;
      RECT 413.27 -903.135 413.6 -902.805 ;
      RECT 413.285 -1025.18 413.585 -902.805 ;
      RECT 413.27 -877.19 413.6 -876.86 ;
      RECT 413.285 -892.16 413.585 -876.86 ;
      RECT 413.27 -892.16 413.6 -891.83 ;
      RECT 413.285 -872.965 413.585 -829.2 ;
      RECT 413.27 -829.575 413.6 -829.245 ;
      RECT 413.27 -872.965 413.6 -872.635 ;
      RECT 395.115 -876.73 395.445 -876.4 ;
      RECT 395.13 -892.16 395.43 -876.4 ;
      RECT 395.115 -892.16 395.445 -891.83 ;
      RECT 395.13 -872.945 395.43 -829.2 ;
      RECT 395.115 -831.175 395.445 -830.845 ;
      RECT 395.115 -872.535 395.445 -872.205 ;
      RECT 394.515 -916.05 394.815 -840.46 ;
      RECT 394.5 -840.835 394.83 -840.505 ;
      RECT 394.5 -860.315 394.83 -859.985 ;
      RECT 394.5 -916.05 394.83 -915.72 ;
      RECT 393.9 -855.655 394.2 -841.09 ;
      RECT 393.885 -841.465 394.215 -841.135 ;
      RECT 393.885 -855.655 394.215 -855.325 ;
      RECT 393.27 -903.135 393.6 -902.805 ;
      RECT 393.285 -1025.18 393.585 -902.805 ;
      RECT 393.27 -877.19 393.6 -876.86 ;
      RECT 393.285 -892.16 393.585 -876.86 ;
      RECT 393.27 -892.16 393.6 -891.83 ;
      RECT 393.285 -872.965 393.585 -829.2 ;
      RECT 393.27 -829.575 393.6 -829.245 ;
      RECT 393.27 -872.965 393.6 -872.635 ;
      RECT 383.245 -908.525 383.575 -908.195 ;
      RECT 383.26 -1017.91 383.56 -908.195 ;
      RECT 383.245 -915.765 383.575 -915.435 ;
      RECT 383.245 -1017.865 383.575 -1017.535 ;
      RECT 382.615 -914.965 382.945 -914.635 ;
      RECT 382.63 -1025.18 382.93 -914.635 ;
      RECT 382 -909.325 382.33 -908.995 ;
      RECT 382.015 -1025.18 382.315 -908.995 ;
      RECT 375.115 -876.73 375.445 -876.4 ;
      RECT 375.13 -892.16 375.43 -876.4 ;
      RECT 375.115 -892.16 375.445 -891.83 ;
      RECT 375.13 -872.945 375.43 -829.2 ;
      RECT 375.115 -831.175 375.445 -830.845 ;
      RECT 375.115 -872.535 375.445 -872.205 ;
      RECT 374.515 -908.04 374.815 -840.46 ;
      RECT 374.5 -840.835 374.83 -840.505 ;
      RECT 374.5 -860.315 374.83 -859.985 ;
      RECT 374.5 -908.04 374.83 -907.71 ;
      RECT 373.9 -855.655 374.2 -841.09 ;
      RECT 373.885 -841.465 374.215 -841.135 ;
      RECT 373.885 -855.655 374.215 -855.325 ;
      RECT 373.27 -903.135 373.6 -902.805 ;
      RECT 373.285 -1025.18 373.585 -902.805 ;
      RECT 373.27 -877.19 373.6 -876.86 ;
      RECT 373.285 -892.16 373.585 -876.86 ;
      RECT 373.27 -892.16 373.6 -891.83 ;
      RECT 373.285 -872.965 373.585 -829.2 ;
      RECT 373.27 -829.575 373.6 -829.245 ;
      RECT 373.27 -872.965 373.6 -872.635 ;
      RECT 356.3 -924.89 356.6 -845.185 ;
      RECT 356.285 -845.56 356.615 -845.23 ;
      RECT 356.285 -924.89 356.615 -924.56 ;
      RECT 355.115 -876.73 355.445 -876.4 ;
      RECT 355.13 -892.16 355.43 -876.4 ;
      RECT 355.115 -892.16 355.445 -891.83 ;
      RECT 355.13 -872.945 355.43 -829.2 ;
      RECT 355.115 -831.175 355.445 -830.845 ;
      RECT 355.115 -872.535 355.445 -872.205 ;
      RECT 354.515 -916.05 354.815 -840.46 ;
      RECT 354.5 -840.835 354.83 -840.505 ;
      RECT 354.5 -860.315 354.83 -859.985 ;
      RECT 354.5 -916.05 354.83 -915.72 ;
      RECT 353.9 -855.655 354.2 -841.09 ;
      RECT 353.885 -841.465 354.215 -841.135 ;
      RECT 353.885 -855.655 354.215 -855.325 ;
      RECT 353.27 -903.135 353.6 -902.805 ;
      RECT 353.285 -1025.18 353.585 -902.805 ;
      RECT 353.27 -877.19 353.6 -876.86 ;
      RECT 353.285 -892.16 353.585 -876.86 ;
      RECT 353.27 -892.16 353.6 -891.83 ;
      RECT 353.285 -872.965 353.585 -829.2 ;
      RECT 353.27 -829.575 353.6 -829.245 ;
      RECT 353.27 -872.965 353.6 -872.635 ;
      RECT 344.11 -925.265 344.44 -924.935 ;
      RECT 344.125 -1025.18 344.425 -924.935 ;
      RECT 343.245 -908.525 343.575 -908.195 ;
      RECT 343.26 -1017.91 343.56 -908.195 ;
      RECT 343.245 -915.765 343.575 -915.435 ;
      RECT 343.245 -924.465 343.575 -924.135 ;
      RECT 343.245 -1017.865 343.575 -1017.535 ;
      RECT 342.615 -914.965 342.945 -914.635 ;
      RECT 342.63 -1025.18 342.93 -914.635 ;
      RECT 342 -909.325 342.33 -908.995 ;
      RECT 342.015 -1025.18 342.315 -908.995 ;
      RECT 335.115 -876.73 335.445 -876.4 ;
      RECT 335.13 -892.16 335.43 -876.4 ;
      RECT 335.115 -892.16 335.445 -891.83 ;
      RECT 335.13 -872.945 335.43 -829.2 ;
      RECT 335.115 -831.175 335.445 -830.845 ;
      RECT 335.115 -872.535 335.445 -872.205 ;
      RECT 334.515 -908.04 334.815 -840.46 ;
      RECT 334.5 -840.835 334.83 -840.505 ;
      RECT 334.5 -860.315 334.83 -859.985 ;
      RECT 334.5 -908.04 334.83 -907.71 ;
      RECT 333.9 -855.655 334.2 -841.09 ;
      RECT 333.885 -841.465 334.215 -841.135 ;
      RECT 333.885 -855.655 334.215 -855.325 ;
      RECT 333.27 -903.135 333.6 -902.805 ;
      RECT 333.285 -1025.18 333.585 -902.805 ;
      RECT 333.27 -877.19 333.6 -876.86 ;
      RECT 333.285 -892.16 333.585 -876.86 ;
      RECT 333.27 -892.16 333.6 -891.83 ;
      RECT 333.285 -872.965 333.585 -829.2 ;
      RECT 333.27 -829.575 333.6 -829.245 ;
      RECT 333.27 -872.965 333.6 -872.635 ;
      RECT 315.115 -876.73 315.445 -876.4 ;
      RECT 315.13 -892.16 315.43 -876.4 ;
      RECT 315.115 -892.16 315.445 -891.83 ;
      RECT 315.13 -872.945 315.43 -829.2 ;
      RECT 315.115 -831.175 315.445 -830.845 ;
      RECT 315.115 -872.535 315.445 -872.205 ;
      RECT 314.515 -916.05 314.815 -840.46 ;
      RECT 314.5 -840.835 314.83 -840.505 ;
      RECT 314.5 -860.315 314.83 -859.985 ;
      RECT 314.5 -916.05 314.83 -915.72 ;
      RECT 313.9 -855.655 314.2 -841.09 ;
      RECT 313.885 -841.465 314.215 -841.135 ;
      RECT 313.885 -855.655 314.215 -855.325 ;
      RECT 313.27 -903.135 313.6 -902.805 ;
      RECT 313.285 -1025.18 313.585 -902.805 ;
      RECT 313.27 -877.19 313.6 -876.86 ;
      RECT 313.285 -892.16 313.585 -876.86 ;
      RECT 313.27 -892.16 313.6 -891.83 ;
      RECT 313.285 -872.965 313.585 -829.2 ;
      RECT 313.27 -829.575 313.6 -829.245 ;
      RECT 313.27 -872.965 313.6 -872.635 ;
      RECT 303.245 -908.525 303.575 -908.195 ;
      RECT 303.26 -1017.91 303.56 -908.195 ;
      RECT 303.245 -915.765 303.575 -915.435 ;
      RECT 303.245 -1017.865 303.575 -1017.535 ;
      RECT 302.615 -914.965 302.945 -914.635 ;
      RECT 302.63 -1025.18 302.93 -914.635 ;
      RECT 302 -909.325 302.33 -908.995 ;
      RECT 302.015 -1025.18 302.315 -908.995 ;
      RECT 295.115 -876.73 295.445 -876.4 ;
      RECT 295.13 -892.16 295.43 -876.4 ;
      RECT 295.115 -892.16 295.445 -891.83 ;
      RECT 295.13 -872.945 295.43 -829.2 ;
      RECT 295.115 -831.175 295.445 -830.845 ;
      RECT 295.115 -872.535 295.445 -872.205 ;
      RECT 294.515 -908.04 294.815 -840.46 ;
      RECT 294.5 -840.835 294.83 -840.505 ;
      RECT 294.5 -860.315 294.83 -859.985 ;
      RECT 294.5 -908.04 294.83 -907.71 ;
      RECT 293.9 -855.655 294.2 -841.09 ;
      RECT 293.885 -841.465 294.215 -841.135 ;
      RECT 293.885 -855.655 294.215 -855.325 ;
      RECT 293.27 -903.135 293.6 -902.805 ;
      RECT 293.285 -1025.18 293.585 -902.805 ;
      RECT 293.27 -877.19 293.6 -876.86 ;
      RECT 293.285 -892.16 293.585 -876.86 ;
      RECT 293.27 -892.16 293.6 -891.83 ;
      RECT 293.285 -872.965 293.585 -829.2 ;
      RECT 293.27 -829.575 293.6 -829.245 ;
      RECT 293.27 -872.965 293.6 -872.635 ;
      RECT 275.115 -876.73 275.445 -876.4 ;
      RECT 275.13 -892.16 275.43 -876.4 ;
      RECT 275.115 -892.16 275.445 -891.83 ;
      RECT 275.13 -872.945 275.43 -829.2 ;
      RECT 275.115 -831.175 275.445 -830.845 ;
      RECT 275.115 -872.535 275.445 -872.205 ;
      RECT 274.515 -916.05 274.815 -840.46 ;
      RECT 274.5 -840.835 274.83 -840.505 ;
      RECT 274.5 -860.315 274.83 -859.985 ;
      RECT 274.5 -916.05 274.83 -915.72 ;
      RECT 273.9 -855.655 274.2 -841.09 ;
      RECT 273.885 -841.465 274.215 -841.135 ;
      RECT 273.885 -855.655 274.215 -855.325 ;
      RECT 273.27 -903.135 273.6 -902.805 ;
      RECT 273.285 -1025.18 273.585 -902.805 ;
      RECT 273.27 -877.19 273.6 -876.86 ;
      RECT 273.285 -892.16 273.585 -876.86 ;
      RECT 273.27 -892.16 273.6 -891.83 ;
      RECT 273.285 -872.965 273.585 -829.2 ;
      RECT 273.27 -829.575 273.6 -829.245 ;
      RECT 273.27 -872.965 273.6 -872.635 ;
      RECT 263.245 -908.525 263.575 -908.195 ;
      RECT 263.26 -1017.91 263.56 -908.195 ;
      RECT 263.245 -915.765 263.575 -915.435 ;
      RECT 263.245 -1017.865 263.575 -1017.535 ;
      RECT 262.615 -914.965 262.945 -914.635 ;
      RECT 262.63 -1025.18 262.93 -914.635 ;
      RECT 262 -909.325 262.33 -908.995 ;
      RECT 262.015 -1025.18 262.315 -908.995 ;
      RECT 255.115 -876.73 255.445 -876.4 ;
      RECT 255.13 -892.16 255.43 -876.4 ;
      RECT 255.115 -892.16 255.445 -891.83 ;
      RECT 255.13 -872.945 255.43 -829.2 ;
      RECT 255.115 -831.175 255.445 -830.845 ;
      RECT 255.115 -872.535 255.445 -872.205 ;
      RECT 254.515 -908.04 254.815 -840.46 ;
      RECT 254.5 -840.835 254.83 -840.505 ;
      RECT 254.5 -860.315 254.83 -859.985 ;
      RECT 254.5 -908.04 254.83 -907.71 ;
      RECT 253.9 -855.655 254.2 -841.09 ;
      RECT 253.885 -841.465 254.215 -841.135 ;
      RECT 253.885 -855.655 254.215 -855.325 ;
      RECT 253.27 -903.135 253.6 -902.805 ;
      RECT 253.285 -1025.18 253.585 -902.805 ;
      RECT 253.27 -877.19 253.6 -876.86 ;
      RECT 253.285 -892.16 253.585 -876.86 ;
      RECT 253.27 -892.16 253.6 -891.83 ;
      RECT 253.285 -872.965 253.585 -829.2 ;
      RECT 253.27 -829.575 253.6 -829.245 ;
      RECT 253.27 -872.965 253.6 -872.635 ;
      RECT 235.115 -876.73 235.445 -876.4 ;
      RECT 235.13 -892.16 235.43 -876.4 ;
      RECT 235.115 -892.16 235.445 -891.83 ;
      RECT 235.13 -872.945 235.43 -829.2 ;
      RECT 235.115 -831.175 235.445 -830.845 ;
      RECT 235.115 -872.535 235.445 -872.205 ;
      RECT 234.515 -916.05 234.815 -840.46 ;
      RECT 234.5 -840.835 234.83 -840.505 ;
      RECT 234.5 -860.315 234.83 -859.985 ;
      RECT 234.5 -916.05 234.83 -915.72 ;
      RECT 233.9 -855.655 234.2 -841.09 ;
      RECT 233.885 -841.465 234.215 -841.135 ;
      RECT 233.885 -855.655 234.215 -855.325 ;
      RECT 233.27 -903.135 233.6 -902.805 ;
      RECT 233.285 -1025.18 233.585 -902.805 ;
      RECT 233.27 -877.19 233.6 -876.86 ;
      RECT 233.285 -892.16 233.585 -876.86 ;
      RECT 233.27 -892.16 233.6 -891.83 ;
      RECT 233.285 -872.965 233.585 -829.2 ;
      RECT 233.27 -829.575 233.6 -829.245 ;
      RECT 233.27 -872.965 233.6 -872.635 ;
      RECT 223.245 -908.525 223.575 -908.195 ;
      RECT 223.26 -1017.91 223.56 -908.195 ;
      RECT 223.245 -915.765 223.575 -915.435 ;
      RECT 223.245 -1017.865 223.575 -1017.535 ;
      RECT 222.615 -914.965 222.945 -914.635 ;
      RECT 222.63 -1025.18 222.93 -914.635 ;
      RECT 222 -909.325 222.33 -908.995 ;
      RECT 222.015 -1025.18 222.315 -908.995 ;
      RECT 215.115 -876.73 215.445 -876.4 ;
      RECT 215.13 -892.16 215.43 -876.4 ;
      RECT 215.115 -892.16 215.445 -891.83 ;
      RECT 215.13 -872.945 215.43 -829.2 ;
      RECT 215.115 -831.175 215.445 -830.845 ;
      RECT 215.115 -872.535 215.445 -872.205 ;
      RECT 214.515 -908.04 214.815 -840.46 ;
      RECT 214.5 -840.835 214.83 -840.505 ;
      RECT 214.5 -860.315 214.83 -859.985 ;
      RECT 214.5 -908.04 214.83 -907.71 ;
      RECT 213.9 -855.655 214.2 -841.09 ;
      RECT 213.885 -841.465 214.215 -841.135 ;
      RECT 213.885 -855.655 214.215 -855.325 ;
      RECT 213.27 -903.135 213.6 -902.805 ;
      RECT 213.285 -1025.18 213.585 -902.805 ;
      RECT 213.27 -877.19 213.6 -876.86 ;
      RECT 213.285 -892.16 213.585 -876.86 ;
      RECT 213.27 -892.16 213.6 -891.83 ;
      RECT 213.285 -872.965 213.585 -829.2 ;
      RECT 213.27 -829.575 213.6 -829.245 ;
      RECT 213.27 -872.965 213.6 -872.635 ;
      RECT 196.3 -924.89 196.6 -845.185 ;
      RECT 196.285 -845.56 196.615 -845.23 ;
      RECT 196.285 -924.89 196.615 -924.56 ;
      RECT 195.115 -876.73 195.445 -876.4 ;
      RECT 195.13 -892.16 195.43 -876.4 ;
      RECT 195.115 -892.16 195.445 -891.83 ;
      RECT 195.13 -872.945 195.43 -829.2 ;
      RECT 195.115 -831.175 195.445 -830.845 ;
      RECT 195.115 -872.535 195.445 -872.205 ;
      RECT 194.515 -916.05 194.815 -840.46 ;
      RECT 194.5 -840.835 194.83 -840.505 ;
      RECT 194.5 -860.315 194.83 -859.985 ;
      RECT 194.5 -916.05 194.83 -915.72 ;
      RECT 193.9 -855.655 194.2 -841.09 ;
      RECT 193.885 -841.465 194.215 -841.135 ;
      RECT 193.885 -855.655 194.215 -855.325 ;
      RECT 193.27 -903.135 193.6 -902.805 ;
      RECT 193.285 -1025.18 193.585 -902.805 ;
      RECT 193.27 -877.19 193.6 -876.86 ;
      RECT 193.285 -892.16 193.585 -876.86 ;
      RECT 193.27 -892.16 193.6 -891.83 ;
      RECT 193.285 -872.965 193.585 -829.2 ;
      RECT 193.27 -829.575 193.6 -829.245 ;
      RECT 193.27 -872.965 193.6 -872.635 ;
      RECT 184.11 -925.265 184.44 -924.935 ;
      RECT 184.125 -1025.18 184.425 -924.935 ;
      RECT 183.245 -908.525 183.575 -908.195 ;
      RECT 183.26 -1017.91 183.56 -908.195 ;
      RECT 183.245 -915.765 183.575 -915.435 ;
      RECT 183.245 -924.465 183.575 -924.135 ;
      RECT 183.245 -1017.865 183.575 -1017.535 ;
      RECT 182.615 -914.965 182.945 -914.635 ;
      RECT 182.63 -1025.18 182.93 -914.635 ;
      RECT 182 -909.325 182.33 -908.995 ;
      RECT 182.015 -1025.18 182.315 -908.995 ;
      RECT 175.115 -876.73 175.445 -876.4 ;
      RECT 175.13 -892.16 175.43 -876.4 ;
      RECT 175.115 -892.16 175.445 -891.83 ;
      RECT 175.13 -872.945 175.43 -829.2 ;
      RECT 175.115 -831.175 175.445 -830.845 ;
      RECT 175.115 -872.535 175.445 -872.205 ;
      RECT 174.515 -908.04 174.815 -840.46 ;
      RECT 174.5 -840.835 174.83 -840.505 ;
      RECT 174.5 -860.315 174.83 -859.985 ;
      RECT 174.5 -908.04 174.83 -907.71 ;
      RECT 173.9 -855.655 174.2 -841.09 ;
      RECT 173.885 -841.465 174.215 -841.135 ;
      RECT 173.885 -855.655 174.215 -855.325 ;
      RECT 173.27 -903.135 173.6 -902.805 ;
      RECT 173.285 -1025.18 173.585 -902.805 ;
      RECT 173.27 -877.19 173.6 -876.86 ;
      RECT 173.285 -892.16 173.585 -876.86 ;
      RECT 173.27 -892.16 173.6 -891.83 ;
      RECT 173.285 -872.965 173.585 -829.2 ;
      RECT 173.27 -829.575 173.6 -829.245 ;
      RECT 173.27 -872.965 173.6 -872.635 ;
      RECT 155.115 -876.73 155.445 -876.4 ;
      RECT 155.13 -892.16 155.43 -876.4 ;
      RECT 155.115 -892.16 155.445 -891.83 ;
      RECT 155.13 -872.945 155.43 -829.2 ;
      RECT 155.115 -831.175 155.445 -830.845 ;
      RECT 155.115 -872.535 155.445 -872.205 ;
      RECT 154.515 -916.05 154.815 -840.46 ;
      RECT 154.5 -840.835 154.83 -840.505 ;
      RECT 154.5 -860.315 154.83 -859.985 ;
      RECT 154.5 -916.05 154.83 -915.72 ;
      RECT 153.9 -855.655 154.2 -841.09 ;
      RECT 153.885 -841.465 154.215 -841.135 ;
      RECT 153.885 -855.655 154.215 -855.325 ;
      RECT 153.27 -903.135 153.6 -902.805 ;
      RECT 153.285 -1025.18 153.585 -902.805 ;
      RECT 153.27 -877.19 153.6 -876.86 ;
      RECT 153.285 -892.16 153.585 -876.86 ;
      RECT 153.27 -892.16 153.6 -891.83 ;
      RECT 153.285 -872.965 153.585 -829.2 ;
      RECT 153.27 -829.575 153.6 -829.245 ;
      RECT 153.27 -872.965 153.6 -872.635 ;
      RECT 143.245 -908.525 143.575 -908.195 ;
      RECT 143.26 -1017.91 143.56 -908.195 ;
      RECT 143.245 -915.765 143.575 -915.435 ;
      RECT 143.245 -1017.865 143.575 -1017.535 ;
      RECT 142.615 -914.965 142.945 -914.635 ;
      RECT 142.63 -1025.18 142.93 -914.635 ;
      RECT 142 -909.325 142.33 -908.995 ;
      RECT 142.015 -1025.18 142.315 -908.995 ;
      RECT 135.115 -876.73 135.445 -876.4 ;
      RECT 135.13 -892.16 135.43 -876.4 ;
      RECT 135.115 -892.16 135.445 -891.83 ;
      RECT 135.13 -872.945 135.43 -829.2 ;
      RECT 135.115 -831.175 135.445 -830.845 ;
      RECT 135.115 -872.535 135.445 -872.205 ;
      RECT 134.515 -908.04 134.815 -840.46 ;
      RECT 134.5 -840.835 134.83 -840.505 ;
      RECT 134.5 -860.315 134.83 -859.985 ;
      RECT 134.5 -908.04 134.83 -907.71 ;
      RECT 133.9 -855.655 134.2 -841.09 ;
      RECT 133.885 -841.465 134.215 -841.135 ;
      RECT 133.885 -855.655 134.215 -855.325 ;
      RECT 133.27 -903.135 133.6 -902.805 ;
      RECT 133.285 -1025.18 133.585 -902.805 ;
      RECT 133.27 -877.19 133.6 -876.86 ;
      RECT 133.285 -892.16 133.585 -876.86 ;
      RECT 133.27 -892.16 133.6 -891.83 ;
      RECT 133.285 -872.965 133.585 -829.2 ;
      RECT 133.27 -829.575 133.6 -829.245 ;
      RECT 133.27 -872.965 133.6 -872.635 ;
      RECT 115.115 -876.73 115.445 -876.4 ;
      RECT 115.13 -892.16 115.43 -876.4 ;
      RECT 115.115 -892.16 115.445 -891.83 ;
      RECT 115.13 -872.945 115.43 -829.2 ;
      RECT 115.115 -831.175 115.445 -830.845 ;
      RECT 115.115 -872.535 115.445 -872.205 ;
      RECT 114.515 -916.05 114.815 -840.46 ;
      RECT 114.5 -840.835 114.83 -840.505 ;
      RECT 114.5 -860.315 114.83 -859.985 ;
      RECT 114.5 -916.05 114.83 -915.72 ;
      RECT 113.9 -855.655 114.2 -841.09 ;
      RECT 113.885 -841.465 114.215 -841.135 ;
      RECT 113.885 -855.655 114.215 -855.325 ;
      RECT 113.27 -903.135 113.6 -902.805 ;
      RECT 113.285 -1025.18 113.585 -902.805 ;
      RECT 113.27 -877.19 113.6 -876.86 ;
      RECT 113.285 -892.16 113.585 -876.86 ;
      RECT 113.27 -892.16 113.6 -891.83 ;
      RECT 113.285 -872.965 113.585 -829.2 ;
      RECT 113.27 -829.575 113.6 -829.245 ;
      RECT 113.27 -872.965 113.6 -872.635 ;
      RECT 103.245 -908.525 103.575 -908.195 ;
      RECT 103.26 -1017.91 103.56 -908.195 ;
      RECT 103.245 -915.765 103.575 -915.435 ;
      RECT 103.245 -1017.865 103.575 -1017.535 ;
      RECT 102.615 -914.965 102.945 -914.635 ;
      RECT 102.63 -1025.18 102.93 -914.635 ;
      RECT 102 -909.325 102.33 -908.995 ;
      RECT 102.015 -1025.18 102.315 -908.995 ;
      RECT 95.115 -876.73 95.445 -876.4 ;
      RECT 95.13 -892.16 95.43 -876.4 ;
      RECT 95.115 -892.16 95.445 -891.83 ;
      RECT 95.13 -872.945 95.43 -829.2 ;
      RECT 95.115 -831.175 95.445 -830.845 ;
      RECT 95.115 -872.535 95.445 -872.205 ;
      RECT 94.515 -908.04 94.815 -840.46 ;
      RECT 94.5 -840.835 94.83 -840.505 ;
      RECT 94.5 -860.315 94.83 -859.985 ;
      RECT 94.5 -908.04 94.83 -907.71 ;
      RECT 93.9 -855.655 94.2 -841.09 ;
      RECT 93.885 -841.465 94.215 -841.135 ;
      RECT 93.885 -855.655 94.215 -855.325 ;
      RECT 93.27 -903.135 93.6 -902.805 ;
      RECT 93.285 -1025.18 93.585 -902.805 ;
      RECT 93.27 -877.19 93.6 -876.86 ;
      RECT 93.285 -892.16 93.585 -876.86 ;
      RECT 93.27 -892.16 93.6 -891.83 ;
      RECT 93.285 -872.965 93.585 -829.2 ;
      RECT 93.27 -829.575 93.6 -829.245 ;
      RECT 93.27 -872.965 93.6 -872.635 ;
      RECT 75.115 -876.73 75.445 -876.4 ;
      RECT 75.13 -892.16 75.43 -876.4 ;
      RECT 75.115 -892.16 75.445 -891.83 ;
      RECT 75.13 -872.945 75.43 -829.2 ;
      RECT 75.115 -831.175 75.445 -830.845 ;
      RECT 75.115 -872.535 75.445 -872.205 ;
      RECT 74.515 -916.05 74.815 -840.46 ;
      RECT 74.5 -840.835 74.83 -840.505 ;
      RECT 74.5 -860.315 74.83 -859.985 ;
      RECT 74.5 -916.05 74.83 -915.72 ;
      RECT 73.9 -855.655 74.2 -841.09 ;
      RECT 73.885 -841.465 74.215 -841.135 ;
      RECT 73.885 -855.655 74.215 -855.325 ;
      RECT 73.27 -903.135 73.6 -902.805 ;
      RECT 73.285 -1025.18 73.585 -902.805 ;
      RECT 73.27 -877.19 73.6 -876.86 ;
      RECT 73.285 -892.16 73.585 -876.86 ;
      RECT 73.27 -892.16 73.6 -891.83 ;
      RECT 73.285 -872.965 73.585 -829.2 ;
      RECT 73.27 -829.575 73.6 -829.245 ;
      RECT 73.27 -872.965 73.6 -872.635 ;
      RECT 63.245 -908.525 63.575 -908.195 ;
      RECT 63.26 -1017.91 63.56 -908.195 ;
      RECT 63.245 -915.765 63.575 -915.435 ;
      RECT 63.245 -1017.865 63.575 -1017.535 ;
      RECT 62.615 -914.965 62.945 -914.635 ;
      RECT 62.63 -1025.18 62.93 -914.635 ;
      RECT 62 -909.325 62.33 -908.995 ;
      RECT 62.015 -1025.18 62.315 -908.995 ;
      RECT 55.115 -876.73 55.445 -876.4 ;
      RECT 55.13 -892.16 55.43 -876.4 ;
      RECT 55.115 -892.16 55.445 -891.83 ;
      RECT 55.13 -872.945 55.43 -829.2 ;
      RECT 55.115 -831.175 55.445 -830.845 ;
      RECT 55.115 -872.535 55.445 -872.205 ;
      RECT 54.515 -908.04 54.815 -840.46 ;
      RECT 54.5 -840.835 54.83 -840.505 ;
      RECT 54.5 -860.315 54.83 -859.985 ;
      RECT 54.5 -908.04 54.83 -907.71 ;
      RECT 53.9 -855.655 54.2 -841.09 ;
      RECT 53.885 -841.465 54.215 -841.135 ;
      RECT 53.885 -855.655 54.215 -855.325 ;
      RECT 53.27 -903.135 53.6 -902.805 ;
      RECT 53.285 -1025.18 53.585 -902.805 ;
      RECT 53.27 -877.19 53.6 -876.86 ;
      RECT 53.285 -892.16 53.585 -876.86 ;
      RECT 53.27 -892.16 53.6 -891.83 ;
      RECT 53.285 -872.965 53.585 -829.2 ;
      RECT 53.27 -829.575 53.6 -829.245 ;
      RECT 53.27 -872.965 53.6 -872.635 ;
      RECT 36.3 -924.89 36.6 -845.185 ;
      RECT 36.285 -845.56 36.615 -845.23 ;
      RECT 36.285 -924.89 36.615 -924.56 ;
      RECT 35.115 -876.73 35.445 -876.4 ;
      RECT 35.13 -892.16 35.43 -876.4 ;
      RECT 35.115 -892.16 35.445 -891.83 ;
      RECT 35.13 -872.945 35.43 -829.2 ;
      RECT 35.115 -831.175 35.445 -830.845 ;
      RECT 35.115 -872.535 35.445 -872.205 ;
      RECT 34.515 -916.05 34.815 -840.46 ;
      RECT 34.5 -840.835 34.83 -840.505 ;
      RECT 34.5 -860.315 34.83 -859.985 ;
      RECT 34.5 -916.05 34.83 -915.72 ;
      RECT 33.9 -855.655 34.2 -841.09 ;
      RECT 33.885 -841.465 34.215 -841.135 ;
      RECT 33.885 -855.655 34.215 -855.325 ;
      RECT 33.27 -903.135 33.6 -902.805 ;
      RECT 33.285 -1025.18 33.585 -902.805 ;
      RECT 33.27 -877.19 33.6 -876.86 ;
      RECT 33.285 -892.16 33.585 -876.86 ;
      RECT 33.27 -892.16 33.6 -891.83 ;
      RECT 33.285 -872.965 33.585 -829.2 ;
      RECT 33.27 -829.575 33.6 -829.245 ;
      RECT 33.27 -872.965 33.6 -872.635 ;
      RECT 24.11 -925.265 24.44 -924.935 ;
      RECT 24.125 -1025.18 24.425 -924.935 ;
      RECT 23.245 -908.525 23.575 -908.195 ;
      RECT 23.26 -1017.91 23.56 -908.195 ;
      RECT 23.245 -915.765 23.575 -915.435 ;
      RECT 23.245 -924.465 23.575 -924.135 ;
      RECT 23.245 -1017.865 23.575 -1017.535 ;
      RECT 22.615 -914.965 22.945 -914.635 ;
      RECT 22.63 -1025.18 22.93 -914.635 ;
      RECT 22 -909.325 22.33 -908.995 ;
      RECT 22.015 -1025.18 22.315 -908.995 ;
      RECT 15.115 -876.73 15.445 -876.4 ;
      RECT 15.13 -892.16 15.43 -876.4 ;
      RECT 15.115 -892.16 15.445 -891.83 ;
      RECT 15.13 -872.945 15.43 -829.2 ;
      RECT 15.115 -831.175 15.445 -830.845 ;
      RECT 15.115 -872.535 15.445 -872.205 ;
      RECT 14.515 -908.04 14.815 -840.46 ;
      RECT 14.5 -840.835 14.83 -840.505 ;
      RECT 14.5 -860.315 14.83 -859.985 ;
      RECT 14.5 -908.04 14.83 -907.71 ;
      RECT 13.9 -855.655 14.2 -841.09 ;
      RECT 13.885 -841.465 14.215 -841.135 ;
      RECT 13.885 -855.655 14.215 -855.325 ;
      RECT 13.27 -903.135 13.6 -902.805 ;
      RECT 13.285 -1025.18 13.585 -902.805 ;
      RECT 13.27 -877.19 13.6 -876.86 ;
      RECT 13.285 -892.16 13.585 -876.86 ;
      RECT 13.27 -892.16 13.6 -891.83 ;
      RECT 13.285 -872.965 13.585 -829.2 ;
      RECT 13.27 -829.575 13.6 -829.245 ;
      RECT 13.27 -872.965 13.6 -872.635 ;
      RECT 11.005 -866.95 11.335 -866.62 ;
      RECT 11.02 -972.98 11.32 -866.62 ;
      RECT 11.005 -972.98 11.335 -972.65 ;
      RECT -5.91 -993.415 -5.58 -993.085 ;
      RECT -5.895 -1013.85 -5.595 -993.085 ;
      RECT -5.91 -1013.85 -5.58 -1013.52 ;
      RECT -9.505 -1013.405 -9.175 -1013.075 ;
      RECT -9.49 -1017.91 -9.19 -1013.075 ;
      RECT -9.505 -1017.865 -9.175 -1017.535 ;
      RECT -10.34 -819.74 -10.01 -819.41 ;
      RECT -10.325 -974.77 -10.025 -819.41 ;
      RECT -10.34 -974.77 -10.01 -974.44 ;
      RECT -10.635 -1014.205 -10.305 -1013.875 ;
      RECT -10.62 -1025.18 -10.32 -1013.875 ;
      RECT -11.75 -998.18 -11.42 -997.85 ;
      RECT -11.735 -1013.85 -11.435 -997.85 ;
      RECT -11.75 -1013.85 -11.42 -1013.52 ;
      RECT -12.385 -997.68 -12.055 -997.35 ;
      RECT -12.37 -1014.605 -12.07 -997.35 ;
      RECT -12.385 -1014.605 -12.055 -1014.275 ;
      RECT -15.345 -1013.405 -15.015 -1013.075 ;
      RECT -15.33 -1017.91 -15.03 -1013.075 ;
      RECT -15.345 -1017.865 -15.015 -1017.535 ;
      RECT -16.475 -1014.205 -16.145 -1013.875 ;
      RECT -16.46 -1025.18 -16.16 -1013.875 ;
      RECT -17.59 -999.18 -17.26 -998.85 ;
      RECT -17.575 -1013.85 -17.275 -998.85 ;
      RECT -17.59 -1013.85 -17.26 -1013.52 ;
      RECT -18.225 -998.68 -17.895 -998.35 ;
      RECT -18.21 -1014.605 -17.91 -998.35 ;
      RECT -18.225 -1014.605 -17.895 -1014.275 ;
      RECT -21.185 -1013.405 -20.855 -1013.075 ;
      RECT -21.17 -1017.91 -20.87 -1013.075 ;
      RECT -21.185 -1017.865 -20.855 -1017.535 ;
      RECT -22.315 -1014.205 -21.985 -1013.875 ;
      RECT -22.3 -1025.18 -22 -1013.875 ;
      RECT -23.43 -1000.18 -23.1 -999.85 ;
      RECT -23.415 -1013.85 -23.115 -999.85 ;
      RECT -23.43 -1013.85 -23.1 -1013.52 ;
      RECT -24.065 -999.68 -23.735 -999.35 ;
      RECT -24.05 -1014.605 -23.75 -999.35 ;
      RECT -24.065 -1014.605 -23.735 -1014.275 ;
      RECT -27.025 -1013.405 -26.695 -1013.075 ;
      RECT -27.01 -1017.91 -26.71 -1013.075 ;
      RECT -27.025 -1017.865 -26.695 -1017.535 ;
      RECT -28.155 -1014.205 -27.825 -1013.875 ;
      RECT -28.14 -1025.18 -27.84 -1013.875 ;
      RECT -29.27 -1001.18 -28.94 -1000.85 ;
      RECT -29.255 -1013.85 -28.955 -1000.85 ;
      RECT -29.27 -1013.85 -28.94 -1013.52 ;
      RECT -29.905 -1000.68 -29.575 -1000.35 ;
      RECT -29.89 -1014.605 -29.59 -1000.35 ;
      RECT -29.905 -1014.605 -29.575 -1014.275 ;
      RECT -32.865 -1013.405 -32.535 -1013.075 ;
      RECT -32.85 -1017.91 -32.55 -1013.075 ;
      RECT -32.865 -1017.865 -32.535 -1017.535 ;
      RECT -33.995 -1014.205 -33.665 -1013.875 ;
      RECT -33.98 -1025.18 -33.68 -1013.875 ;
      RECT -35.11 -1002.18 -34.78 -1001.85 ;
      RECT -35.095 -1013.85 -34.795 -1001.85 ;
      RECT -35.11 -1013.85 -34.78 -1013.52 ;
      RECT -35.745 -1001.68 -35.415 -1001.35 ;
      RECT -35.73 -1014.605 -35.43 -1001.35 ;
      RECT -35.745 -1014.605 -35.415 -1014.275 ;
      RECT -38.705 -1013.405 -38.375 -1013.075 ;
      RECT -38.69 -1017.91 -38.39 -1013.075 ;
      RECT -38.705 -1017.865 -38.375 -1017.535 ;
      RECT -39.835 -1014.205 -39.505 -1013.875 ;
      RECT -39.82 -1025.18 -39.52 -1013.875 ;
      RECT -40.95 -1003.18 -40.62 -1002.85 ;
      RECT -40.935 -1013.85 -40.635 -1002.85 ;
      RECT -40.95 -1013.85 -40.62 -1013.52 ;
      RECT -41.585 -1002.68 -41.255 -1002.35 ;
      RECT -41.57 -1014.605 -41.27 -1002.35 ;
      RECT -41.585 -1014.605 -41.255 -1014.275 ;
      RECT -44.545 -1013.405 -44.215 -1013.075 ;
      RECT -44.53 -1017.91 -44.23 -1013.075 ;
      RECT -44.545 -1017.865 -44.215 -1017.535 ;
      RECT -45.675 -1014.205 -45.345 -1013.875 ;
      RECT -45.66 -1025.18 -45.36 -1013.875 ;
      RECT -46.79 -1004.18 -46.46 -1003.85 ;
      RECT -46.775 -1013.85 -46.475 -1003.85 ;
      RECT -46.79 -1013.85 -46.46 -1013.52 ;
      RECT -47.425 -1003.68 -47.095 -1003.35 ;
      RECT -47.41 -1014.605 -47.11 -1003.35 ;
      RECT -47.425 -1014.605 -47.095 -1014.275 ;
      RECT -50.385 -1013.405 -50.055 -1013.075 ;
      RECT -50.37 -1017.91 -50.07 -1013.075 ;
      RECT -50.385 -1017.865 -50.055 -1017.535 ;
      RECT -51.515 -1014.205 -51.185 -1013.875 ;
      RECT -51.5 -1025.18 -51.2 -1013.875 ;
      RECT -52.63 -1005.18 -52.3 -1004.85 ;
      RECT -52.615 -1013.85 -52.315 -1004.85 ;
      RECT -52.63 -1013.85 -52.3 -1013.52 ;
      RECT -53.265 -1004.68 -52.935 -1004.35 ;
      RECT -53.25 -1014.605 -52.95 -1004.35 ;
      RECT -53.265 -1014.605 -52.935 -1014.275 ;
      RECT -56.225 -1013.405 -55.895 -1013.075 ;
      RECT -56.21 -1017.91 -55.91 -1013.075 ;
      RECT -56.225 -1017.865 -55.895 -1017.535 ;
      RECT -57.355 -1014.205 -57.025 -1013.875 ;
      RECT -57.34 -1025.18 -57.04 -1013.875 ;
      RECT -58.47 -1006.18 -58.14 -1005.85 ;
      RECT -58.455 -1013.85 -58.155 -1005.85 ;
      RECT -58.47 -1013.85 -58.14 -1013.52 ;
      RECT -59.105 -1005.68 -58.775 -1005.35 ;
      RECT -59.09 -1014.605 -58.79 -1005.35 ;
      RECT -59.105 -1014.605 -58.775 -1014.275 ;
      RECT -62.065 -1013.405 -61.735 -1013.075 ;
      RECT -62.05 -1017.91 -61.75 -1013.075 ;
      RECT -62.065 -1017.865 -61.735 -1017.535 ;
      RECT -63.195 -1014.205 -62.865 -1013.875 ;
      RECT -63.18 -1025.18 -62.88 -1013.875 ;
      RECT -64.31 -1007.18 -63.98 -1006.85 ;
      RECT -64.295 -1013.85 -63.995 -1006.85 ;
      RECT -64.31 -1013.85 -63.98 -1013.52 ;
      RECT -64.945 -1006.68 -64.615 -1006.35 ;
      RECT -64.93 -1014.605 -64.63 -1006.35 ;
      RECT -64.945 -1014.605 -64.615 -1014.275 ;
      RECT -67.905 -1013.405 -67.575 -1013.075 ;
      RECT -67.89 -1017.91 -67.59 -1013.075 ;
      RECT -67.905 -1017.865 -67.575 -1017.535 ;
      RECT -69.035 -1014.205 -68.705 -1013.875 ;
      RECT -69.02 -1025.18 -68.72 -1013.875 ;
      RECT -70.15 -1008.18 -69.82 -1007.85 ;
      RECT -70.135 -1013.85 -69.835 -1007.85 ;
      RECT -70.15 -1013.85 -69.82 -1013.52 ;
      RECT -70.785 -1007.68 -70.455 -1007.35 ;
      RECT -70.77 -1014.605 -70.47 -1007.35 ;
      RECT -70.785 -1014.605 -70.455 -1014.275 ;
      RECT -73.745 -1013.405 -73.415 -1013.075 ;
      RECT -73.73 -1017.91 -73.43 -1013.075 ;
      RECT -73.745 -1017.865 -73.415 -1017.535 ;
      RECT -74.875 -1014.205 -74.545 -1013.875 ;
      RECT -74.86 -1025.18 -74.56 -1013.875 ;
      RECT -75.99 -1009.18 -75.66 -1008.85 ;
      RECT -75.975 -1013.85 -75.675 -1008.85 ;
      RECT -75.99 -1013.85 -75.66 -1013.52 ;
      RECT -76.625 -1008.68 -76.295 -1008.35 ;
      RECT -76.61 -1014.605 -76.31 -1008.35 ;
      RECT -76.625 -1014.605 -76.295 -1014.275 ;
      RECT -79.585 -1013.405 -79.255 -1013.075 ;
      RECT -79.57 -1017.91 -79.27 -1013.075 ;
      RECT -79.585 -1017.865 -79.255 -1017.535 ;
      RECT -80.715 -1014.205 -80.385 -1013.875 ;
      RECT -80.7 -1025.18 -80.4 -1013.875 ;
      RECT -81.58 -1017.91 -81.18 -994.725 ;
      RECT -81.72 -1025.06 -81.3 -1017.49 ;
  END
END sramgen_sram_4096x32m8w8_replica_v1

END LIBRARY
